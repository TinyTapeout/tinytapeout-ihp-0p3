module tt_um_a1k0n_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire audio;
 wire hsync;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire \vgademo.a_cos[0] ;
 wire \vgademo.a_cos[10] ;
 wire \vgademo.a_cos[11] ;
 wire \vgademo.a_cos[12] ;
 wire \vgademo.a_cos[13] ;
 wire \vgademo.a_cos[14] ;
 wire \vgademo.a_cos[1] ;
 wire \vgademo.a_cos[2] ;
 wire \vgademo.a_cos[3] ;
 wire \vgademo.a_cos[4] ;
 wire \vgademo.a_cos[5] ;
 wire \vgademo.a_cos[6] ;
 wire \vgademo.a_cos[7] ;
 wire \vgademo.a_cos[8] ;
 wire \vgademo.a_cos[9] ;
 wire \vgademo.a_scrolly[10] ;
 wire \vgademo.a_scrolly[11] ;
 wire \vgademo.a_scrolly[12] ;
 wire \vgademo.a_scrolly[13] ;
 wire \vgademo.a_scrolly[3] ;
 wire \vgademo.a_scrolly[4] ;
 wire \vgademo.a_scrolly[5] ;
 wire \vgademo.a_scrolly[6] ;
 wire \vgademo.a_scrolly[7] ;
 wire \vgademo.a_scrolly[8] ;
 wire \vgademo.a_scrolly[9] ;
 wire \vgademo.a_sin[0] ;
 wire \vgademo.a_sin[10] ;
 wire \vgademo.a_sin[11] ;
 wire \vgademo.a_sin[12] ;
 wire \vgademo.a_sin[13] ;
 wire \vgademo.a_sin[14] ;
 wire \vgademo.a_sin[1] ;
 wire \vgademo.a_sin[2] ;
 wire \vgademo.a_sin[3] ;
 wire \vgademo.a_sin[4] ;
 wire \vgademo.a_sin[5] ;
 wire \vgademo.a_sin[6] ;
 wire \vgademo.a_sin[7] ;
 wire \vgademo.a_sin[8] ;
 wire \vgademo.a_sin[9] ;
 wire \vgademo.audio_beat_out[0] ;
 wire \vgademo.audio_beat_out[1] ;
 wire \vgademo.audio_beat_out[2] ;
 wire \vgademo.audio_beat_out[3] ;
 wire \vgademo.audio_beat_out[4] ;
 wire \vgademo.audio_kick_frames[0] ;
 wire \vgademo.audio_kick_frames[1] ;
 wire \vgademo.audio_kick_frames[2] ;
 wire \vgademo.audio_snare_frames[0] ;
 wire \vgademo.audio_snare_frames[1] ;
 wire \vgademo.audio_snare_frames[2] ;
 wire \vgademo.audio_snare_frames[3] ;
 wire \vgademo.audio_songpos[0] ;
 wire \vgademo.audio_songpos[1] ;
 wire \vgademo.audio_songpos[2] ;
 wire \vgademo.audio_songpos[3] ;
 wire \vgademo.audio_songpos[4] ;
 wire \vgademo.audio_songpos[5] ;
 wire \vgademo.audio_songpos[6] ;
 wire \vgademo.audio_songpos[7] ;
 wire \vgademo.b_cos[0] ;
 wire \vgademo.b_cos[10] ;
 wire \vgademo.b_cos[11] ;
 wire \vgademo.b_cos[1] ;
 wire \vgademo.b_cos[2] ;
 wire \vgademo.b_cos[3] ;
 wire \vgademo.b_cos[4] ;
 wire \vgademo.b_cos[5] ;
 wire \vgademo.b_cos[6] ;
 wire \vgademo.b_cos[7] ;
 wire \vgademo.b_cos[8] ;
 wire \vgademo.b_cos[9] ;
 wire \vgademo.b_sin[0] ;
 wire \vgademo.b_sin[10] ;
 wire \vgademo.b_sin[11] ;
 wire \vgademo.b_sin[1] ;
 wire \vgademo.b_sin[2] ;
 wire \vgademo.b_sin[3] ;
 wire \vgademo.b_sin[4] ;
 wire \vgademo.b_sin[5] ;
 wire \vgademo.b_sin[6] ;
 wire \vgademo.b_sin[7] ;
 wire \vgademo.b_sin[8] ;
 wire \vgademo.b_sin[9] ;
 wire \vgademo.bayer_j[0] ;
 wire \vgademo.bayer_j[1] ;
 wire \vgademo.h_count[0] ;
 wire \vgademo.h_count[10] ;
 wire \vgademo.h_count[1] ;
 wire \vgademo.h_count[2] ;
 wire \vgademo.h_count[3] ;
 wire \vgademo.h_count[4] ;
 wire \vgademo.h_count[5] ;
 wire \vgademo.h_count[6] ;
 wire \vgademo.h_count[7] ;
 wire \vgademo.h_count[8] ;
 wire \vgademo.h_count[9] ;
 wire \vgademo.linelfsr[0] ;
 wire \vgademo.linelfsr[10] ;
 wire \vgademo.linelfsr[11] ;
 wire \vgademo.linelfsr[12] ;
 wire \vgademo.linelfsr[1] ;
 wire \vgademo.linelfsr[2] ;
 wire \vgademo.linelfsr[3] ;
 wire \vgademo.linelfsr[4] ;
 wire \vgademo.linelfsr[5] ;
 wire \vgademo.linelfsr[6] ;
 wire \vgademo.linelfsr[7] ;
 wire \vgademo.linelfsr[8] ;
 wire \vgademo.linelfsr[9] ;
 wire \vgademo.plane_du[0] ;
 wire \vgademo.plane_du[10] ;
 wire \vgademo.plane_du[1] ;
 wire \vgademo.plane_du[2] ;
 wire \vgademo.plane_du[3] ;
 wire \vgademo.plane_du[4] ;
 wire \vgademo.plane_du[5] ;
 wire \vgademo.plane_du[6] ;
 wire \vgademo.plane_du[7] ;
 wire \vgademo.plane_du[8] ;
 wire \vgademo.plane_du[9] ;
 wire \vgademo.plane_dx[0] ;
 wire \vgademo.plane_dx[1] ;
 wire \vgademo.plane_dx[2] ;
 wire \vgademo.plane_dx[3] ;
 wire \vgademo.plane_dx_div.d[16] ;
 wire \vgademo.plane_dx_div.d[17] ;
 wire \vgademo.plane_dx_div.d[18] ;
 wire \vgademo.plane_dx_div.d[19] ;
 wire \vgademo.plane_dx_div.d[20] ;
 wire \vgademo.plane_dx_div.d[21] ;
 wire \vgademo.plane_dx_div.d[22] ;
 wire \vgademo.plane_dx_div.d[23] ;
 wire \vgademo.plane_dx_div.d[24] ;
 wire \vgademo.plane_dx_div.i[0] ;
 wire \vgademo.plane_dx_div.i[1] ;
 wire \vgademo.plane_dx_div.i[2] ;
 wire \vgademo.plane_dx_div.i[3] ;
 wire \vgademo.plane_dx_div.q[3] ;
 wire \vgademo.plane_dx_div.q[4] ;
 wire \vgademo.plane_dx_div.q[5] ;
 wire \vgademo.plane_dx_div.q[6] ;
 wire \vgademo.plane_dx_div.q[7] ;
 wire \vgademo.plane_dx_div.q[8] ;
 wire \vgademo.plane_dx_div.q[9] ;
 wire \vgademo.plane_dx_div.r[16] ;
 wire \vgademo.plane_dx_div.r[17] ;
 wire \vgademo.plane_dx_div.r[18] ;
 wire \vgademo.plane_dx_div.r[19] ;
 wire \vgademo.plane_dx_div.r[20] ;
 wire \vgademo.plane_dx_div.r[21] ;
 wire \vgademo.plane_dx_div.r[22] ;
 wire \vgademo.plane_dx_div.r[23] ;
 wire \vgademo.plane_dx_div.r[24] ;
 wire \vgademo.plane_dx_div.r[25] ;
 wire \vgademo.plane_u[0] ;
 wire \vgademo.plane_u[10] ;
 wire \vgademo.plane_u[11] ;
 wire \vgademo.plane_u[12] ;
 wire \vgademo.plane_u[13] ;
 wire \vgademo.plane_u[14] ;
 wire \vgademo.plane_u[15] ;
 wire \vgademo.plane_u[16] ;
 wire \vgademo.plane_u[17] ;
 wire \vgademo.plane_u[18] ;
 wire \vgademo.plane_u[19] ;
 wire \vgademo.plane_u[1] ;
 wire \vgademo.plane_u[20] ;
 wire \vgademo.plane_u[21] ;
 wire \vgademo.plane_u[2] ;
 wire \vgademo.plane_u[3] ;
 wire \vgademo.plane_u[4] ;
 wire \vgademo.plane_u[5] ;
 wire \vgademo.plane_u[6] ;
 wire \vgademo.plane_u[7] ;
 wire \vgademo.plane_u[8] ;
 wire \vgademo.plane_u[9] ;
 wire \vgademo.scanline_audio_sample[0] ;
 wire \vgademo.scanline_audio_sample[1] ;
 wire \vgademo.scanline_audio_sample[2] ;
 wire \vgademo.scanline_audio_sample[3] ;
 wire \vgademo.scanline_audio_sample[4] ;
 wire \vgademo.scanline_audio_sample[5] ;
 wire \vgademo.scanline_audio_sample[6] ;
 wire \vgademo.soundtrack.noise_lfsr[0] ;
 wire \vgademo.soundtrack.noise_lfsr[10] ;
 wire \vgademo.soundtrack.noise_lfsr[11] ;
 wire \vgademo.soundtrack.noise_lfsr[12] ;
 wire \vgademo.soundtrack.noise_lfsr[13] ;
 wire \vgademo.soundtrack.noise_lfsr[14] ;
 wire \vgademo.soundtrack.noise_lfsr[1] ;
 wire \vgademo.soundtrack.noise_lfsr[2] ;
 wire \vgademo.soundtrack.noise_lfsr[3] ;
 wire \vgademo.soundtrack.noise_lfsr[4] ;
 wire \vgademo.soundtrack.noise_lfsr[5] ;
 wire \vgademo.soundtrack.noise_lfsr[6] ;
 wire \vgademo.soundtrack.noise_lfsr[7] ;
 wire \vgademo.soundtrack.noise_lfsr[8] ;
 wire \vgademo.soundtrack.noise_lfsr[9] ;
 wire \vgademo.soundtrack.pulse_osc_p[0] ;
 wire \vgademo.soundtrack.pulse_osc_p[10] ;
 wire \vgademo.soundtrack.pulse_osc_p[11] ;
 wire \vgademo.soundtrack.pulse_osc_p[12] ;
 wire \vgademo.soundtrack.pulse_osc_p[13] ;
 wire \vgademo.soundtrack.pulse_osc_p[1] ;
 wire \vgademo.soundtrack.pulse_osc_p[2] ;
 wire \vgademo.soundtrack.pulse_osc_p[3] ;
 wire \vgademo.soundtrack.pulse_osc_p[4] ;
 wire \vgademo.soundtrack.pulse_osc_p[5] ;
 wire \vgademo.soundtrack.pulse_osc_p[6] ;
 wire \vgademo.soundtrack.pulse_osc_p[7] ;
 wire \vgademo.soundtrack.pulse_osc_p[8] ;
 wire \vgademo.soundtrack.pulse_osc_p[9] ;
 wire \vgademo.soundtrack.pulse_vol[0] ;
 wire \vgademo.soundtrack.pulse_vol[1] ;
 wire \vgademo.soundtrack.pulse_vol[2] ;
 wire \vgademo.soundtrack.pulse_vol[3] ;
 wire \vgademo.soundtrack.sample_div[0] ;
 wire \vgademo.soundtrack.sample_div[1] ;
 wire \vgademo.soundtrack.sample_div[2] ;
 wire \vgademo.soundtrack.sample_div[3] ;
 wire \vgademo.soundtrack.sample_div[4] ;
 wire \vgademo.soundtrack.sample_div[5] ;
 wire \vgademo.soundtrack.sample_div[6] ;
 wire \vgademo.soundtrack.sample_div[7] ;
 wire \vgademo.soundtrack.sample_div[8] ;
 wire \vgademo.soundtrack.sample_div[9] ;
 wire \vgademo.soundtrack.sample_div_[0] ;
 wire \vgademo.soundtrack.sample_div_[1] ;
 wire \vgademo.soundtrack.sample_div_[2] ;
 wire \vgademo.soundtrack.sample_div_[3] ;
 wire \vgademo.soundtrack.sample_div_[4] ;
 wire \vgademo.soundtrack.sample_div_[5] ;
 wire \vgademo.soundtrack.sample_div_[6] ;
 wire \vgademo.soundtrack.sample_div_[7] ;
 wire \vgademo.soundtrack.sample_div_[8] ;
 wire \vgademo.soundtrack.sample_div_[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[9] ;
 wire \vgademo.soundtrack.tick_div[0] ;
 wire \vgademo.soundtrack.tick_div[1] ;
 wire \vgademo.soundtrack.tick_div[2] ;
 wire \vgademo.soundtrack.tick_div[3] ;
 wire \vgademo.soundtrack.tick_div[4] ;
 wire \vgademo.soundtrack.tick_div[5] ;
 wire \vgademo.soundtrack.tick_div[6] ;
 wire \vgademo.soundtrack.tick_div[7] ;
 wire \vgademo.soundtrack.tick_div_[0] ;
 wire \vgademo.soundtrack.tri_osc_i[0] ;
 wire \vgademo.soundtrack.tri_osc_i[1] ;
 wire \vgademo.soundtrack.tri_osc_i[2] ;
 wire \vgademo.soundtrack.tri_osc_i[3] ;
 wire \vgademo.soundtrack.tri_osc_i[4] ;
 wire \vgademo.soundtrack.tri_osc_i[5] ;
 wire \vgademo.soundtrack.tri_osc_i[6] ;
 wire \vgademo.soundtrack.tri_osc_i[7] ;
 wire \vgademo.soundtrack.tri_osc_i[8] ;
 wire \vgademo.soundtrack.tri_osc_p[0] ;
 wire \vgademo.soundtrack.tri_osc_p[10] ;
 wire \vgademo.soundtrack.tri_osc_p[11] ;
 wire \vgademo.soundtrack.tri_osc_p[12] ;
 wire \vgademo.soundtrack.tri_osc_p[13] ;
 wire \vgademo.soundtrack.tri_osc_p[14] ;
 wire \vgademo.soundtrack.tri_osc_p[15] ;
 wire \vgademo.soundtrack.tri_osc_p[1] ;
 wire \vgademo.soundtrack.tri_osc_p[2] ;
 wire \vgademo.soundtrack.tri_osc_p[3] ;
 wire \vgademo.soundtrack.tri_osc_p[4] ;
 wire \vgademo.soundtrack.tri_osc_p[5] ;
 wire \vgademo.soundtrack.tri_osc_p[6] ;
 wire \vgademo.soundtrack.tri_osc_p[7] ;
 wire \vgademo.soundtrack.tri_osc_p[8] ;
 wire \vgademo.soundtrack.tri_osc_p[9] ;
 wire \vgademo.v_count[2] ;
 wire \vgademo.v_count[3] ;
 wire \vgademo.v_count[4] ;
 wire \vgademo.v_count[5] ;
 wire \vgademo.v_count[6] ;
 wire \vgademo.v_count[7] ;
 wire \vgademo.v_count[8] ;
 wire \vgademo.v_count[9] ;
 wire \vgademo.vsync ;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;

 sg13g2_inv_1 _3729_ (.Y(_3084_),
    .A(net220));
 sg13g2_inv_1 _3730_ (.Y(_3085_),
    .A(net192));
 sg13g2_inv_1 _3731_ (.Y(_3086_),
    .A(net245));
 sg13g2_inv_1 _3732_ (.Y(_3087_),
    .A(net258));
 sg13g2_inv_1 _3733_ (.Y(_3088_),
    .A(net199));
 sg13g2_inv_1 _3734_ (.Y(_3089_),
    .A(\vgademo.soundtrack.noise_lfsr[2] ));
 sg13g2_inv_1 _3735_ (.Y(_3090_),
    .A(\vgademo.soundtrack.noise_lfsr[1] ));
 sg13g2_inv_1 _3736_ (.Y(_3091_),
    .A(net168));
 sg13g2_inv_2 _3737_ (.Y(_3092_),
    .A(net1037));
 sg13g2_inv_1 _3738_ (.Y(_3093_),
    .A(net411));
 sg13g2_inv_1 _3739_ (.Y(_3094_),
    .A(net538));
 sg13g2_inv_1 _3740_ (.Y(_3095_),
    .A(net559));
 sg13g2_inv_1 _3741_ (.Y(_3096_),
    .A(net567));
 sg13g2_inv_1 _3742_ (.Y(_3097_),
    .A(net335));
 sg13g2_inv_2 _3743_ (.Y(_3098_),
    .A(net1062));
 sg13g2_inv_1 _3744_ (.Y(_3099_),
    .A(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_inv_1 _3745_ (.Y(_3100_),
    .A(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_inv_1 _3746_ (.Y(_3101_),
    .A(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_inv_1 _3747_ (.Y(_3102_),
    .A(\vgademo.audio_beat_out[2] ));
 sg13g2_inv_1 _3748_ (.Y(_3103_),
    .A(net1049));
 sg13g2_inv_2 _3749_ (.Y(_3104_),
    .A(net1054));
 sg13g2_inv_1 _3750_ (.Y(_3105_),
    .A(net1056));
 sg13g2_inv_1 _3751_ (.Y(_3106_),
    .A(net1048));
 sg13g2_inv_2 _3752_ (.Y(_3107_),
    .A(\vgademo.audio_songpos[6] ));
 sg13g2_inv_2 _3753_ (.Y(_3108_),
    .A(_0060_));
 sg13g2_inv_1 _3754_ (.Y(_3109_),
    .A(net979));
 sg13g2_inv_1 _3755_ (.Y(_3110_),
    .A(\vgademo.v_count[3] ));
 sg13g2_inv_1 _3756_ (.Y(_3111_),
    .A(\vgademo.v_count[2] ));
 sg13g2_inv_1 _3757_ (.Y(_3112_),
    .A(\vgademo.v_count[4] ));
 sg13g2_inv_1 _3758_ (.Y(_3113_),
    .A(net976));
 sg13g2_inv_1 _3759_ (.Y(_3114_),
    .A(net1014));
 sg13g2_inv_1 _3760_ (.Y(_3115_),
    .A(\vgademo.h_count[0] ));
 sg13g2_inv_1 _3761_ (.Y(_3116_),
    .A(net1011));
 sg13g2_inv_1 _3762_ (.Y(_3117_),
    .A(net1012));
 sg13g2_inv_1 _3763_ (.Y(_3118_),
    .A(\vgademo.h_count[5] ));
 sg13g2_inv_1 _3764_ (.Y(_3119_),
    .A(net1009));
 sg13g2_inv_2 _3765_ (.Y(_3120_),
    .A(\vgademo.h_count[7] ));
 sg13g2_inv_1 _3766_ (.Y(_3121_),
    .A(\vgademo.h_count[9] ));
 sg13g2_inv_4 _3767_ (.A(\vgademo.audio_songpos[7] ),
    .Y(_3122_));
 sg13g2_inv_2 _3768_ (.Y(_3123_),
    .A(net1003));
 sg13g2_inv_1 _3769_ (.Y(_3124_),
    .A(net983));
 sg13g2_inv_2 _3770_ (.Y(_3125_),
    .A(net986));
 sg13g2_inv_1 _3771_ (.Y(_3126_),
    .A(net987));
 sg13g2_inv_2 _3772_ (.Y(_3127_),
    .A(net990));
 sg13g2_inv_2 _3773_ (.Y(_3128_),
    .A(net992));
 sg13g2_inv_4 _3774_ (.A(net995),
    .Y(_3129_));
 sg13g2_inv_4 _3775_ (.A(net1002),
    .Y(_3130_));
 sg13g2_inv_2 _3776_ (.Y(_3131_),
    .A(_0066_));
 sg13g2_inv_1 _3777_ (.Y(_3132_),
    .A(_0064_));
 sg13g2_inv_1 _3778_ (.Y(_3133_),
    .A(_0069_));
 sg13g2_inv_1 _3779_ (.Y(_3134_),
    .A(net270));
 sg13g2_inv_1 _3780_ (.Y(_3135_),
    .A(_0018_));
 sg13g2_inv_1 _3781_ (.Y(_3136_),
    .A(_0020_));
 sg13g2_inv_1 _3782_ (.Y(_3137_),
    .A(net404));
 sg13g2_inv_1 _3783_ (.Y(_3138_),
    .A(net315));
 sg13g2_inv_1 _3784_ (.Y(_3139_),
    .A(net586));
 sg13g2_inv_1 _3785_ (.Y(_3140_),
    .A(net566));
 sg13g2_inv_1 _3786_ (.Y(_3141_),
    .A(net557));
 sg13g2_inv_1 _3787_ (.Y(_3142_),
    .A(\vgademo.soundtrack.pulse_vol[0] ));
 sg13g2_inv_1 _3788_ (.Y(_3143_),
    .A(\vgademo.soundtrack.pulse_vol[2] ));
 sg13g2_inv_2 _3789_ (.Y(_3144_),
    .A(net1018));
 sg13g2_inv_1 _3790_ (.Y(_3145_),
    .A(net1030));
 sg13g2_inv_2 _3791_ (.Y(_3146_),
    .A(net1023));
 sg13g2_inv_4 _3792_ (.A(net1026),
    .Y(_3147_));
 sg13g2_inv_1 _3793_ (.Y(_3148_),
    .A(net267));
 sg13g2_inv_1 _3794_ (.Y(_3149_),
    .A(net459));
 sg13g2_inv_1 _3795_ (.Y(_3150_),
    .A(\vgademo.b_sin[8] ));
 sg13g2_inv_1 _3796_ (.Y(_3151_),
    .A(\vgademo.b_sin[9] ));
 sg13g2_inv_1 _3797_ (.Y(_3152_),
    .A(\vgademo.b_sin[10] ));
 sg13g2_inv_1 _3798_ (.Y(_3153_),
    .A(\vgademo.a_cos[6] ));
 sg13g2_inv_2 _3799_ (.Y(_3154_),
    .A(net964));
 sg13g2_inv_1 _3800_ (.Y(_3155_),
    .A(net571));
 sg13g2_inv_1 _3801_ (.Y(_3156_),
    .A(\vgademo.b_cos[7] ));
 sg13g2_inv_1 _3802_ (.Y(_3157_),
    .A(\vgademo.b_cos[8] ));
 sg13g2_inv_4 _3803_ (.A(\vgademo.b_cos[9] ),
    .Y(_3158_));
 sg13g2_inv_1 _3804_ (.Y(_3159_),
    .A(net970));
 sg13g2_inv_1 _3805_ (.Y(_3160_),
    .A(net558));
 sg13g2_inv_1 _3806_ (.Y(_3161_),
    .A(net406));
 sg13g2_inv_1 _3807_ (.Y(_3162_),
    .A(net341));
 sg13g2_inv_1 _3808_ (.Y(_3163_),
    .A(net550));
 sg13g2_inv_1 _3809_ (.Y(_3164_),
    .A(net574));
 sg13g2_inv_1 _3810_ (.Y(_3165_),
    .A(\vgademo.a_sin[9] ));
 sg13g2_inv_1 _3811_ (.Y(_3166_),
    .A(net549));
 sg13g2_inv_1 _3812_ (.Y(_3167_),
    .A(\vgademo.a_sin[12] ));
 sg13g2_inv_2 _3813_ (.Y(_3168_),
    .A(net502));
 sg13g2_inv_1 _3814_ (.Y(_3169_),
    .A(net345));
 sg13g2_inv_1 _3815_ (.Y(_3170_),
    .A(net292));
 sg13g2_inv_1 _3816_ (.Y(_3171_),
    .A(\vgademo.plane_du[4] ));
 sg13g2_inv_1 _3817_ (.Y(_3172_),
    .A(net314));
 sg13g2_inv_2 _3818_ (.Y(_3173_),
    .A(net547));
 sg13g2_inv_1 _3819_ (.Y(_3174_),
    .A(net304));
 sg13g2_inv_1 _3820_ (.Y(_3175_),
    .A(net344));
 sg13g2_inv_1 _3821_ (.Y(_3176_),
    .A(\vgademo.plane_du[7] ));
 sg13g2_inv_1 _3822_ (.Y(_3177_),
    .A(net338));
 sg13g2_inv_1 _3823_ (.Y(_3178_),
    .A(_0025_));
 sg13g2_inv_1 _3824_ (.Y(_3179_),
    .A(net353));
 sg13g2_inv_1 _3825_ (.Y(_3180_),
    .A(net409));
 sg13g2_inv_1 _3826_ (.Y(_3181_),
    .A(net278));
 sg13g2_inv_1 _3827_ (.Y(_3182_),
    .A(net434));
 sg13g2_inv_1 _3828_ (.Y(_3183_),
    .A(\vgademo.plane_u[14] ));
 sg13g2_inv_1 _3829_ (.Y(_3184_),
    .A(net492));
 sg13g2_inv_1 _3830_ (.Y(_3185_),
    .A(net426));
 sg13g2_inv_1 _3831_ (.Y(_3186_),
    .A(net513));
 sg13g2_inv_1 _3832_ (.Y(_3187_),
    .A(net255));
 sg13g2_inv_1 _3833_ (.Y(_3188_),
    .A(net399));
 sg13g2_inv_1 _3834_ (.Y(_3189_),
    .A(net235));
 sg13g2_inv_1 _3835_ (.Y(_3190_),
    .A(net1063));
 sg13g2_inv_1 _3836_ (.Y(_3191_),
    .A(net396));
 sg13g2_inv_1 _3837_ (.Y(_3192_),
    .A(net405));
 sg13g2_inv_1 _3838_ (.Y(_3193_),
    .A(net376));
 sg13g2_inv_1 _3839_ (.Y(_3194_),
    .A(net354));
 sg13g2_inv_1 _3840_ (.Y(_3195_),
    .A(net447));
 sg13g2_inv_1 _3841_ (.Y(_3196_),
    .A(net417));
 sg13g2_inv_1 _3842_ (.Y(_3197_),
    .A(net190));
 sg13g2_inv_1 _3843_ (.Y(_3198_),
    .A(net309));
 sg13g2_inv_1 _3844_ (.Y(_3199_),
    .A(net352));
 sg13g2_inv_1 _3845_ (.Y(_3200_),
    .A(net369));
 sg13g2_inv_1 _3846_ (.Y(_3201_),
    .A(\vgademo.scanline_audio_sample[4] ));
 sg13g2_inv_1 _3847_ (.Y(_3202_),
    .A(_0050_));
 sg13g2_nand2_2 _3848_ (.Y(_3203_),
    .A(\vgademo.h_count[7] ),
    .B(\vgademo.h_count[6] ));
 sg13g2_nor3_1 _3849_ (.A(net957),
    .B(_3119_),
    .C(_3203_),
    .Y(_3204_));
 sg13g2_nand4_1 _3850_ (.B(net1009),
    .C(\vgademo.h_count[7] ),
    .A(\vgademo.h_count[5] ),
    .Y(_3205_),
    .D(net1008));
 sg13g2_nor2_1 _3851_ (.A(\vgademo.h_count[9] ),
    .B(_0061_),
    .Y(_3206_));
 sg13g2_nand2_1 _3852_ (.Y(_3207_),
    .A(net1007),
    .B(_3206_));
 sg13g2_nor3_1 _3853_ (.A(net1015),
    .B(\vgademo.h_count[0] ),
    .C(net1011),
    .Y(_3208_));
 sg13g2_and2_1 _3854_ (.A(net1012),
    .B(_3208_),
    .X(_3209_));
 sg13g2_nand2_2 _3855_ (.Y(_3210_),
    .A(net1012),
    .B(_3208_));
 sg13g2_nor3_2 _3856_ (.A(_3205_),
    .B(_3207_),
    .C(_3210_),
    .Y(_3211_));
 sg13g2_nand4_1 _3857_ (.B(_3204_),
    .C(_3206_),
    .A(net1007),
    .Y(_3212_),
    .D(_3209_));
 sg13g2_nor3_2 _3858_ (.A(_3205_),
    .B(_3207_),
    .C(_3210_),
    .Y(_3213_));
 sg13g2_nor2_1 _3859_ (.A(net546),
    .B(_3211_),
    .Y(_0000_));
 sg13g2_nand2_1 _3860_ (.Y(_3214_),
    .A(net1015),
    .B(\vgademo.h_count[0] ));
 sg13g2_inv_1 _3861_ (.Y(_3215_),
    .A(_3214_));
 sg13g2_xor2_1 _3862_ (.B(net546),
    .A(net1014),
    .X(_0002_));
 sg13g2_nor2_1 _3863_ (.A(net506),
    .B(_3214_),
    .Y(_3216_));
 sg13g2_and2_1 _3864_ (.A(net506),
    .B(_3214_),
    .X(_3217_));
 sg13g2_nor3_1 _3865_ (.A(_3211_),
    .B(_3216_),
    .C(_3217_),
    .Y(_0003_));
 sg13g2_xor2_1 _3866_ (.B(_3216_),
    .A(net329),
    .X(_3218_));
 sg13g2_nor2_1 _3867_ (.A(_3211_),
    .B(net330),
    .Y(_0004_));
 sg13g2_nor3_1 _3868_ (.A(_3116_),
    .B(_3117_),
    .C(_3214_),
    .Y(_3219_));
 sg13g2_and2_1 _3869_ (.A(net507),
    .B(_3219_),
    .X(_3220_));
 sg13g2_nor2_1 _3870_ (.A(net1009),
    .B(_3219_),
    .Y(_3221_));
 sg13g2_nor3_1 _3871_ (.A(_3211_),
    .B(_3220_),
    .C(_3221_),
    .Y(_0005_));
 sg13g2_xor2_1 _3872_ (.B(_3220_),
    .A(net460),
    .X(_3222_));
 sg13g2_nor2_1 _3873_ (.A(_3213_),
    .B(net461),
    .Y(_0006_));
 sg13g2_nand2_2 _3874_ (.Y(_3223_),
    .A(\vgademo.h_count[5] ),
    .B(_3220_));
 sg13g2_and2_1 _3875_ (.A(net576),
    .B(_3223_),
    .X(_3224_));
 sg13g2_nor2_1 _3876_ (.A(net576),
    .B(_3223_),
    .Y(_3225_));
 sg13g2_nor3_1 _3877_ (.A(_3211_),
    .B(net577),
    .C(_3225_),
    .Y(_0007_));
 sg13g2_xor2_1 _3878_ (.B(_3225_),
    .A(net445),
    .X(_3226_));
 sg13g2_nor2_1 _3879_ (.A(_3213_),
    .B(net446),
    .Y(_0008_));
 sg13g2_nor2_1 _3880_ (.A(_3203_),
    .B(_3223_),
    .Y(_3227_));
 sg13g2_nor2b_1 _3881_ (.A(_3227_),
    .B_N(net580),
    .Y(_3228_));
 sg13g2_nor3_2 _3882_ (.A(net580),
    .B(_3203_),
    .C(_3223_),
    .Y(_3229_));
 sg13g2_nor3_1 _3883_ (.A(_3213_),
    .B(net581),
    .C(_3229_),
    .Y(_0009_));
 sg13g2_o21ai_1 _3884_ (.B1(_3212_),
    .Y(_3230_),
    .A1(_3189_),
    .A2(_3229_));
 sg13g2_a21oi_1 _3885_ (.A1(_3189_),
    .A2(_3229_),
    .Y(_0010_),
    .B1(_3230_));
 sg13g2_nand3_1 _3886_ (.B(net1007),
    .C(_3227_),
    .A(net591),
    .Y(_3231_));
 sg13g2_a21oi_1 _3887_ (.A1(net1006),
    .A2(_3231_),
    .Y(_3232_),
    .B1(_3213_));
 sg13g2_o21ai_1 _3888_ (.B1(_3232_),
    .Y(_3233_),
    .A1(net1006),
    .A2(_3231_));
 sg13g2_inv_1 _3889_ (.Y(_0001_),
    .A(net592));
 sg13g2_nand2_2 _3890_ (.Y(_3234_),
    .A(net287),
    .B(\vgademo.v_count[6] ));
 sg13g2_nor2_1 _3891_ (.A(_0063_),
    .B(_3234_),
    .Y(_3235_));
 sg13g2_nand2_2 _3892_ (.Y(_3236_),
    .A(\vgademo.v_count[3] ),
    .B(\vgademo.v_count[2] ));
 sg13g2_nor2_2 _3893_ (.A(\vgademo.bayer_j[1] ),
    .B(net979),
    .Y(_3237_));
 sg13g2_o21ai_1 _3894_ (.B1(_3235_),
    .Y(_3238_),
    .A1(_3236_),
    .A2(_3237_));
 sg13g2_or3_1 _3895_ (.A(net979),
    .B(\vgademo.v_count[2] ),
    .C(_3235_),
    .X(_3239_));
 sg13g2_nor3_1 _3896_ (.A(net978),
    .B(_3113_),
    .C(_3234_),
    .Y(_3240_));
 sg13g2_nor2b_2 _3897_ (.A(\vgademo.v_count[9] ),
    .B_N(\vgademo.v_count[8] ),
    .Y(_3241_));
 sg13g2_nand4_1 _3898_ (.B(net473),
    .C(_3240_),
    .A(\vgademo.bayer_j[1] ),
    .Y(_3242_),
    .D(_3241_));
 sg13g2_a21o_1 _3899_ (.A2(_3239_),
    .A1(_3238_),
    .B1(_3242_),
    .X(_0012_));
 sg13g2_nor2_1 _3900_ (.A(net1014),
    .B(net1012),
    .Y(_3243_));
 sg13g2_nor3_1 _3901_ (.A(_3116_),
    .B(_3119_),
    .C(_3243_),
    .Y(_3244_));
 sg13g2_nor3_1 _3902_ (.A(\vgademo.h_count[5] ),
    .B(net1008),
    .C(_3244_),
    .Y(_3245_));
 sg13g2_o21ai_1 _3903_ (.B1(\vgademo.h_count[10] ),
    .Y(_3246_),
    .A1(_3120_),
    .A2(_3245_));
 sg13g2_o21ai_1 _3904_ (.B1(\vgademo.h_count[10] ),
    .Y(_3247_),
    .A1(net593),
    .A2(_3204_));
 sg13g2_nor3_1 _3905_ (.A(net1011),
    .B(net1013),
    .C(_0061_),
    .Y(_3248_));
 sg13g2_nor3_1 _3906_ (.A(net1011),
    .B(net1013),
    .C(_3215_),
    .Y(_3249_));
 sg13g2_nor4_1 _3907_ (.A(_3118_),
    .B(net1009),
    .C(_3203_),
    .D(_3249_),
    .Y(_3250_));
 sg13g2_o21ai_1 _3908_ (.B1(_3250_),
    .Y(_3251_),
    .A1(\vgademo.h_count[10] ),
    .A2(_3248_));
 sg13g2_a22oi_1 _3909_ (.Y(_3252_),
    .B1(_3247_),
    .B2(_3251_),
    .A2(_3246_),
    .A1(net1007));
 sg13g2_nand2_2 _3910_ (.Y(_0011_),
    .A(_3121_),
    .B(_3252_));
 sg13g2_nor2b_2 _3911_ (.A(net1056),
    .B_N(net1058),
    .Y(_3253_));
 sg13g2_nand2_1 _3912_ (.Y(_3254_),
    .A(net1058),
    .B(net959));
 sg13g2_nand2_1 _3913_ (.Y(_3255_),
    .A(net1052),
    .B(_3253_));
 sg13g2_nor2b_1 _3914_ (.A(net1061),
    .B_N(net1059),
    .Y(_3256_));
 sg13g2_nand2b_1 _3915_ (.Y(_3257_),
    .B(net1062),
    .A_N(net1060));
 sg13g2_nor2_2 _3916_ (.A(net1062),
    .B(net1056),
    .Y(_3258_));
 sg13g2_nor2b_2 _3917_ (.A(net1054),
    .B_N(net1060),
    .Y(_3259_));
 sg13g2_nor2_1 _3918_ (.A(_3258_),
    .B(_3259_),
    .Y(_3260_));
 sg13g2_nand2_1 _3919_ (.Y(_3261_),
    .A(_3257_),
    .B(_3260_));
 sg13g2_nor2_2 _3920_ (.A(net1052),
    .B(net1055),
    .Y(_3262_));
 sg13g2_nand2_2 _3921_ (.Y(_3263_),
    .A(_3104_),
    .B(net959));
 sg13g2_nor2_1 _3922_ (.A(net1049),
    .B(_3262_),
    .Y(_3264_));
 sg13g2_nand3b_1 _3923_ (.B(net1059),
    .C(net1055),
    .Y(_3265_),
    .A_N(net1061));
 sg13g2_and2_1 _3924_ (.A(net1053),
    .B(_3265_),
    .X(_3266_));
 sg13g2_xnor2_1 _3925_ (.Y(_3267_),
    .A(net1061),
    .B(net1060));
 sg13g2_nor2_2 _3926_ (.A(net1062),
    .B(net1059),
    .Y(_3268_));
 sg13g2_or2_1 _3927_ (.X(_3269_),
    .B(net1059),
    .A(net1061));
 sg13g2_and2_1 _3928_ (.A(net1061),
    .B(\vgademo.audio_songpos[1] ),
    .X(_3270_));
 sg13g2_nand2_2 _3929_ (.Y(_3271_),
    .A(net1062),
    .B(net1058));
 sg13g2_nor2_1 _3930_ (.A(_3098_),
    .B(_3105_),
    .Y(_3272_));
 sg13g2_a21oi_2 _3931_ (.B1(net1052),
    .Y(_3273_),
    .A2(net1059),
    .A1(net1061));
 sg13g2_or2_1 _3932_ (.X(_3274_),
    .B(_3273_),
    .A(_3262_));
 sg13g2_a21oi_2 _3933_ (.B1(_3262_),
    .Y(_3275_),
    .A2(_3273_),
    .A1(_3269_));
 sg13g2_a221oi_1 _3934_ (.B2(_3273_),
    .C1(_3262_),
    .B1(_3269_),
    .A1(net1053),
    .Y(_3276_),
    .A2(_3265_));
 sg13g2_nor2_1 _3935_ (.A(net1055),
    .B(_3256_),
    .Y(_3277_));
 sg13g2_nand2_2 _3936_ (.Y(_3278_),
    .A(_3105_),
    .B(_3267_));
 sg13g2_nand2_1 _3937_ (.Y(_3279_),
    .A(_3266_),
    .B(_3278_));
 sg13g2_o21ai_1 _3938_ (.B1(_3279_),
    .Y(_3280_),
    .A1(\vgademo.audio_songpos[3] ),
    .A2(_3278_));
 sg13g2_nor3_1 _3939_ (.A(net1050),
    .B(net1046),
    .C(_3262_),
    .Y(_3281_));
 sg13g2_nor2_1 _3940_ (.A(net960),
    .B(net1047),
    .Y(_3282_));
 sg13g2_nand2_2 _3941_ (.Y(_3283_),
    .A(net1050),
    .B(net958));
 sg13g2_mux2_1 _3942_ (.A0(net1061),
    .A1(_3256_),
    .S(_3255_),
    .X(_3284_));
 sg13g2_a221oi_1 _3943_ (.B2(_3284_),
    .C1(_3122_),
    .B1(_3282_),
    .A1(_3261_),
    .Y(_3285_),
    .A2(_3281_));
 sg13g2_o21ai_1 _3944_ (.B1(net960),
    .Y(_3286_),
    .A1(_3276_),
    .A2(_3277_));
 sg13g2_a221oi_1 _3945_ (.B2(_3266_),
    .C1(net960),
    .B1(_3278_),
    .A1(_3262_),
    .Y(_3287_),
    .A2(_3267_));
 sg13g2_nand3b_1 _3946_ (.B(net1047),
    .C(_3286_),
    .Y(_3288_),
    .A_N(_3287_));
 sg13g2_nor3_1 _3947_ (.A(net958),
    .B(_3264_),
    .C(_3268_),
    .Y(_3289_));
 sg13g2_nor2_2 _3948_ (.A(net1051),
    .B(net1047),
    .Y(_3290_));
 sg13g2_nand2_2 _3949_ (.Y(_3291_),
    .A(net1054),
    .B(net1056));
 sg13g2_o21ai_1 _3950_ (.B1(net1052),
    .Y(_3292_),
    .A1(net1059),
    .A2(net1055));
 sg13g2_inv_1 _3951_ (.Y(_3293_),
    .A(_3292_));
 sg13g2_nand2_1 _3952_ (.Y(_3294_),
    .A(net954),
    .B(_3292_));
 sg13g2_nand2b_2 _3953_ (.Y(_3295_),
    .B(net1052),
    .A_N(net1059));
 sg13g2_nand2b_2 _3954_ (.Y(_3296_),
    .B(net959),
    .A_N(_3295_));
 sg13g2_nand2_1 _3955_ (.Y(_3297_),
    .A(net1062),
    .B(net959));
 sg13g2_nor3_1 _3956_ (.A(_3098_),
    .B(_3283_),
    .C(_3296_),
    .Y(_3298_));
 sg13g2_nor3_1 _3957_ (.A(net1045),
    .B(_3289_),
    .C(_3298_),
    .Y(_3299_));
 sg13g2_a221oi_1 _3958_ (.B2(_3299_),
    .C1(_3107_),
    .B1(_3294_),
    .A1(_3285_),
    .Y(_3300_),
    .A2(_3288_));
 sg13g2_mux2_2 _3959_ (.A0(\vgademo.soundtrack.pulse_osc_p[13] ),
    .A1(\vgademo.soundtrack.pulse_osc_p[12] ),
    .S(_3300_),
    .X(_3301_));
 sg13g2_nand2b_1 _3960_ (.Y(_3302_),
    .B(\vgademo.soundtrack.pulse_vol[0] ),
    .A_N(_3301_));
 sg13g2_inv_1 _3961_ (.Y(_3303_),
    .A(_3302_));
 sg13g2_nor2_1 _3962_ (.A(net1020),
    .B(_3143_),
    .Y(_3304_));
 sg13g2_o21ai_1 _3963_ (.B1(_3304_),
    .Y(_3305_),
    .A1(_3142_),
    .A2(_3301_));
 sg13g2_nor2_2 _3964_ (.A(_3144_),
    .B(_3305_),
    .Y(_3306_));
 sg13g2_nor2_1 _3965_ (.A(net1034),
    .B(_0040_),
    .Y(_3307_));
 sg13g2_a21oi_1 _3966_ (.A1(net1034),
    .A2(\vgademo.soundtrack.noise_lfsr[5] ),
    .Y(_3308_),
    .B1(_3307_));
 sg13g2_mux2_1 _3967_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(\vgademo.soundtrack.noise_lfsr[7] ),
    .S(net1034),
    .X(_3309_));
 sg13g2_nand2_1 _3968_ (.Y(_3310_),
    .A(net1030),
    .B(_3309_));
 sg13g2_o21ai_1 _3969_ (.B1(_3310_),
    .Y(_3311_),
    .A1(net1029),
    .A2(_3308_));
 sg13g2_nor2_1 _3970_ (.A(_3089_),
    .B(net1033),
    .Y(_3312_));
 sg13g2_a21oi_1 _3971_ (.A1(\vgademo.soundtrack.noise_lfsr[3] ),
    .A2(net1033),
    .Y(_3313_),
    .B1(_3312_));
 sg13g2_a21oi_1 _3972_ (.A1(_3090_),
    .A2(net1033),
    .Y(_3314_),
    .B1(net1030));
 sg13g2_o21ai_1 _3973_ (.B1(_3314_),
    .Y(_3315_),
    .A1(net1033),
    .A2(\vgademo.soundtrack.noise_lfsr[0] ));
 sg13g2_o21ai_1 _3974_ (.B1(_3315_),
    .Y(_3316_),
    .A1(_3145_),
    .A2(_3313_));
 sg13g2_mux2_1 _3975_ (.A0(\vgademo.soundtrack.noise_lfsr[10] ),
    .A1(\vgademo.soundtrack.noise_lfsr[11] ),
    .S(net1032),
    .X(_3317_));
 sg13g2_nand2_1 _3976_ (.Y(_3318_),
    .A(net1029),
    .B(_3317_));
 sg13g2_nand2b_1 _3977_ (.Y(_3319_),
    .B(net1032),
    .A_N(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_o21ai_1 _3978_ (.B1(_3319_),
    .Y(_3320_),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .A2(net1032));
 sg13g2_o21ai_1 _3979_ (.B1(_3318_),
    .Y(_3321_),
    .A1(net1028),
    .A2(_3320_));
 sg13g2_nand2b_1 _3980_ (.Y(_3322_),
    .B(\vgademo.soundtrack.noise_lfsr[12] ),
    .A_N(net1032));
 sg13g2_nor2_1 _3981_ (.A(net1028),
    .B(_3322_),
    .Y(_3323_));
 sg13g2_mux2_1 _3982_ (.A0(_3321_),
    .A1(_3323_),
    .S(net1024),
    .X(_3324_));
 sg13g2_nand2_1 _3983_ (.Y(_3325_),
    .A(net1022),
    .B(_3324_));
 sg13g2_nor2_1 _3984_ (.A(net1025),
    .B(_3316_),
    .Y(_3326_));
 sg13g2_o21ai_1 _3985_ (.B1(_3146_),
    .Y(_3327_),
    .A1(_3147_),
    .A2(_3311_));
 sg13g2_o21ai_1 _3986_ (.B1(_3325_),
    .Y(_3328_),
    .A1(_3326_),
    .A2(_3327_));
 sg13g2_nand2_1 _3987_ (.Y(_3329_),
    .A(_3306_),
    .B(_3328_));
 sg13g2_xnor2_1 _3988_ (.Y(_3330_),
    .A(_3306_),
    .B(_3328_));
 sg13g2_xnor2_1 _3989_ (.Y(_3331_),
    .A(net1017),
    .B(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_xor2_1 _3990_ (.B(_3331_),
    .A(_3330_),
    .X(_3332_));
 sg13g2_nand2_1 _3991_ (.Y(_3333_),
    .A(net214),
    .B(_3332_));
 sg13g2_xor2_1 _3992_ (.B(_3332_),
    .A(net214),
    .X(\vgademo.soundtrack.sigma_delta_accum_[0] ));
 sg13g2_and2_1 _3993_ (.A(net1020),
    .B(\vgademo.soundtrack.pulse_vol[2] ),
    .X(_3334_));
 sg13g2_nand2_2 _3994_ (.Y(_3335_),
    .A(net1020),
    .B(\vgademo.soundtrack.pulse_vol[2] ));
 sg13g2_nor2_1 _3995_ (.A(_3144_),
    .B(_3335_),
    .Y(_3336_));
 sg13g2_xnor2_1 _3996_ (.Y(_3337_),
    .A(net1019),
    .B(_3334_));
 sg13g2_nor2_1 _3997_ (.A(net1020),
    .B(\vgademo.soundtrack.pulse_vol[2] ),
    .Y(_3338_));
 sg13g2_inv_1 _3998_ (.Y(_3339_),
    .A(_3338_));
 sg13g2_and2_1 _3999_ (.A(net1020),
    .B(\vgademo.soundtrack.pulse_vol[0] ),
    .X(_3340_));
 sg13g2_nor2_1 _4000_ (.A(net1020),
    .B(\vgademo.soundtrack.pulse_vol[0] ),
    .Y(_3341_));
 sg13g2_nor2_1 _4001_ (.A(_3340_),
    .B(_3341_),
    .Y(_3342_));
 sg13g2_a21o_1 _4002_ (.A2(_3341_),
    .A1(_3301_),
    .B1(_3340_),
    .X(_3343_));
 sg13g2_nand4_1 _4003_ (.B(_3335_),
    .C(_3339_),
    .A(net1019),
    .Y(_3344_),
    .D(_3343_));
 sg13g2_nor2b_1 _4004_ (.A(net1034),
    .B_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Y(_3345_));
 sg13g2_a21oi_1 _4005_ (.A1(\vgademo.soundtrack.noise_lfsr[6] ),
    .A2(net1034),
    .Y(_3346_),
    .B1(_3345_));
 sg13g2_mux2_1 _4006_ (.A0(\vgademo.soundtrack.noise_lfsr[7] ),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .S(net1034),
    .X(_3347_));
 sg13g2_nand2_1 _4007_ (.Y(_3348_),
    .A(net1030),
    .B(_3347_));
 sg13g2_o21ai_1 _4008_ (.B1(_3348_),
    .Y(_3349_),
    .A1(net1029),
    .A2(_3346_));
 sg13g2_nand2b_1 _4009_ (.Y(_3350_),
    .B(net1025),
    .A_N(_3349_));
 sg13g2_nor2_1 _4010_ (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .B(net1033),
    .Y(_3351_));
 sg13g2_a21oi_1 _4011_ (.A1(net1032),
    .A2(_0040_),
    .Y(_3352_),
    .B1(_3351_));
 sg13g2_a21oi_1 _4012_ (.A1(_3089_),
    .A2(net1033),
    .Y(_3353_),
    .B1(net1030));
 sg13g2_o21ai_1 _4013_ (.B1(_3353_),
    .Y(_3354_),
    .A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(net1033));
 sg13g2_a21oi_1 _4014_ (.A1(net1031),
    .A2(_3352_),
    .Y(_3355_),
    .B1(net1025));
 sg13g2_a21oi_1 _4015_ (.A1(_3354_),
    .A2(_3355_),
    .Y(_3356_),
    .B1(net1021));
 sg13g2_nor2b_1 _4016_ (.A(net1032),
    .B_N(\vgademo.soundtrack.noise_lfsr[9] ),
    .Y(_3357_));
 sg13g2_a21oi_1 _4017_ (.A1(net1032),
    .A2(\vgademo.soundtrack.noise_lfsr[10] ),
    .Y(_3358_),
    .B1(_3357_));
 sg13g2_mux2_1 _4018_ (.A0(\vgademo.soundtrack.noise_lfsr[11] ),
    .A1(\vgademo.soundtrack.noise_lfsr[12] ),
    .S(net1032),
    .X(_3359_));
 sg13g2_nand2_1 _4019_ (.Y(_3360_),
    .A(net1028),
    .B(_3359_));
 sg13g2_o21ai_1 _4020_ (.B1(_3360_),
    .Y(_3361_),
    .A1(net1028),
    .A2(_3358_));
 sg13g2_and2_1 _4021_ (.A(_3147_),
    .B(_3361_),
    .X(_3362_));
 sg13g2_a22oi_1 _4022_ (.Y(_3363_),
    .B1(_3362_),
    .B2(net1021),
    .A2(_3356_),
    .A1(_3350_));
 sg13g2_nor2_1 _4023_ (.A(_3344_),
    .B(_3363_),
    .Y(_3364_));
 sg13g2_xor2_1 _4024_ (.B(_3363_),
    .A(_3344_),
    .X(_3365_));
 sg13g2_xor2_1 _4025_ (.B(\vgademo.soundtrack.tri_osc_p[2] ),
    .A(net1017),
    .X(_3366_));
 sg13g2_xnor2_1 _4026_ (.Y(_3367_),
    .A(_3365_),
    .B(_3366_));
 sg13g2_o21ai_1 _4027_ (.B1(_3329_),
    .Y(_3368_),
    .A1(_3330_),
    .A2(_3331_));
 sg13g2_nand2b_1 _4028_ (.Y(_3369_),
    .B(_3368_),
    .A_N(_3367_));
 sg13g2_xnor2_1 _4029_ (.Y(_3370_),
    .A(_3367_),
    .B(_3368_));
 sg13g2_nand2_1 _4030_ (.Y(_3371_),
    .A(net381),
    .B(_3370_));
 sg13g2_xnor2_1 _4031_ (.Y(_3372_),
    .A(net381),
    .B(_3370_));
 sg13g2_xor2_1 _4032_ (.B(_3372_),
    .A(_3333_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[1] ));
 sg13g2_o21ai_1 _4033_ (.B1(_3371_),
    .Y(_3373_),
    .A1(_3333_),
    .A2(_3372_));
 sg13g2_a21oi_2 _4034_ (.B1(_3364_),
    .Y(_3374_),
    .A2(_3366_),
    .A1(_3365_));
 sg13g2_nand4_1 _4035_ (.B(_3143_),
    .C(net1018),
    .A(\vgademo.soundtrack.pulse_vol[1] ),
    .Y(_3375_),
    .D(_3302_));
 sg13g2_nor2_1 _4036_ (.A(net1029),
    .B(_3309_),
    .Y(_3376_));
 sg13g2_a21oi_2 _4037_ (.B1(_3376_),
    .Y(_3377_),
    .A2(_3320_),
    .A1(net1028));
 sg13g2_mux2_1 _4038_ (.A0(_3313_),
    .A1(_3308_),
    .S(net1030),
    .X(_3378_));
 sg13g2_nor2_1 _4039_ (.A(net1024),
    .B(_3378_),
    .Y(_3379_));
 sg13g2_a21oi_1 _4040_ (.A1(net1024),
    .A2(_3377_),
    .Y(_3380_),
    .B1(_3379_));
 sg13g2_nor2_1 _4041_ (.A(net1028),
    .B(_3317_),
    .Y(_3381_));
 sg13g2_a21oi_2 _4042_ (.B1(_3381_),
    .Y(_3382_),
    .A2(_3322_),
    .A1(net1028));
 sg13g2_inv_1 _4043_ (.Y(_3383_),
    .A(_3382_));
 sg13g2_nand3_1 _4044_ (.B(_3147_),
    .C(_3382_),
    .A(net1021),
    .Y(_3384_));
 sg13g2_o21ai_1 _4045_ (.B1(_3384_),
    .Y(_3385_),
    .A1(net1021),
    .A2(_3380_));
 sg13g2_nand2b_1 _4046_ (.Y(_3386_),
    .B(_3385_),
    .A_N(_3375_));
 sg13g2_xor2_1 _4047_ (.B(_3385_),
    .A(_3375_),
    .X(_3387_));
 sg13g2_xnor2_1 _4048_ (.Y(_3388_),
    .A(net1017),
    .B(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_xnor2_1 _4049_ (.Y(_0366_),
    .A(_3387_),
    .B(_3388_));
 sg13g2_or2_1 _4050_ (.X(_0367_),
    .B(_0366_),
    .A(_3374_));
 sg13g2_and2_1 _4051_ (.A(_3374_),
    .B(_0366_),
    .X(_0368_));
 sg13g2_xor2_1 _4052_ (.B(_0366_),
    .A(_3374_),
    .X(_0369_));
 sg13g2_xnor2_1 _4053_ (.Y(_0370_),
    .A(_3369_),
    .B(_0369_));
 sg13g2_and2_1 _4054_ (.A(net570),
    .B(_0370_),
    .X(_0371_));
 sg13g2_or2_1 _4055_ (.X(_0372_),
    .B(_0370_),
    .A(net570));
 sg13g2_nand2b_1 _4056_ (.Y(_0373_),
    .B(_0372_),
    .A_N(_0371_));
 sg13g2_xnor2_1 _4057_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .A(_3373_),
    .B(_0373_));
 sg13g2_a21oi_1 _4058_ (.A1(_3373_),
    .A2(_0372_),
    .Y(_0374_),
    .B1(_0371_));
 sg13g2_o21ai_1 _4059_ (.B1(_0367_),
    .Y(_0375_),
    .A1(_3369_),
    .A2(_0368_));
 sg13g2_o21ai_1 _4060_ (.B1(_3386_),
    .Y(_0376_),
    .A1(_3387_),
    .A2(_3388_));
 sg13g2_nor3_1 _4061_ (.A(\vgademo.soundtrack.pulse_vol[2] ),
    .B(_3340_),
    .C(_3341_),
    .Y(_0377_));
 sg13g2_o21ai_1 _4062_ (.B1(_0377_),
    .Y(_0378_),
    .A1(\vgademo.soundtrack.pulse_vol[0] ),
    .A2(_3301_));
 sg13g2_nor2_2 _4063_ (.A(_3337_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_nor2_1 _4064_ (.A(net1030),
    .B(_3347_),
    .Y(_0380_));
 sg13g2_a21oi_1 _4065_ (.A1(net1029),
    .A2(_3358_),
    .Y(_0381_),
    .B1(_0380_));
 sg13g2_or2_1 _4066_ (.X(_0382_),
    .B(_3352_),
    .A(net1029));
 sg13g2_a21oi_1 _4067_ (.A1(net1029),
    .A2(_3346_),
    .Y(_0383_),
    .B1(net1024));
 sg13g2_a221oi_1 _4068_ (.B2(_0383_),
    .C1(net1021),
    .B1(_0382_),
    .A1(net1024),
    .Y(_0384_),
    .A2(_0381_));
 sg13g2_nand2b_1 _4069_ (.Y(_0385_),
    .B(_3359_),
    .A_N(net1028));
 sg13g2_nand2b_1 _4070_ (.Y(_0386_),
    .B(_3147_),
    .A_N(_0385_));
 sg13g2_a21o_1 _4071_ (.A2(_0386_),
    .A1(net1021),
    .B1(_0384_),
    .X(_0387_));
 sg13g2_inv_1 _4072_ (.Y(_0388_),
    .A(_0387_));
 sg13g2_xnor2_1 _4073_ (.Y(_0389_),
    .A(_0379_),
    .B(_0388_));
 sg13g2_xor2_1 _4074_ (.B(\vgademo.soundtrack.tri_osc_p[4] ),
    .A(net1017),
    .X(_0390_));
 sg13g2_nor2b_1 _4075_ (.A(_0389_),
    .B_N(_0390_),
    .Y(_0391_));
 sg13g2_xnor2_1 _4076_ (.Y(_0392_),
    .A(_0389_),
    .B(_0390_));
 sg13g2_and2_1 _4077_ (.A(_0376_),
    .B(_0392_),
    .X(_0393_));
 sg13g2_or2_1 _4078_ (.X(_0394_),
    .B(_0392_),
    .A(_0376_));
 sg13g2_nand2b_1 _4079_ (.Y(_0395_),
    .B(_0394_),
    .A_N(_0393_));
 sg13g2_xnor2_1 _4080_ (.Y(_0396_),
    .A(_0375_),
    .B(_0395_));
 sg13g2_nand2_1 _4081_ (.Y(_0397_),
    .A(net536),
    .B(_0396_));
 sg13g2_xnor2_1 _4082_ (.Y(_0398_),
    .A(net536),
    .B(_0396_));
 sg13g2_xor2_1 _4083_ (.B(_0398_),
    .A(_0374_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[3] ));
 sg13g2_o21ai_1 _4084_ (.B1(_0397_),
    .Y(_0399_),
    .A1(_0374_),
    .A2(_0398_));
 sg13g2_a21o_1 _4085_ (.A2(_0394_),
    .A1(_0375_),
    .B1(_0393_),
    .X(_0400_));
 sg13g2_a21oi_1 _4086_ (.A1(_0379_),
    .A2(_0388_),
    .Y(_0401_),
    .B1(_0391_));
 sg13g2_nand3_1 _4087_ (.B(_3302_),
    .C(_3338_),
    .A(net1018),
    .Y(_0402_));
 sg13g2_nand2_1 _4088_ (.Y(_0403_),
    .A(_3147_),
    .B(_3323_));
 sg13g2_nand2_1 _4089_ (.Y(_0404_),
    .A(net1024),
    .B(_3321_));
 sg13g2_a21oi_1 _4090_ (.A1(_3147_),
    .A2(_3311_),
    .Y(_0405_),
    .B1(net1022));
 sg13g2_a22oi_1 _4091_ (.Y(_0406_),
    .B1(_0404_),
    .B2(_0405_),
    .A2(_0403_),
    .A1(net1021));
 sg13g2_nand2b_1 _4092_ (.Y(_0407_),
    .B(_0406_),
    .A_N(_0402_));
 sg13g2_xnor2_1 _4093_ (.Y(_0408_),
    .A(_0402_),
    .B(_0406_));
 sg13g2_inv_1 _4094_ (.Y(_0409_),
    .A(_0408_));
 sg13g2_xnor2_1 _4095_ (.Y(_0410_),
    .A(net1017),
    .B(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_xor2_1 _4096_ (.B(_0410_),
    .A(_0408_),
    .X(_0411_));
 sg13g2_nor2_1 _4097_ (.A(_0401_),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_xor2_1 _4098_ (.B(_0411_),
    .A(_0401_),
    .X(_0413_));
 sg13g2_xor2_1 _4099_ (.B(_0413_),
    .A(_0400_),
    .X(_0414_));
 sg13g2_and2_1 _4100_ (.A(net579),
    .B(_0414_),
    .X(_0415_));
 sg13g2_or2_1 _4101_ (.X(_0416_),
    .B(_0414_),
    .A(net579));
 sg13g2_nand2b_1 _4102_ (.Y(_0417_),
    .B(_0416_),
    .A_N(_0415_));
 sg13g2_xnor2_1 _4103_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .A(_0399_),
    .B(_0417_));
 sg13g2_a21oi_1 _4104_ (.A1(_0399_),
    .A2(_0416_),
    .Y(_0418_),
    .B1(_0415_));
 sg13g2_a21oi_1 _4105_ (.A1(_0400_),
    .A2(_0413_),
    .Y(_0419_),
    .B1(_0412_));
 sg13g2_o21ai_1 _4106_ (.B1(_0407_),
    .Y(_0420_),
    .A1(_0409_),
    .A2(_0410_));
 sg13g2_nor2_1 _4107_ (.A(net1024),
    .B(_3349_),
    .Y(_0421_));
 sg13g2_nor2_1 _4108_ (.A(net1022),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_o21ai_1 _4109_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_3147_),
    .A2(_3361_));
 sg13g2_o21ai_1 _4110_ (.B1(_3343_),
    .Y(_0424_),
    .A1(_3334_),
    .A2(_3338_));
 sg13g2_or2_1 _4111_ (.X(_0425_),
    .B(_0424_),
    .A(_3337_));
 sg13g2_xor2_1 _4112_ (.B(_0425_),
    .A(_0423_),
    .X(_0426_));
 sg13g2_xnor2_1 _4113_ (.Y(_0427_),
    .A(net1017),
    .B(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_nand2b_1 _4114_ (.Y(_0428_),
    .B(_0426_),
    .A_N(_0427_));
 sg13g2_xnor2_1 _4115_ (.Y(_0429_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_nand2_1 _4116_ (.Y(_0430_),
    .A(_0420_),
    .B(_0429_));
 sg13g2_xnor2_1 _4117_ (.Y(_0431_),
    .A(_0420_),
    .B(_0429_));
 sg13g2_xor2_1 _4118_ (.B(_0431_),
    .A(_0419_),
    .X(_0432_));
 sg13g2_nand2_1 _4119_ (.Y(_0433_),
    .A(net532),
    .B(_0432_));
 sg13g2_xnor2_1 _4120_ (.Y(_0434_),
    .A(net532),
    .B(_0432_));
 sg13g2_xor2_1 _4121_ (.B(_0434_),
    .A(_0418_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[5] ));
 sg13g2_o21ai_1 _4122_ (.B1(_0433_),
    .Y(_0435_),
    .A1(_0418_),
    .A2(_0434_));
 sg13g2_o21ai_1 _4123_ (.B1(_0430_),
    .Y(_0436_),
    .A1(_0419_),
    .A2(_0431_));
 sg13g2_o21ai_1 _4124_ (.B1(_0428_),
    .Y(_0437_),
    .A1(_0423_),
    .A2(_0425_));
 sg13g2_a21oi_1 _4125_ (.A1(net1027),
    .A2(_3383_),
    .Y(_0438_),
    .B1(net1023));
 sg13g2_o21ai_1 _4126_ (.B1(_0438_),
    .Y(_0439_),
    .A1(net1027),
    .A2(_3377_));
 sg13g2_nor3_1 _4127_ (.A(net1018),
    .B(_3303_),
    .C(_3335_),
    .Y(_0440_));
 sg13g2_nor2b_1 _4128_ (.A(_0439_),
    .B_N(_0440_),
    .Y(_0441_));
 sg13g2_xnor2_1 _4129_ (.Y(_0442_),
    .A(_0439_),
    .B(_0440_));
 sg13g2_xnor2_1 _4130_ (.Y(_0443_),
    .A(net1017),
    .B(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_inv_1 _4131_ (.Y(_0444_),
    .A(_0443_));
 sg13g2_xnor2_1 _4132_ (.Y(_0445_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_and2_1 _4133_ (.A(_0437_),
    .B(_0445_),
    .X(_0446_));
 sg13g2_xnor2_1 _4134_ (.Y(_0447_),
    .A(_0437_),
    .B(_0445_));
 sg13g2_inv_1 _4135_ (.Y(_0448_),
    .A(_0447_));
 sg13g2_xnor2_1 _4136_ (.Y(_0449_),
    .A(_0436_),
    .B(_0447_));
 sg13g2_and2_1 _4137_ (.A(net565),
    .B(_0449_),
    .X(_0450_));
 sg13g2_or2_1 _4138_ (.X(_0451_),
    .B(_0449_),
    .A(net565));
 sg13g2_nand2b_1 _4139_ (.Y(_0452_),
    .B(_0451_),
    .A_N(_0450_));
 sg13g2_xnor2_1 _4140_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[6] ),
    .A(_0435_),
    .B(_0452_));
 sg13g2_a21oi_1 _4141_ (.A1(_0435_),
    .A2(_0451_),
    .Y(_0453_),
    .B1(_0450_));
 sg13g2_a21oi_1 _4142_ (.A1(_0436_),
    .A2(_0448_),
    .Y(_0454_),
    .B1(_0446_));
 sg13g2_a21oi_1 _4143_ (.A1(_0442_),
    .A2(_0444_),
    .Y(_0455_),
    .B1(_0441_));
 sg13g2_o21ai_1 _4144_ (.B1(_3146_),
    .Y(_0456_),
    .A1(net1025),
    .A2(_0381_));
 sg13g2_a21oi_2 _4145_ (.B1(_0456_),
    .Y(_0457_),
    .A2(_0385_),
    .A1(net1024));
 sg13g2_nor3_1 _4146_ (.A(net1020),
    .B(_3142_),
    .C(_3143_),
    .Y(_0458_));
 sg13g2_nor3_1 _4147_ (.A(\vgademo.soundtrack.pulse_vol[0] ),
    .B(net1018),
    .C(_3335_),
    .Y(_0459_));
 sg13g2_a22oi_1 _4148_ (.Y(_0460_),
    .B1(_0459_),
    .B2(_3301_),
    .A2(_0458_),
    .A1(_3144_));
 sg13g2_nor2b_1 _4149_ (.A(_0460_),
    .B_N(_0457_),
    .Y(_0461_));
 sg13g2_xnor2_1 _4150_ (.Y(_0462_),
    .A(_0457_),
    .B(_0460_));
 sg13g2_xnor2_1 _4151_ (.Y(_0463_),
    .A(net1017),
    .B(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_inv_1 _4152_ (.Y(_0464_),
    .A(_0463_));
 sg13g2_xnor2_1 _4153_ (.Y(_0465_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_nand2b_1 _4154_ (.Y(_0466_),
    .B(_0465_),
    .A_N(_0455_));
 sg13g2_xnor2_1 _4155_ (.Y(_0467_),
    .A(_0455_),
    .B(_0465_));
 sg13g2_nand2b_1 _4156_ (.Y(_0468_),
    .B(_0467_),
    .A_N(_0454_));
 sg13g2_xnor2_1 _4157_ (.Y(_0469_),
    .A(_0454_),
    .B(_0467_));
 sg13g2_nand2_1 _4158_ (.Y(_0470_),
    .A(\vgademo.soundtrack.sigma_delta_accum[7] ),
    .B(_0469_));
 sg13g2_xnor2_1 _4159_ (.Y(_0471_),
    .A(net527),
    .B(_0469_));
 sg13g2_xor2_1 _4160_ (.B(_0471_),
    .A(_0453_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[7] ));
 sg13g2_o21ai_1 _4161_ (.B1(_0470_),
    .Y(_0472_),
    .A1(_0453_),
    .A2(_0471_));
 sg13g2_nand2_1 _4162_ (.Y(_0473_),
    .A(_0466_),
    .B(_0468_));
 sg13g2_a21oi_1 _4163_ (.A1(_0462_),
    .A2(_0464_),
    .Y(_0474_),
    .B1(_0461_));
 sg13g2_and2_1 _4164_ (.A(_3146_),
    .B(_3324_),
    .X(_0475_));
 sg13g2_nor2_1 _4165_ (.A(net1018),
    .B(_3305_),
    .Y(_0476_));
 sg13g2_nand2_1 _4166_ (.Y(_0477_),
    .A(_0475_),
    .B(_0476_));
 sg13g2_xnor2_1 _4167_ (.Y(_0478_),
    .A(_0475_),
    .B(_0476_));
 sg13g2_xnor2_1 _4168_ (.Y(_0479_),
    .A(net1016),
    .B(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_xnor2_1 _4169_ (.Y(_0480_),
    .A(_0478_),
    .B(_0479_));
 sg13g2_xor2_1 _4170_ (.B(_0480_),
    .A(_0474_),
    .X(_0481_));
 sg13g2_nand2_1 _4171_ (.Y(_0482_),
    .A(_0473_),
    .B(_0481_));
 sg13g2_xor2_1 _4172_ (.B(_0481_),
    .A(_0473_),
    .X(_0483_));
 sg13g2_xnor2_1 _4173_ (.Y(_0484_),
    .A(net516),
    .B(_0483_));
 sg13g2_nor2b_1 _4174_ (.A(_0484_),
    .B_N(_0472_),
    .Y(_0485_));
 sg13g2_xnor2_1 _4175_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[8] ),
    .A(_0472_),
    .B(_0484_));
 sg13g2_a21o_1 _4176_ (.A2(_0483_),
    .A1(net516),
    .B1(_0485_),
    .X(_0486_));
 sg13g2_o21ai_1 _4177_ (.B1(_0482_),
    .Y(_0487_),
    .A1(_0474_),
    .A2(_0480_));
 sg13g2_o21ai_1 _4178_ (.B1(_0477_),
    .Y(_0488_),
    .A1(_0478_),
    .A2(_0479_));
 sg13g2_nand2_1 _4179_ (.Y(_0489_),
    .A(_3146_),
    .B(_3362_));
 sg13g2_inv_1 _4180_ (.Y(_0490_),
    .A(_0489_));
 sg13g2_and4_1 _4181_ (.A(_3144_),
    .B(_3335_),
    .C(_3339_),
    .D(_3343_),
    .X(_0491_));
 sg13g2_xnor2_1 _4182_ (.Y(_0492_),
    .A(_0490_),
    .B(_0491_));
 sg13g2_xnor2_1 _4183_ (.Y(_0493_),
    .A(net1016),
    .B(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_nor2_1 _4184_ (.A(_0492_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_xor2_1 _4185_ (.B(_0493_),
    .A(_0492_),
    .X(_0495_));
 sg13g2_and2_1 _4186_ (.A(_0488_),
    .B(_0495_),
    .X(_0496_));
 sg13g2_xor2_1 _4187_ (.B(_0495_),
    .A(_0488_),
    .X(_0497_));
 sg13g2_xor2_1 _4188_ (.B(_0497_),
    .A(_0487_),
    .X(_0498_));
 sg13g2_xnor2_1 _4189_ (.Y(_0499_),
    .A(net526),
    .B(_0498_));
 sg13g2_nor2b_1 _4190_ (.A(_0499_),
    .B_N(_0486_),
    .Y(_0500_));
 sg13g2_xnor2_1 _4191_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .A(_0486_),
    .B(_0499_));
 sg13g2_a21o_1 _4192_ (.A2(_0498_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[9] ),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_a21o_1 _4193_ (.A2(_0497_),
    .A1(_0487_),
    .B1(_0496_),
    .X(_0502_));
 sg13g2_a21oi_1 _4194_ (.A1(_0490_),
    .A2(_0491_),
    .Y(_0503_),
    .B1(_0494_));
 sg13g2_nor3_2 _4195_ (.A(net1023),
    .B(net1027),
    .C(_3383_),
    .Y(_0504_));
 sg13g2_and4_1 _4196_ (.A(net1020),
    .B(_3143_),
    .C(_3144_),
    .D(_3302_),
    .X(_0505_));
 sg13g2_xnor2_1 _4197_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_xor2_1 _4198_ (.B(\vgademo.soundtrack.tri_osc_p[11] ),
    .A(net1016),
    .X(_0507_));
 sg13g2_nor2b_1 _4199_ (.A(_0506_),
    .B_N(_0507_),
    .Y(_0508_));
 sg13g2_xnor2_1 _4200_ (.Y(_0509_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_nor2b_1 _4201_ (.A(_0503_),
    .B_N(_0509_),
    .Y(_0510_));
 sg13g2_xnor2_1 _4202_ (.Y(_0511_),
    .A(_0503_),
    .B(_0509_));
 sg13g2_xor2_1 _4203_ (.B(_0511_),
    .A(_0502_),
    .X(_0512_));
 sg13g2_xnor2_1 _4204_ (.Y(_0513_),
    .A(net504),
    .B(_0512_));
 sg13g2_nor2b_1 _4205_ (.A(_0513_),
    .B_N(_0501_),
    .Y(_0514_));
 sg13g2_xnor2_1 _4206_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .A(_0501_),
    .B(_0513_));
 sg13g2_a21o_1 _4207_ (.A2(_0512_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .B1(_0514_),
    .X(_0515_));
 sg13g2_a21oi_1 _4208_ (.A1(_0502_),
    .A2(_0511_),
    .Y(_0516_),
    .B1(_0510_));
 sg13g2_a21o_1 _4209_ (.A2(_0505_),
    .A1(_0504_),
    .B1(_0508_),
    .X(_0517_));
 sg13g2_nand2b_2 _4210_ (.Y(_0518_),
    .B(_3146_),
    .A_N(_0386_));
 sg13g2_nand2b_1 _4211_ (.Y(_0519_),
    .B(_3337_),
    .A_N(_0378_));
 sg13g2_nor2_1 _4212_ (.A(_0518_),
    .B(_0519_),
    .Y(_0520_));
 sg13g2_xor2_1 _4213_ (.B(_0519_),
    .A(_0518_),
    .X(_0521_));
 sg13g2_xor2_1 _4214_ (.B(\vgademo.soundtrack.tri_osc_p[12] ),
    .A(net1016),
    .X(_0522_));
 sg13g2_xor2_1 _4215_ (.B(_0522_),
    .A(_0521_),
    .X(_0523_));
 sg13g2_nand2_1 _4216_ (.Y(_0524_),
    .A(_0517_),
    .B(_0523_));
 sg13g2_xnor2_1 _4217_ (.Y(_0525_),
    .A(_0517_),
    .B(_0523_));
 sg13g2_xor2_1 _4218_ (.B(_0525_),
    .A(_0516_),
    .X(_0526_));
 sg13g2_xnor2_1 _4219_ (.Y(_0527_),
    .A(net494),
    .B(_0526_));
 sg13g2_nor2b_1 _4220_ (.A(_0527_),
    .B_N(_0515_),
    .Y(_0528_));
 sg13g2_xnor2_1 _4221_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .A(_0515_),
    .B(_0527_));
 sg13g2_a21o_1 _4222_ (.A2(_0526_),
    .A1(net494),
    .B1(_0528_),
    .X(_0529_));
 sg13g2_o21ai_1 _4223_ (.B1(_0524_),
    .Y(_0530_),
    .A1(_0516_),
    .A2(_0525_));
 sg13g2_a21oi_1 _4224_ (.A1(_0521_),
    .A2(_0522_),
    .Y(_0531_),
    .B1(_0520_));
 sg13g2_nor2_2 _4225_ (.A(net1021),
    .B(_0403_),
    .Y(_0532_));
 sg13g2_nor3_2 _4226_ (.A(net1018),
    .B(_3303_),
    .C(_3339_),
    .Y(_0533_));
 sg13g2_and2_1 _4227_ (.A(_0532_),
    .B(_0533_),
    .X(_0534_));
 sg13g2_xnor2_1 _4228_ (.Y(_0535_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_xnor2_1 _4229_ (.Y(_0536_),
    .A(net1016),
    .B(\vgademo.soundtrack.tri_osc_p[13] ));
 sg13g2_nor2_1 _4230_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_xor2_1 _4231_ (.B(_0536_),
    .A(_0535_),
    .X(_0538_));
 sg13g2_nor2b_1 _4232_ (.A(_0531_),
    .B_N(_0538_),
    .Y(_0539_));
 sg13g2_nand2b_1 _4233_ (.Y(_0540_),
    .B(_0531_),
    .A_N(_0538_));
 sg13g2_nand2b_1 _4234_ (.Y(_0541_),
    .B(_0540_),
    .A_N(_0539_));
 sg13g2_xnor2_1 _4235_ (.Y(_0542_),
    .A(_0530_),
    .B(_0541_));
 sg13g2_xnor2_1 _4236_ (.Y(_0543_),
    .A(net512),
    .B(_0542_));
 sg13g2_nor2b_1 _4237_ (.A(_0543_),
    .B_N(_0529_),
    .Y(_0544_));
 sg13g2_xnor2_1 _4238_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .A(_0529_),
    .B(_0543_));
 sg13g2_a21o_1 _4239_ (.A2(_0542_),
    .A1(net512),
    .B1(_0544_),
    .X(_0545_));
 sg13g2_nor3_2 _4240_ (.A(net1018),
    .B(_3334_),
    .C(_0424_),
    .Y(_0546_));
 sg13g2_nand2b_1 _4241_ (.Y(_0547_),
    .B(net354),
    .A_N(net1016));
 sg13g2_xor2_1 _4242_ (.B(net1016),
    .A(\vgademo.soundtrack.tri_osc_p[14] ),
    .X(_0548_));
 sg13g2_nor2_1 _4243_ (.A(_0546_),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_xnor2_1 _4244_ (.Y(_0550_),
    .A(_0546_),
    .B(_0548_));
 sg13g2_o21ai_1 _4245_ (.B1(_0550_),
    .Y(_0551_),
    .A1(_0534_),
    .A2(_0537_));
 sg13g2_or3_1 _4246_ (.A(_0534_),
    .B(_0537_),
    .C(_0550_),
    .X(_0552_));
 sg13g2_and2_1 _4247_ (.A(_0551_),
    .B(_0552_),
    .X(_0553_));
 sg13g2_a21o_1 _4248_ (.A2(_0540_),
    .A1(_0530_),
    .B1(_0539_),
    .X(_0554_));
 sg13g2_nand2_1 _4249_ (.Y(_0555_),
    .A(_0553_),
    .B(_0554_));
 sg13g2_xor2_1 _4250_ (.B(_0554_),
    .A(_0553_),
    .X(_0556_));
 sg13g2_xnor2_1 _4251_ (.Y(_0557_),
    .A(net515),
    .B(_0556_));
 sg13g2_nor2b_1 _4252_ (.A(_0557_),
    .B_N(_0545_),
    .Y(_0558_));
 sg13g2_xnor2_1 _4253_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .A(_0545_),
    .B(_0557_));
 sg13g2_a21o_1 _4254_ (.A2(_0556_),
    .A1(net515),
    .B1(_0558_),
    .X(_0559_));
 sg13g2_nand3_1 _4255_ (.B(_0551_),
    .C(_0555_),
    .A(_0549_),
    .Y(_0560_));
 sg13g2_a21o_1 _4256_ (.A2(_0555_),
    .A1(_0551_),
    .B1(_0549_),
    .X(_0561_));
 sg13g2_nand2_2 _4257_ (.Y(_0562_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_and2_1 _4258_ (.A(net548),
    .B(_0562_),
    .X(_0563_));
 sg13g2_xor2_1 _4259_ (.B(_0562_),
    .A(net548),
    .X(_0564_));
 sg13g2_xor2_1 _4260_ (.B(_0564_),
    .A(_0559_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[14] ));
 sg13g2_a21o_1 _4261_ (.A2(_0564_),
    .A1(_0559_),
    .B1(_0563_),
    .X(_0565_));
 sg13g2_and2_1 _4262_ (.A(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .B(_0560_),
    .X(_0566_));
 sg13g2_xor2_1 _4263_ (.B(_0560_),
    .A(net578),
    .X(_0567_));
 sg13g2_xor2_1 _4264_ (.B(_0567_),
    .A(_0565_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[15] ));
 sg13g2_xor2_1 _4265_ (.B(net253),
    .A(\vgademo.soundtrack.sample_div[1] ),
    .X(\vgademo.soundtrack.sample_div_[1] ));
 sg13g2_nand3_1 _4266_ (.B(\vgademo.soundtrack.sample_div[1] ),
    .C(net253),
    .A(net475),
    .Y(_0568_));
 sg13g2_a21o_1 _4267_ (.A2(net253),
    .A1(\vgademo.soundtrack.sample_div[1] ),
    .B1(net475),
    .X(_0569_));
 sg13g2_and2_1 _4268_ (.A(_0568_),
    .B(net476),
    .X(\vgademo.soundtrack.sample_div_[2] ));
 sg13g2_nor2_1 _4269_ (.A(_3100_),
    .B(_0568_),
    .Y(_0570_));
 sg13g2_xnor2_1 _4270_ (.Y(\vgademo.soundtrack.sample_div_[3] ),
    .A(net239),
    .B(_0568_));
 sg13g2_and2_1 _4271_ (.A(net226),
    .B(_0570_),
    .X(_0571_));
 sg13g2_xor2_1 _4272_ (.B(_0570_),
    .A(net226),
    .X(\vgademo.soundtrack.sample_div_[4] ));
 sg13g2_xor2_1 _4273_ (.B(_0571_),
    .A(net268),
    .X(\vgademo.soundtrack.sample_div_[5] ));
 sg13g2_nand3_1 _4274_ (.B(net268),
    .C(_0571_),
    .A(net462),
    .Y(_0572_));
 sg13g2_a21o_1 _4275_ (.A2(_0571_),
    .A1(net268),
    .B1(net462),
    .X(_0573_));
 sg13g2_and2_1 _4276_ (.A(_0572_),
    .B(_0573_),
    .X(\vgademo.soundtrack.sample_div_[6] ));
 sg13g2_nor2_1 _4277_ (.A(_3099_),
    .B(_0572_),
    .Y(_0574_));
 sg13g2_xnor2_1 _4278_ (.Y(\vgademo.soundtrack.sample_div_[7] ),
    .A(net247),
    .B(_0572_));
 sg13g2_and2_1 _4279_ (.A(net218),
    .B(_0574_),
    .X(_0575_));
 sg13g2_xor2_1 _4280_ (.B(_0574_),
    .A(net218),
    .X(\vgademo.soundtrack.sample_div_[8] ));
 sg13g2_and2_1 _4281_ (.A(\vgademo.soundtrack.sample_div[9] ),
    .B(_0575_),
    .X(_0576_));
 sg13g2_nand2_1 _4282_ (.Y(_0577_),
    .A(\vgademo.soundtrack.sample_div[9] ),
    .B(_0575_));
 sg13g2_xor2_1 _4283_ (.B(_0575_),
    .A(net266),
    .X(\vgademo.soundtrack.sample_div_[9] ));
 sg13g2_nor4_2 _4284_ (.A(\vgademo.h_count[5] ),
    .B(net1009),
    .C(_3203_),
    .Y(_0578_),
    .D(_3210_));
 sg13g2_nor2_1 _4285_ (.A(\vgademo.h_count[9] ),
    .B(net1007),
    .Y(_0579_));
 sg13g2_nor3_2 _4286_ (.A(\vgademo.h_count[9] ),
    .B(net1007),
    .C(_0061_),
    .Y(_0580_));
 sg13g2_and2_1 _4287_ (.A(_0578_),
    .B(_0580_),
    .X(_0581_));
 sg13g2_nand2_1 _4288_ (.Y(_0582_),
    .A(_0578_),
    .B(_0580_));
 sg13g2_and2_2 _4289_ (.A(net1091),
    .B(net948),
    .X(_0583_));
 sg13g2_nand2_1 _4290_ (.Y(_0584_),
    .A(net1091),
    .B(net948));
 sg13g2_nor2_1 _4291_ (.A(net932),
    .B(net928),
    .Y(_0585_));
 sg13g2_nor3_1 _4292_ (.A(net974),
    .B(net975),
    .C(\vgademo.v_count[8] ),
    .Y(_0586_));
 sg13g2_nand2_1 _4293_ (.Y(_0587_),
    .A(net973),
    .B(_0586_));
 sg13g2_nor3_1 _4294_ (.A(net978),
    .B(net976),
    .C(_3236_),
    .Y(_0588_));
 sg13g2_nand4_1 _4295_ (.B(_3237_),
    .C(_0586_),
    .A(net973),
    .Y(_0589_),
    .D(_0588_));
 sg13g2_nor2_1 _4296_ (.A(net948),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_or2_1 _4297_ (.X(_0591_),
    .B(_0589_),
    .A(net948));
 sg13g2_nor3_1 _4298_ (.A(net978),
    .B(_3236_),
    .C(_0587_),
    .Y(_0592_));
 sg13g2_and4_2 _4299_ (.A(_3113_),
    .B(_3213_),
    .C(_3237_),
    .D(_0592_),
    .X(_0593_));
 sg13g2_a21oi_2 _4300_ (.B1(net905),
    .Y(_0594_),
    .A2(_0593_),
    .A1(net1091));
 sg13g2_nor2_1 _4301_ (.A(_3190_),
    .B(net894),
    .Y(_0595_));
 sg13g2_nor2_1 _4302_ (.A(net1066),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_nor2_1 _4303_ (.A(net1064),
    .B(net931),
    .Y(_0597_));
 sg13g2_nor2_1 _4304_ (.A(net1066),
    .B(net930),
    .Y(_0598_));
 sg13g2_nor3_1 _4305_ (.A(net893),
    .B(_0597_),
    .C(_0598_),
    .Y(_0599_));
 sg13g2_nor2_1 _4306_ (.A(_0596_),
    .B(_0599_),
    .Y(_0112_));
 sg13g2_nor3_1 _4307_ (.A(net552),
    .B(net930),
    .C(net891),
    .Y(_0600_));
 sg13g2_a21oi_1 _4308_ (.A1(_3190_),
    .A2(net891),
    .Y(_0113_),
    .B1(_0600_));
 sg13g2_nand2_1 _4309_ (.Y(_0601_),
    .A(\vgademo.linelfsr[2] ),
    .B(net891));
 sg13g2_nand2_1 _4310_ (.Y(_0602_),
    .A(net388),
    .B(net941));
 sg13g2_o21ai_1 _4311_ (.B1(_0601_),
    .Y(_0114_),
    .A1(net891),
    .A2(_0602_));
 sg13g2_xnor2_1 _4312_ (.Y(_0603_),
    .A(net1065),
    .B(net361));
 sg13g2_a21oi_1 _4313_ (.A1(net941),
    .A2(_0603_),
    .Y(_0604_),
    .B1(net891));
 sg13g2_a21o_1 _4314_ (.A2(net891),
    .A1(net388),
    .B1(_0604_),
    .X(_0115_));
 sg13g2_xnor2_1 _4315_ (.Y(_0605_),
    .A(net1065),
    .B(\vgademo.linelfsr[5] ));
 sg13g2_a21oi_1 _4316_ (.A1(net941),
    .A2(_0605_),
    .Y(_0606_),
    .B1(net891));
 sg13g2_a21o_1 _4317_ (.A2(net891),
    .A1(net361),
    .B1(_0606_),
    .X(_0116_));
 sg13g2_nor3_1 _4318_ (.A(net390),
    .B(net930),
    .C(net892),
    .Y(_0607_));
 sg13g2_a21oi_1 _4319_ (.A1(_3191_),
    .A2(net892),
    .Y(_0117_),
    .B1(_0607_));
 sg13g2_xnor2_1 _4320_ (.Y(_0608_),
    .A(net1065),
    .B(\vgademo.linelfsr[7] ));
 sg13g2_a21oi_1 _4321_ (.A1(net941),
    .A2(_0608_),
    .Y(_0609_),
    .B1(net892));
 sg13g2_a21o_1 _4322_ (.A2(net892),
    .A1(net390),
    .B1(_0609_),
    .X(_0118_));
 sg13g2_nor3_1 _4323_ (.A(net366),
    .B(net930),
    .C(net894),
    .Y(_0610_));
 sg13g2_a21oi_1 _4324_ (.A1(_3192_),
    .A2(net892),
    .Y(_0119_),
    .B1(_0610_));
 sg13g2_xnor2_1 _4325_ (.Y(_0611_),
    .A(net1066),
    .B(\vgademo.linelfsr[9] ));
 sg13g2_nor3_1 _4326_ (.A(net930),
    .B(net894),
    .C(_0611_),
    .Y(_0612_));
 sg13g2_a21o_1 _4327_ (.A2(net894),
    .A1(net366),
    .B1(_0612_),
    .X(_0120_));
 sg13g2_nor3_1 _4328_ (.A(\vgademo.linelfsr[10] ),
    .B(net930),
    .C(net893),
    .Y(_0613_));
 sg13g2_a21oi_1 _4329_ (.A1(_3193_),
    .A2(net893),
    .Y(_0121_),
    .B1(_0613_));
 sg13g2_nor3_1 _4330_ (.A(_3097_),
    .B(net930),
    .C(net893),
    .Y(_0614_));
 sg13g2_a21o_1 _4331_ (.A2(net894),
    .A1(net393),
    .B1(_0614_),
    .X(_0122_));
 sg13g2_nor3_1 _4332_ (.A(net299),
    .B(net930),
    .C(net893),
    .Y(_0615_));
 sg13g2_a21oi_1 _4333_ (.A1(_3097_),
    .A2(net893),
    .Y(_0123_),
    .B1(_0615_));
 sg13g2_nand2_1 _4334_ (.Y(_0616_),
    .A(net299),
    .B(net893));
 sg13g2_o21ai_1 _4335_ (.B1(_0616_),
    .Y(_0124_),
    .A1(net893),
    .A2(_0598_));
 sg13g2_nand3_1 _4336_ (.B(net496),
    .C(net888),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0617_));
 sg13g2_nand4_1 _4337_ (.B(\vgademo.soundtrack.tick_div[2] ),
    .C(\vgademo.soundtrack.tick_div[1] ),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0618_),
    .D(net888));
 sg13g2_nor2_1 _4338_ (.A(_3101_),
    .B(_0618_),
    .Y(_0619_));
 sg13g2_and2_1 _4339_ (.A(net209),
    .B(_0619_),
    .X(_0620_));
 sg13g2_and3_1 _4340_ (.X(_0621_),
    .A(net203),
    .B(\vgademo.soundtrack.tick_div[5] ),
    .C(_0620_));
 sg13g2_and2_2 _4341_ (.A(net230),
    .B(_0621_),
    .X(_0622_));
 sg13g2_or2_1 _4342_ (.X(_0623_),
    .B(\vgademo.audio_beat_out[0] ),
    .A(\vgademo.audio_beat_out[1] ));
 sg13g2_nor4_2 _4343_ (.A(net595),
    .B(\vgademo.audio_beat_out[2] ),
    .C(net479),
    .Y(_0624_),
    .D(_0623_));
 sg13g2_or4_2 _4344_ (.A(\vgademo.audio_beat_out[3] ),
    .B(\vgademo.audio_beat_out[2] ),
    .C(\vgademo.audio_beat_out[4] ),
    .D(_0623_),
    .X(_0625_));
 sg13g2_nand2_1 _4345_ (.Y(_0626_),
    .A(_0622_),
    .B(_0624_));
 sg13g2_nand3_1 _4346_ (.B(_0622_),
    .C(_0624_),
    .A(_3098_),
    .Y(_0627_));
 sg13g2_mux2_1 _4347_ (.A0(net1061),
    .A1(net274),
    .S(net869),
    .X(_0125_));
 sg13g2_mux2_1 _4348_ (.A0(_3267_),
    .A1(net269),
    .S(net869),
    .X(_0126_));
 sg13g2_xnor2_1 _4349_ (.Y(_0628_),
    .A(net1055),
    .B(_3270_));
 sg13g2_mux2_1 _4350_ (.A0(_0628_),
    .A1(net272),
    .S(net869),
    .X(_0127_));
 sg13g2_nor2_2 _4351_ (.A(_3271_),
    .B(_3291_),
    .Y(_0629_));
 sg13g2_nor2_2 _4352_ (.A(_3274_),
    .B(_0629_),
    .Y(_0630_));
 sg13g2_nand2_1 _4353_ (.Y(_0631_),
    .A(net189),
    .B(net870));
 sg13g2_o21ai_1 _4354_ (.B1(_0631_),
    .Y(_0128_),
    .A1(net870),
    .A2(_0630_));
 sg13g2_nand2_1 _4355_ (.Y(_0632_),
    .A(net1050),
    .B(_0629_));
 sg13g2_o21ai_1 _4356_ (.B1(net961),
    .Y(_0633_),
    .A1(_3271_),
    .A2(_3291_));
 sg13g2_and2_2 _4357_ (.A(_0632_),
    .B(_0633_),
    .X(_0634_));
 sg13g2_nand2_1 _4358_ (.Y(_0635_),
    .A(_0632_),
    .B(_0633_));
 sg13g2_nand2_1 _4359_ (.Y(_0636_),
    .A(net184),
    .B(net869));
 sg13g2_o21ai_1 _4360_ (.B1(_0636_),
    .Y(_0129_),
    .A1(net869),
    .A2(_0634_));
 sg13g2_nor3_2 _4361_ (.A(net960),
    .B(_3104_),
    .C(net958),
    .Y(_0637_));
 sg13g2_nand3_1 _4362_ (.B(_3270_),
    .C(_0637_),
    .A(net1055),
    .Y(_0638_));
 sg13g2_xnor2_1 _4363_ (.Y(_0639_),
    .A(net958),
    .B(_0632_));
 sg13g2_mux2_1 _4364_ (.A0(_0639_),
    .A1(net273),
    .S(net869),
    .X(_0130_));
 sg13g2_or2_1 _4365_ (.X(_0640_),
    .B(_0638_),
    .A(_3107_));
 sg13g2_xnor2_1 _4366_ (.Y(_0641_),
    .A(_3107_),
    .B(_0638_));
 sg13g2_mux2_1 _4367_ (.A0(_0641_),
    .A1(net280),
    .S(net870),
    .X(_0131_));
 sg13g2_xnor2_1 _4368_ (.Y(_0642_),
    .A(_3122_),
    .B(_0640_));
 sg13g2_mux2_1 _4369_ (.A0(_0642_),
    .A1(net271),
    .S(net869),
    .X(_0132_));
 sg13g2_nor4_2 _4370_ (.A(\vgademo.plane_dx_div.i[3] ),
    .B(\vgademo.plane_dx_div.i[2] ),
    .C(\vgademo.plane_dx_div.i[1] ),
    .Y(_0643_),
    .D(\vgademo.plane_dx_div.i[0] ));
 sg13g2_nor4_1 _4371_ (.A(_3118_),
    .B(_3119_),
    .C(_3120_),
    .D(net1008),
    .Y(_0644_));
 sg13g2_and3_2 _4372_ (.X(_0645_),
    .A(_3209_),
    .B(_0580_),
    .C(_0644_));
 sg13g2_nand3_1 _4373_ (.B(_0580_),
    .C(_0644_),
    .A(_3209_),
    .Y(_0646_));
 sg13g2_nor2_1 _4374_ (.A(_0643_),
    .B(net947),
    .Y(_0647_));
 sg13g2_and2_1 _4375_ (.A(_0643_),
    .B(net944),
    .X(_0648_));
 sg13g2_nand2_2 _4376_ (.Y(_0649_),
    .A(_0643_),
    .B(net944));
 sg13g2_a22oi_1 _4377_ (.Y(_0133_),
    .B1(net914),
    .B2(_3095_),
    .A2(net916),
    .A1(_3096_));
 sg13g2_a22oi_1 _4378_ (.Y(_0650_),
    .B1(net914),
    .B2(\vgademo.plane_dx[2] ),
    .A2(net916),
    .A1(net559));
 sg13g2_inv_1 _4379_ (.Y(_0134_),
    .A(net560));
 sg13g2_a22oi_1 _4380_ (.Y(_0651_),
    .B1(net913),
    .B2(net538),
    .A2(net915),
    .A1(\vgademo.plane_dx[2] ));
 sg13g2_inv_1 _4381_ (.Y(_0135_),
    .A(net539));
 sg13g2_a22oi_1 _4382_ (.Y(_0652_),
    .B1(net913),
    .B2(net187),
    .A2(net915),
    .A1(\vgademo.plane_dx[3] ));
 sg13g2_inv_1 _4383_ (.Y(_0136_),
    .A(net188));
 sg13g2_a22oi_1 _4384_ (.Y(_0653_),
    .B1(net913),
    .B2(net1042),
    .A2(net915),
    .A1(net187));
 sg13g2_inv_1 _4385_ (.Y(_0137_),
    .A(_0653_));
 sg13g2_a22oi_1 _4386_ (.Y(_0654_),
    .B1(net913),
    .B2(net1041),
    .A2(net915),
    .A1(net1042));
 sg13g2_inv_1 _4387_ (.Y(_0138_),
    .A(_0654_));
 sg13g2_a22oi_1 _4388_ (.Y(_0655_),
    .B1(net913),
    .B2(net1040),
    .A2(net915),
    .A1(net1041));
 sg13g2_inv_1 _4389_ (.Y(_0139_),
    .A(_0655_));
 sg13g2_a22oi_1 _4390_ (.Y(_0656_),
    .B1(net913),
    .B2(net216),
    .A2(net915),
    .A1(net1040));
 sg13g2_inv_1 _4391_ (.Y(_0140_),
    .A(net217));
 sg13g2_a22oi_1 _4392_ (.Y(_0657_),
    .B1(net913),
    .B2(net1038),
    .A2(net915),
    .A1(net216));
 sg13g2_inv_1 _4393_ (.Y(_0141_),
    .A(_0657_));
 sg13g2_a22oi_1 _4394_ (.Y(_0658_),
    .B1(net913),
    .B2(net1036),
    .A2(net915),
    .A1(net1038));
 sg13g2_inv_1 _4395_ (.Y(_0142_),
    .A(_0658_));
 sg13g2_o21ai_1 _4396_ (.B1(net944),
    .Y(_0143_),
    .A1(_3091_),
    .A2(_0643_));
 sg13g2_xnor2_1 _4397_ (.Y(_0659_),
    .A(\vgademo.plane_dx_div.i[1] ),
    .B(net394));
 sg13g2_nor2_1 _4398_ (.A(net947),
    .B(net395),
    .Y(_0144_));
 sg13g2_a21o_1 _4399_ (.A2(net394),
    .A1(\vgademo.plane_dx_div.i[1] ),
    .B1(net542),
    .X(_0660_));
 sg13g2_nand3_1 _4400_ (.B(\vgademo.plane_dx_div.i[1] ),
    .C(net394),
    .A(net542),
    .Y(_0661_));
 sg13g2_and3_1 _4401_ (.X(_0145_),
    .A(net944),
    .B(net543),
    .C(_0661_));
 sg13g2_xor2_1 _4402_ (.B(_0661_),
    .A(net407),
    .X(_0662_));
 sg13g2_nor2_1 _4403_ (.A(net947),
    .B(net408),
    .Y(_0146_));
 sg13g2_and2_2 _4404_ (.A(net877),
    .B(_0625_),
    .X(_0663_));
 sg13g2_nand2_2 _4405_ (.Y(_0664_),
    .A(net877),
    .B(_0625_));
 sg13g2_nor2_1 _4406_ (.A(net351),
    .B(_0663_),
    .Y(_0665_));
 sg13g2_a21oi_1 _4407_ (.A1(net351),
    .A2(_0622_),
    .Y(_0147_),
    .B1(_0665_));
 sg13g2_and3_2 _4408_ (.X(_0666_),
    .A(\vgademo.audio_beat_out[1] ),
    .B(\vgademo.audio_beat_out[0] ),
    .C(net877));
 sg13g2_nand3_1 _4409_ (.B(net351),
    .C(net877),
    .A(net374),
    .Y(_0667_));
 sg13g2_a21oi_1 _4410_ (.A1(net351),
    .A2(net877),
    .Y(_0668_),
    .B1(net374));
 sg13g2_o21ai_1 _4411_ (.B1(_0627_),
    .Y(_0148_),
    .A1(_0666_),
    .A2(_0668_));
 sg13g2_o21ai_1 _4412_ (.B1(net870),
    .Y(_0669_),
    .A1(net465),
    .A2(_0667_));
 sg13g2_mux2_1 _4413_ (.A0(_3102_),
    .A1(net465),
    .S(net877),
    .X(_0670_));
 sg13g2_a21oi_1 _4414_ (.A1(_0667_),
    .A2(_0670_),
    .Y(_0149_),
    .B1(_0669_));
 sg13g2_nand3b_1 _4415_ (.B(_0666_),
    .C(net518),
    .Y(_0671_),
    .A_N(net465));
 sg13g2_o21ai_1 _4416_ (.B1(_0671_),
    .Y(_0672_),
    .A1(net518),
    .A2(_0669_));
 sg13g2_nor2b_1 _4417_ (.A(_0672_),
    .B_N(_0627_),
    .Y(_0150_));
 sg13g2_nand3_1 _4418_ (.B(\vgademo.audio_beat_out[2] ),
    .C(_0666_),
    .A(\vgademo.audio_beat_out[3] ),
    .Y(_0673_));
 sg13g2_xor2_1 _4419_ (.B(_0673_),
    .A(net479),
    .X(_0674_));
 sg13g2_nand2_1 _4420_ (.Y(_0151_),
    .A(_0627_),
    .B(net480));
 sg13g2_nand2_1 _4421_ (.Y(_0675_),
    .A(net1047),
    .B(_0630_));
 sg13g2_a21oi_1 _4422_ (.A1(net1058),
    .A2(net1056),
    .Y(_0676_),
    .B1(net1053));
 sg13g2_nand3b_1 _4423_ (.B(_0634_),
    .C(_0675_),
    .Y(_0677_),
    .A_N(_0676_));
 sg13g2_or2_1 _4424_ (.X(_0678_),
    .B(_0639_),
    .A(_3107_));
 sg13g2_nand3_1 _4425_ (.B(_0630_),
    .C(_0639_),
    .A(_3278_),
    .Y(_0679_));
 sg13g2_nand2_1 _4426_ (.Y(_0680_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_a22oi_1 _4427_ (.Y(_0681_),
    .B1(_0680_),
    .B2(_0634_),
    .A2(_0677_),
    .A1(_3271_));
 sg13g2_o21ai_1 _4428_ (.B1(net877),
    .Y(_0682_),
    .A1(_0625_),
    .A2(_0681_));
 sg13g2_nand3_1 _4429_ (.B(net1053),
    .C(_3254_),
    .A(net1050),
    .Y(_0683_));
 sg13g2_nand4_1 _4430_ (.B(net961),
    .C(_3263_),
    .A(net1058),
    .Y(_0684_),
    .D(_3291_));
 sg13g2_and2_1 _4431_ (.A(net1047),
    .B(_0684_),
    .X(_0685_));
 sg13g2_nor2_1 _4432_ (.A(net1058),
    .B(net959),
    .Y(_0686_));
 sg13g2_nor2_2 _4433_ (.A(net961),
    .B(net1053),
    .Y(_0687_));
 sg13g2_and2_1 _4434_ (.A(_0686_),
    .B(_0687_),
    .X(_0688_));
 sg13g2_a21oi_1 _4435_ (.A1(net961),
    .A2(_3254_),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_a22oi_1 _4436_ (.Y(_0690_),
    .B1(_0689_),
    .B2(_3106_),
    .A2(_0685_),
    .A1(_0683_));
 sg13g2_inv_1 _4437_ (.Y(_0691_),
    .A(_0690_));
 sg13g2_nor2_2 _4438_ (.A(_3290_),
    .B(_0691_),
    .Y(_0692_));
 sg13g2_nor3_2 _4439_ (.A(\vgademo.audio_kick_frames[1] ),
    .B(\vgademo.audio_kick_frames[0] ),
    .C(_3108_),
    .Y(_0693_));
 sg13g2_or3_2 _4440_ (.A(\vgademo.audio_kick_frames[1] ),
    .B(\vgademo.audio_kick_frames[0] ),
    .C(_3108_),
    .X(_0694_));
 sg13g2_nand2_1 _4441_ (.Y(_0695_),
    .A(_3254_),
    .B(_0687_));
 sg13g2_nand2_1 _4442_ (.Y(_0696_),
    .A(net1047),
    .B(_0687_));
 sg13g2_nor2_1 _4443_ (.A(_3253_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_nor2_1 _4444_ (.A(_0690_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_nor3_1 _4445_ (.A(_0692_),
    .B(_0694_),
    .C(_0698_),
    .Y(_0699_));
 sg13g2_nor2_1 _4446_ (.A(_0624_),
    .B(_0694_),
    .Y(_0700_));
 sg13g2_nor2b_1 _4447_ (.A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[3] ),
    .Y(_0701_));
 sg13g2_xor2_1 _4448_ (.B(\vgademo.soundtrack.tri_osc_i[3] ),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(_0702_));
 sg13g2_o21ai_1 _4449_ (.B1(_0625_),
    .Y(_0703_),
    .A1(_0693_),
    .A2(_0702_));
 sg13g2_a21oi_1 _4450_ (.A1(net1058),
    .A2(net1053),
    .Y(_0704_),
    .B1(_0676_));
 sg13g2_nor2_1 _4451_ (.A(_3253_),
    .B(_0686_),
    .Y(_0705_));
 sg13g2_or2_2 _4452_ (.X(_0706_),
    .B(_0686_),
    .A(_3253_));
 sg13g2_a22oi_1 _4453_ (.Y(_0707_),
    .B1(_0706_),
    .B2(net1049),
    .A2(_3295_),
    .A1(_3264_));
 sg13g2_nand2_1 _4454_ (.Y(_0708_),
    .A(net1047),
    .B(_0707_));
 sg13g2_o21ai_1 _4455_ (.B1(_0708_),
    .Y(_0709_),
    .A1(_3283_),
    .A2(_0704_));
 sg13g2_o21ai_1 _4456_ (.B1(_3290_),
    .Y(_0710_),
    .A1(net1053),
    .A2(_0705_));
 sg13g2_nand2b_2 _4457_ (.Y(_0711_),
    .B(_0710_),
    .A_N(_0709_));
 sg13g2_nor2_2 _4458_ (.A(net950),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_nor4_1 _4459_ (.A(net868),
    .B(_0699_),
    .C(_0703_),
    .D(_0712_),
    .Y(_0713_));
 sg13g2_a21o_1 _4460_ (.A2(net868),
    .A1(net485),
    .B1(_0713_),
    .X(_0152_));
 sg13g2_nand2_1 _4461_ (.Y(_0714_),
    .A(net486),
    .B(net868));
 sg13g2_nor2b_1 _4462_ (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[1] ),
    .Y(_0715_));
 sg13g2_xnor2_1 _4463_ (.Y(_0716_),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .B(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_nor2b_1 _4464_ (.A(_0701_),
    .B_N(_0716_),
    .Y(_0717_));
 sg13g2_xnor2_1 _4465_ (.Y(_0718_),
    .A(_0701_),
    .B(_0716_));
 sg13g2_or3_1 _4466_ (.A(_0692_),
    .B(_0698_),
    .C(_0711_),
    .X(_0719_));
 sg13g2_a21oi_1 _4467_ (.A1(_0692_),
    .A2(_0709_),
    .Y(_0720_),
    .B1(net950));
 sg13g2_a22oi_1 _4468_ (.Y(_0721_),
    .B1(_0719_),
    .B2(_0720_),
    .A2(_0718_),
    .A1(_0694_));
 sg13g2_o21ai_1 _4469_ (.B1(_0714_),
    .Y(_0153_),
    .A1(_0664_),
    .A2(_0721_));
 sg13g2_nand2_1 _4470_ (.Y(_0722_),
    .A(net451),
    .B(net867));
 sg13g2_nand2b_1 _4471_ (.Y(_0723_),
    .B(\vgademo.soundtrack.tri_osc_i[2] ),
    .A_N(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_xnor2_1 _4472_ (.Y(_0724_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_o21ai_1 _4473_ (.B1(_0724_),
    .Y(_0725_),
    .A1(_0715_),
    .A2(_0717_));
 sg13g2_or3_1 _4474_ (.A(_0715_),
    .B(_0717_),
    .C(_0724_),
    .X(_0726_));
 sg13g2_a21oi_1 _4475_ (.A1(_0725_),
    .A2(_0726_),
    .Y(_0727_),
    .B1(_0693_));
 sg13g2_a21oi_1 _4476_ (.A1(_3263_),
    .A2(_3292_),
    .Y(_0728_),
    .B1(net960));
 sg13g2_nor2_1 _4477_ (.A(net1046),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_a21oi_1 _4478_ (.A1(_0695_),
    .A2(_0729_),
    .Y(_0730_),
    .B1(_0697_));
 sg13g2_nand2_1 _4479_ (.Y(_0731_),
    .A(_3253_),
    .B(_0687_));
 sg13g2_a22oi_1 _4480_ (.Y(_0732_),
    .B1(_0731_),
    .B2(_0685_),
    .A2(_0688_),
    .A1(net958));
 sg13g2_nor2b_1 _4481_ (.A(_0732_),
    .B_N(_0730_),
    .Y(_0733_));
 sg13g2_and2_1 _4482_ (.A(_0691_),
    .B(_0733_),
    .X(_0734_));
 sg13g2_o21ai_1 _4483_ (.B1(_0693_),
    .Y(_0735_),
    .A1(_0692_),
    .A2(_0711_));
 sg13g2_o21ai_1 _4484_ (.B1(_0663_),
    .Y(_0736_),
    .A1(_0734_),
    .A2(_0735_));
 sg13g2_o21ai_1 _4485_ (.B1(_0722_),
    .Y(_0154_),
    .A1(_0727_),
    .A2(_0736_));
 sg13g2_nand2_1 _4486_ (.Y(_0737_),
    .A(net510),
    .B(net868));
 sg13g2_and2_1 _4487_ (.A(_0730_),
    .B(_0732_),
    .X(_0738_));
 sg13g2_or2_1 _4488_ (.X(_0739_),
    .B(_0738_),
    .A(_0690_));
 sg13g2_inv_1 _4489_ (.Y(_0740_),
    .A(_0739_));
 sg13g2_nor2_1 _4490_ (.A(_0687_),
    .B(_0739_),
    .Y(_0741_));
 sg13g2_a21oi_1 _4491_ (.A1(_0690_),
    .A2(_0738_),
    .Y(_0742_),
    .B1(_0741_));
 sg13g2_and2_1 _4492_ (.A(_0693_),
    .B(_0711_),
    .X(_0743_));
 sg13g2_nand2_1 _4493_ (.Y(_0744_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(_3139_));
 sg13g2_xor2_1 _4494_ (.B(\vgademo.soundtrack.tri_osc_i[6] ),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .X(_0745_));
 sg13g2_a21o_1 _4495_ (.A2(_0725_),
    .A1(_0723_),
    .B1(_0745_),
    .X(_0746_));
 sg13g2_nand3_1 _4496_ (.B(_0725_),
    .C(_0745_),
    .A(_0723_),
    .Y(_0747_));
 sg13g2_and3_1 _4497_ (.X(_0748_),
    .A(net950),
    .B(_0746_),
    .C(_0747_));
 sg13g2_a221oi_1 _4498_ (.B2(_0743_),
    .C1(_0748_),
    .B1(_0742_),
    .A1(_0712_),
    .Y(_0749_),
    .A2(_0734_));
 sg13g2_o21ai_1 _4499_ (.B1(_0737_),
    .Y(_0155_),
    .A1(_0664_),
    .A2(_0749_));
 sg13g2_nand2_1 _4500_ (.Y(_0750_),
    .A(net519),
    .B(net867));
 sg13g2_xor2_1 _4501_ (.B(\vgademo.soundtrack.tri_osc_i[7] ),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(_0751_));
 sg13g2_a21oi_1 _4502_ (.A1(_0744_),
    .A2(_0746_),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_and3_1 _4503_ (.X(_0753_),
    .A(_0744_),
    .B(_0746_),
    .C(_0751_));
 sg13g2_nor3_1 _4504_ (.A(_0693_),
    .B(_0752_),
    .C(_0753_),
    .Y(_0754_));
 sg13g2_nor2_1 _4505_ (.A(_0692_),
    .B(_0733_),
    .Y(_0755_));
 sg13g2_a221oi_1 _4506_ (.B2(_0755_),
    .C1(_0754_),
    .B1(_0743_),
    .A1(_0712_),
    .Y(_0756_),
    .A2(_0742_));
 sg13g2_o21ai_1 _4507_ (.B1(_0750_),
    .Y(_0156_),
    .A1(_0664_),
    .A2(_0756_));
 sg13g2_nand2_1 _4508_ (.Y(_0757_),
    .A(net540),
    .B(net867));
 sg13g2_a21oi_1 _4509_ (.A1(\vgademo.soundtrack.tri_osc_i[4] ),
    .A2(_3140_),
    .Y(_0758_),
    .B1(_0752_));
 sg13g2_nor2_1 _4510_ (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(_3141_),
    .Y(_0759_));
 sg13g2_nand2_1 _4511_ (.Y(_0760_),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(_3141_));
 sg13g2_nand2b_1 _4512_ (.Y(_0761_),
    .B(_0760_),
    .A_N(_0759_));
 sg13g2_o21ai_1 _4513_ (.B1(net950),
    .Y(_0762_),
    .A1(_0758_),
    .A2(_0761_));
 sg13g2_a21oi_1 _4514_ (.A1(_0758_),
    .A2(_0761_),
    .Y(_0763_),
    .B1(_0762_));
 sg13g2_a221oi_1 _4515_ (.B2(_0712_),
    .C1(_0763_),
    .B1(_0755_),
    .A1(_0740_),
    .Y(_0764_),
    .A2(_0743_));
 sg13g2_o21ai_1 _4516_ (.B1(_0757_),
    .Y(_0157_),
    .A1(_0664_),
    .A2(_0764_));
 sg13g2_o21ai_1 _4517_ (.B1(_0760_),
    .Y(_0765_),
    .A1(_0758_),
    .A2(_0759_));
 sg13g2_xnor2_1 _4518_ (.Y(_0766_),
    .A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(_0765_));
 sg13g2_nand2b_1 _4519_ (.Y(_0767_),
    .B(_0738_),
    .A_N(_0711_));
 sg13g2_nor2_1 _4520_ (.A(_0690_),
    .B(net950),
    .Y(_0768_));
 sg13g2_a22oi_1 _4521_ (.Y(_0769_),
    .B1(_0767_),
    .B2(_0768_),
    .A2(_0766_),
    .A1(net950));
 sg13g2_a22oi_1 _4522_ (.Y(_0158_),
    .B1(_0769_),
    .B2(_0663_),
    .A2(net867),
    .A1(_3139_));
 sg13g2_nor3_1 _4523_ (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(\vgademo.soundtrack.tri_osc_i[7] ),
    .C(_0765_),
    .Y(_0770_));
 sg13g2_o21ai_1 _4524_ (.B1(\vgademo.soundtrack.tri_osc_i[7] ),
    .Y(_0771_),
    .A1(\vgademo.soundtrack.tri_osc_i[6] ),
    .A2(_0765_));
 sg13g2_nand2b_1 _4525_ (.Y(_0772_),
    .B(_0771_),
    .A_N(_0770_));
 sg13g2_nor2_1 _4526_ (.A(_0743_),
    .B(_0768_),
    .Y(_0773_));
 sg13g2_a21oi_1 _4527_ (.A1(_0691_),
    .A2(_0711_),
    .Y(_0774_),
    .B1(_0773_));
 sg13g2_a21oi_1 _4528_ (.A1(net950),
    .A2(_0772_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_a22oi_1 _4529_ (.Y(_0159_),
    .B1(_0775_),
    .B2(_0663_),
    .A2(net867),
    .A1(_3140_));
 sg13g2_o21ai_1 _4530_ (.B1(net950),
    .Y(_0776_),
    .A1(_3141_),
    .A2(_0770_));
 sg13g2_nand2_1 _4531_ (.Y(_0777_),
    .A(_0773_),
    .B(_0776_));
 sg13g2_a22oi_1 _4532_ (.Y(_0160_),
    .B1(_0777_),
    .B2(_0663_),
    .A2(net867),
    .A1(_3141_));
 sg13g2_nor2_1 _4533_ (.A(net1079),
    .B(net197),
    .Y(_0778_));
 sg13g2_a21oi_2 _4534_ (.B1(_0566_),
    .Y(_0779_),
    .A2(_0567_),
    .A1(_0565_));
 sg13g2_a21oi_1 _4535_ (.A1(net1077),
    .A2(_0779_),
    .Y(_0161_),
    .B1(_0778_));
 sg13g2_mux2_1 _4536_ (.A0(\vgademo.soundtrack.tick_div[0] ),
    .A1(net178),
    .S(net888),
    .X(_0162_));
 sg13g2_a21o_1 _4537_ (.A2(net888),
    .A1(\vgademo.soundtrack.tick_div[0] ),
    .B1(net496),
    .X(_0780_));
 sg13g2_and2_1 _4538_ (.A(_0617_),
    .B(net497),
    .X(_0163_));
 sg13g2_xnor2_1 _4539_ (.Y(_0164_),
    .A(net264),
    .B(_0617_));
 sg13g2_xnor2_1 _4540_ (.Y(_0165_),
    .A(net243),
    .B(_0618_));
 sg13g2_xor2_1 _4541_ (.B(_0619_),
    .A(net209),
    .X(_0166_));
 sg13g2_xor2_1 _4542_ (.B(_0620_),
    .A(net262),
    .X(_0167_));
 sg13g2_a21oi_1 _4543_ (.A1(\vgademo.soundtrack.tick_div[5] ),
    .A2(_0620_),
    .Y(_0781_),
    .B1(net203));
 sg13g2_nor2_1 _4544_ (.A(_0621_),
    .B(net204),
    .Y(_0168_));
 sg13g2_xor2_1 _4545_ (.B(_0621_),
    .A(net230),
    .X(_0169_));
 sg13g2_nand2_1 _4546_ (.Y(_0782_),
    .A(_0094_),
    .B(net887));
 sg13g2_o21ai_1 _4547_ (.B1(_0782_),
    .Y(_0170_),
    .A1(net170),
    .A2(net887));
 sg13g2_nand2_1 _4548_ (.Y(_0783_),
    .A(_0095_),
    .B(net886));
 sg13g2_o21ai_1 _4549_ (.B1(_0783_),
    .Y(_0171_),
    .A1(net166),
    .A2(net887));
 sg13g2_nand2_1 _4550_ (.Y(_0784_),
    .A(_0096_),
    .B(net887));
 sg13g2_o21ai_1 _4551_ (.B1(_0784_),
    .Y(_0172_),
    .A1(net182),
    .A2(net886));
 sg13g2_mux2_1 _4552_ (.A0(net228),
    .A1(_0040_),
    .S(net888),
    .X(_0173_));
 sg13g2_mux2_1 _4553_ (.A0(net233),
    .A1(\vgademo.soundtrack.noise_lfsr[5] ),
    .S(net888),
    .X(_0174_));
 sg13g2_mux2_1 _4554_ (.A0(_0098_),
    .A1(net174),
    .S(net888),
    .X(_0175_));
 sg13g2_mux2_1 _4555_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(net276),
    .S(net889),
    .X(_0176_));
 sg13g2_mux2_1 _4556_ (.A0(_0099_),
    .A1(net176),
    .S(net889),
    .X(_0177_));
 sg13g2_mux2_1 _4557_ (.A0(net323),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net889),
    .X(_0178_));
 sg13g2_mux2_1 _4558_ (.A0(net185),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net886),
    .X(_0179_));
 sg13g2_nand2_1 _4559_ (.Y(_0785_),
    .A(_0100_),
    .B(net886));
 sg13g2_o21ai_1 _4560_ (.B1(_0785_),
    .Y(_0180_),
    .A1(net180),
    .A2(net886));
 sg13g2_nand2_1 _4561_ (.Y(_0786_),
    .A(_0101_),
    .B(net886));
 sg13g2_o21ai_1 _4562_ (.B1(_0786_),
    .Y(_0181_),
    .A1(net172),
    .A2(net886));
 sg13g2_mux2_1 _4563_ (.A0(_0102_),
    .A1(net201),
    .S(net888),
    .X(_0182_));
 sg13g2_xor2_1 _4564_ (.B(\vgademo.soundtrack.noise_lfsr[14] ),
    .A(\vgademo.soundtrack.noise_lfsr[0] ),
    .X(_0787_));
 sg13g2_mux2_1 _4565_ (.A0(net241),
    .A1(_0787_),
    .S(net889),
    .X(_0183_));
 sg13g2_mux2_1 _4566_ (.A0(\vgademo.soundtrack.noise_lfsr[0] ),
    .A1(net332),
    .S(net886),
    .X(_0184_));
 sg13g2_nand3_1 _4567_ (.B(net1035),
    .C(net1026),
    .A(net1031),
    .Y(_0788_));
 sg13g2_or2_1 _4568_ (.X(_0789_),
    .B(_0788_),
    .A(_3146_));
 sg13g2_nand2_1 _4569_ (.Y(_0790_),
    .A(net1035),
    .B(_0789_));
 sg13g2_nand3_1 _4570_ (.B(_3265_),
    .C(_0630_),
    .A(_3257_),
    .Y(_0791_));
 sg13g2_nand2_1 _4571_ (.Y(_0792_),
    .A(net1051),
    .B(_0630_));
 sg13g2_o21ai_1 _4572_ (.B1(_0792_),
    .Y(_0793_),
    .A1(net1060),
    .A2(_3258_));
 sg13g2_a21oi_1 _4573_ (.A1(_0791_),
    .A2(_0793_),
    .Y(_0794_),
    .B1(_0641_));
 sg13g2_nand2_1 _4574_ (.Y(_0795_),
    .A(_3098_),
    .B(_3291_));
 sg13g2_nand4_1 _4575_ (.B(net1048),
    .C(_3271_),
    .A(net1050),
    .Y(_0796_),
    .D(_0795_));
 sg13g2_a21oi_1 _4576_ (.A1(_0678_),
    .A2(_0796_),
    .Y(_0797_),
    .B1(_0794_));
 sg13g2_a21oi_1 _4577_ (.A1(_3257_),
    .A2(_3296_),
    .Y(_0798_),
    .B1(net1048));
 sg13g2_or3_1 _4578_ (.A(net1060),
    .B(net1051),
    .C(_3258_),
    .X(_0799_));
 sg13g2_a21oi_1 _4579_ (.A1(_0634_),
    .A2(_0798_),
    .Y(_0800_),
    .B1(_0797_));
 sg13g2_a21oi_2 _4580_ (.B1(net869),
    .Y(_0801_),
    .A2(_0800_),
    .A1(_0799_));
 sg13g2_nor2_2 _4581_ (.A(_0666_),
    .B(_0801_),
    .Y(_0802_));
 sg13g2_a22oi_1 _4582_ (.Y(_0185_),
    .B1(_0802_),
    .B2(_3088_),
    .A2(_0790_),
    .A1(_0666_));
 sg13g2_xnor2_1 _4583_ (.Y(_0803_),
    .A(net1031),
    .B(net1035));
 sg13g2_nand2_1 _4584_ (.Y(_0804_),
    .A(_0789_),
    .B(_0803_));
 sg13g2_a22oi_1 _4585_ (.Y(_0186_),
    .B1(_0804_),
    .B2(_0666_),
    .A2(_0802_),
    .A1(_3087_));
 sg13g2_a21oi_1 _4586_ (.A1(net1031),
    .A2(net1035),
    .Y(_0805_),
    .B1(net1026));
 sg13g2_nor2_1 _4587_ (.A(net1023),
    .B(_0788_),
    .Y(_0806_));
 sg13g2_nor2_1 _4588_ (.A(_0805_),
    .B(_0806_),
    .Y(_0807_));
 sg13g2_a22oi_1 _4589_ (.Y(_0187_),
    .B1(_0807_),
    .B2(_0666_),
    .A2(_0802_),
    .A1(_3086_));
 sg13g2_a21oi_1 _4590_ (.A1(_3146_),
    .A2(_0788_),
    .Y(_0808_),
    .B1(_0667_));
 sg13g2_a21oi_1 _4591_ (.A1(_3085_),
    .A2(_0802_),
    .Y(_0188_),
    .B1(_0808_));
 sg13g2_and2_1 _4592_ (.A(net1071),
    .B(net889),
    .X(_0809_));
 sg13g2_nand2_1 _4593_ (.Y(_0810_),
    .A(net1071),
    .B(net889));
 sg13g2_a21o_1 _4594_ (.A2(net1056),
    .A1(net1058),
    .B1(_3104_),
    .X(_0811_));
 sg13g2_a22oi_1 _4595_ (.Y(_0812_),
    .B1(_3275_),
    .B2(_0811_),
    .A2(_3271_),
    .A1(net959));
 sg13g2_nor2b_1 _4596_ (.A(_3259_),
    .B_N(_3295_),
    .Y(_0813_));
 sg13g2_o21ai_1 _4597_ (.B1(net1050),
    .Y(_0814_),
    .A1(_0628_),
    .A2(_0813_));
 sg13g2_o21ai_1 _4598_ (.B1(_0814_),
    .Y(_0815_),
    .A1(net1049),
    .A2(_0812_));
 sg13g2_nand2_1 _4599_ (.Y(_0816_),
    .A(net1062),
    .B(_3104_));
 sg13g2_and2_1 _4600_ (.A(net954),
    .B(_0686_),
    .X(_0817_));
 sg13g2_a22oi_1 _4601_ (.Y(_0818_),
    .B1(_0816_),
    .B2(_0817_),
    .A2(_0815_),
    .A1(net1046));
 sg13g2_nor2_1 _4602_ (.A(net1054),
    .B(net959),
    .Y(_0819_));
 sg13g2_nor2_1 _4603_ (.A(_3268_),
    .B(_0819_),
    .Y(_0820_));
 sg13g2_nor3_1 _4604_ (.A(net958),
    .B(_3268_),
    .C(_0819_),
    .Y(_0821_));
 sg13g2_a21oi_1 _4605_ (.A1(_0633_),
    .A2(_0821_),
    .Y(_0822_),
    .B1(net1045));
 sg13g2_nand3_1 _4606_ (.B(_3263_),
    .C(_3292_),
    .A(net1049),
    .Y(_0823_));
 sg13g2_nand2_1 _4607_ (.Y(_0824_),
    .A(net958),
    .B(_0823_));
 sg13g2_a21oi_1 _4608_ (.A1(_0822_),
    .A2(_0824_),
    .Y(_0825_),
    .B1(_3107_));
 sg13g2_o21ai_1 _4609_ (.B1(_0825_),
    .Y(_0826_),
    .A1(_3122_),
    .A2(_0818_));
 sg13g2_o21ai_1 _4610_ (.B1(_0826_),
    .Y(_0827_),
    .A1(net1046),
    .A2(\vgademo.audio_songpos[6] ));
 sg13g2_nor2_1 _4611_ (.A(_3098_),
    .B(_0819_),
    .Y(_0828_));
 sg13g2_a221oi_1 _4612_ (.B2(_0828_),
    .C1(net1049),
    .B1(_0705_),
    .A1(_3256_),
    .Y(_0829_),
    .A2(_3262_));
 sg13g2_nand2_2 _4613_ (.Y(_0830_),
    .A(_3104_),
    .B(_3272_));
 sg13g2_nor2_1 _4614_ (.A(_3259_),
    .B(_3270_),
    .Y(_0831_));
 sg13g2_nand3_1 _4615_ (.B(_0830_),
    .C(_0831_),
    .A(_3296_),
    .Y(_0832_));
 sg13g2_o21ai_1 _4616_ (.B1(_0637_),
    .Y(_0833_),
    .A1(net959),
    .A2(_3271_));
 sg13g2_o21ai_1 _4617_ (.B1(_3282_),
    .Y(_0834_),
    .A1(net1055),
    .A2(_0813_));
 sg13g2_nand2b_1 _4618_ (.Y(_0835_),
    .B(_0830_),
    .A_N(_0834_));
 sg13g2_nand2_1 _4619_ (.Y(_0836_),
    .A(_0833_),
    .B(_0835_));
 sg13g2_a221oi_1 _4620_ (.B2(net954),
    .C1(_0836_),
    .B1(_0832_),
    .A1(net1046),
    .Y(_0837_),
    .A2(_0829_));
 sg13g2_nand2_2 _4621_ (.Y(_0838_),
    .A(_3102_),
    .B(\vgademo.audio_songpos[6] ));
 sg13g2_o21ai_1 _4622_ (.B1(net1048),
    .Y(_0839_),
    .A1(net961),
    .A2(_3104_));
 sg13g2_nor2b_1 _4623_ (.A(_0839_),
    .B_N(_0633_),
    .Y(_0840_));
 sg13g2_nor2_1 _4624_ (.A(net1045),
    .B(_0840_),
    .Y(_0841_));
 sg13g2_nand3_1 _4625_ (.B(net1052),
    .C(_0706_),
    .A(net960),
    .Y(_0842_));
 sg13g2_nand2_1 _4626_ (.Y(_0843_),
    .A(_0729_),
    .B(_0842_));
 sg13g2_a21oi_1 _4627_ (.A1(_0841_),
    .A2(_0843_),
    .Y(_0844_),
    .B1(_0838_));
 sg13g2_o21ai_1 _4628_ (.B1(_0844_),
    .Y(_0845_),
    .A1(_3122_),
    .A2(_0837_));
 sg13g2_nor2_1 _4629_ (.A(\vgademo.audio_beat_out[2] ),
    .B(\vgademo.audio_songpos[6] ),
    .Y(_0846_));
 sg13g2_nor2b_1 _4630_ (.A(_0696_),
    .B_N(_0846_),
    .Y(_0847_));
 sg13g2_a21oi_1 _4631_ (.A1(\vgademo.audio_beat_out[2] ),
    .A2(_0827_),
    .Y(_0848_),
    .B1(_0847_));
 sg13g2_nand2_2 _4632_ (.Y(_0849_),
    .A(_0845_),
    .B(_0848_));
 sg13g2_inv_2 _4633_ (.Y(_0850_),
    .A(_0849_));
 sg13g2_nand3_1 _4634_ (.B(net954),
    .C(_0706_),
    .A(net1052),
    .Y(_0851_));
 sg13g2_nand4_1 _4635_ (.B(_3296_),
    .C(_0830_),
    .A(net954),
    .Y(_0852_),
    .D(_0831_));
 sg13g2_a21o_1 _4636_ (.A2(_0687_),
    .A1(_3265_),
    .B1(net958),
    .X(_0853_));
 sg13g2_inv_1 _4637_ (.Y(_0854_),
    .A(_0853_));
 sg13g2_o21ai_1 _4638_ (.B1(_3282_),
    .Y(_0855_),
    .A1(_3274_),
    .A2(_3293_));
 sg13g2_nand3_1 _4639_ (.B(_0853_),
    .C(_0855_),
    .A(_0852_),
    .Y(_0856_));
 sg13g2_a22oi_1 _4640_ (.Y(_0857_),
    .B1(_0856_),
    .B2(net1045),
    .A2(_0851_),
    .A1(_0841_));
 sg13g2_nor2b_1 _4641_ (.A(net954),
    .B_N(_0846_),
    .Y(_0858_));
 sg13g2_nand3_1 _4642_ (.B(_3263_),
    .C(_3295_),
    .A(net1049),
    .Y(_0859_));
 sg13g2_nand3_1 _4643_ (.B(_0812_),
    .C(_0859_),
    .A(net1046),
    .Y(_0860_));
 sg13g2_nor3_1 _4644_ (.A(_3253_),
    .B(_3283_),
    .C(_0629_),
    .Y(_0861_));
 sg13g2_a221oi_1 _4645_ (.B2(_3275_),
    .C1(_3122_),
    .B1(_0861_),
    .A1(net954),
    .Y(_0862_),
    .A2(_0629_));
 sg13g2_nor2_1 _4646_ (.A(_3266_),
    .B(_0819_),
    .Y(_0863_));
 sg13g2_o21ai_1 _4647_ (.B1(_0822_),
    .Y(_0864_),
    .A1(_3283_),
    .A2(_0863_));
 sg13g2_nand3_1 _4648_ (.B(\vgademo.audio_songpos[6] ),
    .C(_0864_),
    .A(\vgademo.audio_beat_out[2] ),
    .Y(_0865_));
 sg13g2_a21oi_1 _4649_ (.A1(_0860_),
    .A2(_0862_),
    .Y(_0866_),
    .B1(_0865_));
 sg13g2_a21oi_1 _4650_ (.A1(_0696_),
    .A2(_0858_),
    .Y(_0867_),
    .B1(_0866_));
 sg13g2_o21ai_1 _4651_ (.B1(_0867_),
    .Y(_0868_),
    .A1(_0838_),
    .A2(_0857_));
 sg13g2_o21ai_1 _4652_ (.B1(_0854_),
    .Y(_0869_),
    .A1(net1049),
    .A2(_0812_));
 sg13g2_a21oi_1 _4653_ (.A1(_0824_),
    .A2(_0839_),
    .Y(_0870_),
    .B1(net1045));
 sg13g2_a21oi_1 _4654_ (.A1(net1045),
    .A2(_0869_),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_o21ai_1 _4655_ (.B1(_0871_),
    .Y(_0872_),
    .A1(\vgademo.audio_songpos[6] ),
    .A2(_0637_));
 sg13g2_o21ai_1 _4656_ (.B1(net1046),
    .Y(_0873_),
    .A1(net1052),
    .A2(_3265_));
 sg13g2_o21ai_1 _4657_ (.B1(net1045),
    .Y(_0874_),
    .A1(_0829_),
    .A2(_0873_));
 sg13g2_inv_1 _4658_ (.Y(_0875_),
    .A(_0874_));
 sg13g2_a21oi_1 _4659_ (.A1(net1046),
    .A2(_0634_),
    .Y(_0876_),
    .B1(_0728_));
 sg13g2_a22oi_1 _4660_ (.Y(_0877_),
    .B1(_0876_),
    .B2(_3122_),
    .A2(_0875_),
    .A1(_0835_));
 sg13g2_a22oi_1 _4661_ (.Y(_0878_),
    .B1(_0872_),
    .B2(\vgademo.audio_beat_out[2] ),
    .A2(_0846_),
    .A1(net960));
 sg13g2_o21ai_1 _4662_ (.B1(_0878_),
    .Y(_0879_),
    .A1(_0838_),
    .A2(_0877_));
 sg13g2_nand2b_1 _4663_ (.Y(_0880_),
    .B(_0879_),
    .A_N(_0868_));
 sg13g2_nand2_2 _4664_ (.Y(_0881_),
    .A(_0850_),
    .B(_0880_));
 sg13g2_o21ai_1 _4665_ (.B1(_0849_),
    .Y(_0882_),
    .A1(_0868_),
    .A2(_0879_));
 sg13g2_nand2_1 _4666_ (.Y(_0883_),
    .A(_0881_),
    .B(_0882_));
 sg13g2_nand2_1 _4667_ (.Y(_0884_),
    .A(net882),
    .B(_0883_));
 sg13g2_xnor2_1 _4668_ (.Y(_0189_),
    .A(net286),
    .B(_0884_));
 sg13g2_nand2b_1 _4669_ (.Y(_0885_),
    .B(_0881_),
    .A_N(_0042_));
 sg13g2_xnor2_1 _4670_ (.Y(_0886_),
    .A(_0042_),
    .B(_0881_));
 sg13g2_nand3_1 _4671_ (.B(_0883_),
    .C(_0886_),
    .A(\vgademo.soundtrack.pulse_osc_p[0] ),
    .Y(_0887_));
 sg13g2_a21o_1 _4672_ (.A2(_0883_),
    .A1(\vgademo.soundtrack.pulse_osc_p[0] ),
    .B1(_0886_),
    .X(_0888_));
 sg13g2_a21oi_1 _4673_ (.A1(_0887_),
    .A2(_0888_),
    .Y(_0889_),
    .B1(net880));
 sg13g2_a21oi_1 _4674_ (.A1(_3197_),
    .A2(net880),
    .Y(_0190_),
    .B1(_0889_));
 sg13g2_nor2_1 _4675_ (.A(net313),
    .B(net881),
    .Y(_0890_));
 sg13g2_nand2_1 _4676_ (.Y(_0891_),
    .A(_0885_),
    .B(_0887_));
 sg13g2_o21ai_1 _4677_ (.B1(_0850_),
    .Y(_0892_),
    .A1(_0868_),
    .A2(_0879_));
 sg13g2_nand2b_1 _4678_ (.Y(_0893_),
    .B(_0868_),
    .A_N(_0879_));
 sg13g2_nand2_1 _4679_ (.Y(_0894_),
    .A(_0849_),
    .B(_0893_));
 sg13g2_and2_1 _4680_ (.A(_0892_),
    .B(_0894_),
    .X(_0895_));
 sg13g2_nand2_1 _4681_ (.Y(_0896_),
    .A(\vgademo.soundtrack.pulse_osc_p[2] ),
    .B(_0895_));
 sg13g2_xnor2_1 _4682_ (.Y(_0897_),
    .A(net313),
    .B(_0895_));
 sg13g2_nand2b_1 _4683_ (.Y(_0898_),
    .B(_0891_),
    .A_N(_0897_));
 sg13g2_xor2_1 _4684_ (.B(_0897_),
    .A(_0891_),
    .X(_0899_));
 sg13g2_a21oi_1 _4685_ (.A1(net881),
    .A2(_0899_),
    .Y(_0191_),
    .B1(_0890_));
 sg13g2_nand2_1 _4686_ (.Y(_0900_),
    .A(_0868_),
    .B(_0879_));
 sg13g2_nand2_1 _4687_ (.Y(_0901_),
    .A(_0882_),
    .B(_0900_));
 sg13g2_o21ai_1 _4688_ (.B1(_0901_),
    .Y(_0902_),
    .A1(_0850_),
    .A2(_0900_));
 sg13g2_and2_1 _4689_ (.A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .B(_0902_),
    .X(_0903_));
 sg13g2_xnor2_1 _4690_ (.Y(_0904_),
    .A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .B(_0902_));
 sg13g2_a21oi_1 _4691_ (.A1(_0896_),
    .A2(_0898_),
    .Y(_0905_),
    .B1(_0904_));
 sg13g2_and3_1 _4692_ (.X(_0906_),
    .A(_0896_),
    .B(_0898_),
    .C(_0904_));
 sg13g2_nor3_1 _4693_ (.A(net880),
    .B(_0905_),
    .C(_0906_),
    .Y(_0907_));
 sg13g2_a21o_1 _4694_ (.A2(net880),
    .A1(net339),
    .B1(_0907_),
    .X(_0192_));
 sg13g2_nand3_1 _4695_ (.B(_0881_),
    .C(_0893_),
    .A(net309),
    .Y(_0908_));
 sg13g2_nand3_1 _4696_ (.B(_0880_),
    .C(_0894_),
    .A(_3198_),
    .Y(_0909_));
 sg13g2_and2_1 _4697_ (.A(_0908_),
    .B(_0909_),
    .X(_0910_));
 sg13g2_o21ai_1 _4698_ (.B1(_0910_),
    .Y(_0911_),
    .A1(_0903_),
    .A2(_0905_));
 sg13g2_or3_1 _4699_ (.A(_0903_),
    .B(_0905_),
    .C(_0910_),
    .X(_0912_));
 sg13g2_nand3_1 _4700_ (.B(_0911_),
    .C(_0912_),
    .A(net881),
    .Y(_0913_));
 sg13g2_o21ai_1 _4701_ (.B1(_0913_),
    .Y(_0193_),
    .A1(_3198_),
    .A2(net881));
 sg13g2_nand2_1 _4702_ (.Y(_0914_),
    .A(_0892_),
    .B(_0900_));
 sg13g2_nor2_1 _4703_ (.A(_3199_),
    .B(_0914_),
    .Y(_0915_));
 sg13g2_xnor2_1 _4704_ (.Y(_0916_),
    .A(_3199_),
    .B(_0914_));
 sg13g2_a21oi_1 _4705_ (.A1(_0908_),
    .A2(_0911_),
    .Y(_0917_),
    .B1(_0916_));
 sg13g2_nand3_1 _4706_ (.B(_0911_),
    .C(_0916_),
    .A(_0908_),
    .Y(_0918_));
 sg13g2_nand3b_1 _4707_ (.B(_0918_),
    .C(net881),
    .Y(_0919_),
    .A_N(_0917_));
 sg13g2_o21ai_1 _4708_ (.B1(_0919_),
    .Y(_0194_),
    .A1(_3199_),
    .A2(net881));
 sg13g2_xnor2_1 _4709_ (.Y(_0920_),
    .A(_3200_),
    .B(_0849_));
 sg13g2_o21ai_1 _4710_ (.B1(_0920_),
    .Y(_0921_),
    .A1(_0915_),
    .A2(_0917_));
 sg13g2_or3_1 _4711_ (.A(_0915_),
    .B(_0917_),
    .C(_0920_),
    .X(_0922_));
 sg13g2_nand3_1 _4712_ (.B(_0921_),
    .C(_0922_),
    .A(net882),
    .Y(_0923_));
 sg13g2_o21ai_1 _4713_ (.B1(_0923_),
    .Y(_0195_),
    .A1(_3200_),
    .A2(net882));
 sg13g2_nor2_1 _4714_ (.A(net350),
    .B(net881),
    .Y(_0924_));
 sg13g2_nor2_1 _4715_ (.A(\vgademo.soundtrack.pulse_osc_p[7] ),
    .B(_0850_),
    .Y(_0925_));
 sg13g2_o21ai_1 _4716_ (.B1(_0921_),
    .Y(_0926_),
    .A1(_3200_),
    .A2(_0850_));
 sg13g2_a21oi_1 _4717_ (.A1(\vgademo.soundtrack.pulse_osc_p[7] ),
    .A2(_0850_),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_xnor2_1 _4718_ (.Y(_0928_),
    .A(net350),
    .B(_0849_));
 sg13g2_xnor2_1 _4719_ (.Y(_0929_),
    .A(_0926_),
    .B(_0928_));
 sg13g2_a21oi_1 _4720_ (.A1(net881),
    .A2(_0929_),
    .Y(_0196_),
    .B1(_0924_));
 sg13g2_nor3_2 _4721_ (.A(net880),
    .B(_0925_),
    .C(_0927_),
    .Y(_0930_));
 sg13g2_and2_1 _4722_ (.A(net224),
    .B(_0930_),
    .X(_0931_));
 sg13g2_xor2_1 _4723_ (.B(_0930_),
    .A(net224),
    .X(_0197_));
 sg13g2_xor2_1 _4724_ (.B(_0931_),
    .A(net256),
    .X(_0198_));
 sg13g2_and3_2 _4725_ (.X(_0932_),
    .A(net256),
    .B(net194),
    .C(_0931_));
 sg13g2_a21oi_1 _4726_ (.A1(\vgademo.soundtrack.pulse_osc_p[9] ),
    .A2(_0931_),
    .Y(_0933_),
    .B1(net194));
 sg13g2_nor2_1 _4727_ (.A(_0932_),
    .B(net195),
    .Y(_0199_));
 sg13g2_xor2_1 _4728_ (.B(_0932_),
    .A(net257),
    .X(_0200_));
 sg13g2_nand3_1 _4729_ (.B(net257),
    .C(_0932_),
    .A(net508),
    .Y(_0934_));
 sg13g2_a21o_1 _4730_ (.A2(_0932_),
    .A1(net257),
    .B1(net508),
    .X(_0935_));
 sg13g2_and2_1 _4731_ (.A(_0934_),
    .B(_0935_),
    .X(_0201_));
 sg13g2_xnor2_1 _4732_ (.Y(_0202_),
    .A(net251),
    .B(_0934_));
 sg13g2_nor3_1 _4733_ (.A(\vgademo.audio_kick_frames[0] ),
    .B(net867),
    .C(_0700_),
    .Y(_0936_));
 sg13g2_a21o_1 _4734_ (.A2(_0664_),
    .A1(net587),
    .B1(_0936_),
    .X(_0203_));
 sg13g2_nand2b_1 _4735_ (.Y(_0937_),
    .B(_0936_),
    .A_N(net454));
 sg13g2_o21ai_1 _4736_ (.B1(net454),
    .Y(_0938_),
    .A1(\vgademo.audio_kick_frames[0] ),
    .A2(net867));
 sg13g2_nand3_1 _4737_ (.B(_0624_),
    .C(_0681_),
    .A(net877),
    .Y(_0939_));
 sg13g2_nand3_1 _4738_ (.B(_0938_),
    .C(_0939_),
    .A(_0937_),
    .Y(_0204_));
 sg13g2_xor2_1 _4739_ (.B(_0937_),
    .A(net385),
    .X(_0940_));
 sg13g2_nand2_1 _4740_ (.Y(_0205_),
    .A(_0939_),
    .B(net386));
 sg13g2_o21ai_1 _4741_ (.B1(_0791_),
    .Y(_0941_),
    .A1(_3280_),
    .A2(_0630_));
 sg13g2_a21oi_1 _4742_ (.A1(net1055),
    .A2(_3259_),
    .Y(_0942_),
    .B1(_3267_));
 sg13g2_o21ai_1 _4743_ (.B1(_0830_),
    .Y(_0943_),
    .A1(_3269_),
    .A2(_3291_));
 sg13g2_nor3_1 _4744_ (.A(net1060),
    .B(_3258_),
    .C(_3272_),
    .Y(_0944_));
 sg13g2_mux4_1 _4745_ (.S0(_0634_),
    .A0(_0943_),
    .A1(_0944_),
    .A2(_0941_),
    .A3(_0942_),
    .S1(_0642_),
    .X(_0945_));
 sg13g2_xnor2_1 _4746_ (.Y(_0946_),
    .A(_3104_),
    .B(_3253_));
 sg13g2_nand2_1 _4747_ (.Y(_0947_),
    .A(net1062),
    .B(_0946_));
 sg13g2_nand2_1 _4748_ (.Y(_0948_),
    .A(_0635_),
    .B(_0947_));
 sg13g2_nand2_1 _4749_ (.Y(_0949_),
    .A(net1050),
    .B(_3271_));
 sg13g2_a21oi_1 _4750_ (.A1(_0948_),
    .A2(_0949_),
    .Y(_0950_),
    .B1(\vgademo.audio_songpos[6] ));
 sg13g2_or3_1 _4751_ (.A(_0639_),
    .B(_0945_),
    .C(_0950_),
    .X(_0951_));
 sg13g2_nand3_1 _4752_ (.B(_3259_),
    .C(_3297_),
    .A(net960),
    .Y(_0952_));
 sg13g2_o21ai_1 _4753_ (.B1(_0952_),
    .Y(_0953_),
    .A1(_0792_),
    .A2(_0820_));
 sg13g2_nand2_1 _4754_ (.Y(_0954_),
    .A(_3098_),
    .B(_0706_));
 sg13g2_nand4_1 _4755_ (.B(_0946_),
    .C(_0948_),
    .A(_0642_),
    .Y(_0955_),
    .D(_0954_));
 sg13g2_o21ai_1 _4756_ (.B1(_0955_),
    .Y(_0956_),
    .A1(_0642_),
    .A2(_0953_));
 sg13g2_nand2_1 _4757_ (.Y(_0957_),
    .A(_0641_),
    .B(_0947_));
 sg13g2_nand3_1 _4758_ (.B(_0956_),
    .C(_0957_),
    .A(_0639_),
    .Y(_0958_));
 sg13g2_nand3_1 _4759_ (.B(_0951_),
    .C(_0958_),
    .A(_0624_),
    .Y(_0959_));
 sg13g2_and2_2 _4760_ (.A(_0669_),
    .B(_0959_),
    .X(_0960_));
 sg13g2_o21ai_1 _4761_ (.B1(_0625_),
    .Y(_0961_),
    .A1(_3142_),
    .A2(_3336_));
 sg13g2_mux2_1 _4762_ (.A0(net222),
    .A1(_0961_),
    .S(_0960_),
    .X(_0206_));
 sg13g2_o21ai_1 _4763_ (.B1(_0625_),
    .Y(_0962_),
    .A1(_3336_),
    .A2(_3342_));
 sg13g2_mux2_1 _4764_ (.A0(net208),
    .A1(_0962_),
    .S(_0960_),
    .X(_0207_));
 sg13g2_xnor2_1 _4765_ (.Y(_0963_),
    .A(_3143_),
    .B(_3340_));
 sg13g2_o21ai_1 _4766_ (.B1(_0625_),
    .Y(_0964_),
    .A1(_3336_),
    .A2(_0963_));
 sg13g2_mux2_1 _4767_ (.A0(net223),
    .A1(_0964_),
    .S(_0960_),
    .X(_0208_));
 sg13g2_a21oi_1 _4768_ (.A1(\vgademo.soundtrack.pulse_vol[2] ),
    .A2(_3340_),
    .Y(_0965_),
    .B1(net1019));
 sg13g2_o21ai_1 _4769_ (.B1(_0960_),
    .Y(_0966_),
    .A1(_0624_),
    .A2(_0965_));
 sg13g2_o21ai_1 _4770_ (.B1(_0966_),
    .Y(_0209_),
    .A1(_3084_),
    .A2(_0960_));
 sg13g2_nand2_1 _4771_ (.Y(_0967_),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B(net883));
 sg13g2_xnor2_1 _4772_ (.Y(_0210_),
    .A(net206),
    .B(_0967_));
 sg13g2_nand2_1 _4773_ (.Y(_0968_),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B(net206));
 sg13g2_xor2_1 _4774_ (.B(\vgademo.soundtrack.tri_osc_p[1] ),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(_0969_));
 sg13g2_nor2b_1 _4775_ (.A(_0968_),
    .B_N(_0969_),
    .Y(_0970_));
 sg13g2_xor2_1 _4776_ (.B(_0969_),
    .A(_0968_),
    .X(_0971_));
 sg13g2_nand2_1 _4777_ (.Y(_0972_),
    .A(net348),
    .B(_0810_));
 sg13g2_o21ai_1 _4778_ (.B1(_0972_),
    .Y(_0211_),
    .A1(_0810_),
    .A2(_0971_));
 sg13g2_nor2_1 _4779_ (.A(net401),
    .B(net884),
    .Y(_0973_));
 sg13g2_nand2_1 _4780_ (.Y(_0974_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_xnor2_1 _4781_ (.Y(_0975_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_a21oi_1 _4782_ (.A1(\vgademo.soundtrack.tri_osc_i[1] ),
    .A2(net348),
    .Y(_0976_),
    .B1(_0970_));
 sg13g2_or2_1 _4783_ (.X(_0977_),
    .B(_0976_),
    .A(_0975_));
 sg13g2_xnor2_1 _4784_ (.Y(_0978_),
    .A(_0975_),
    .B(_0976_));
 sg13g2_a21oi_1 _4785_ (.A1(net884),
    .A2(_0978_),
    .Y(_0212_),
    .B1(_0973_));
 sg13g2_nor2_1 _4786_ (.A(net397),
    .B(net884),
    .Y(_0979_));
 sg13g2_xnor2_1 _4787_ (.Y(_0980_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_a21oi_1 _4788_ (.A1(_0974_),
    .A2(_0977_),
    .Y(_0981_),
    .B1(_0980_));
 sg13g2_nand3_1 _4789_ (.B(_0977_),
    .C(_0980_),
    .A(_0974_),
    .Y(_0982_));
 sg13g2_nand2b_1 _4790_ (.Y(_0983_),
    .B(_0982_),
    .A_N(_0981_));
 sg13g2_a21oi_1 _4791_ (.A1(net884),
    .A2(_0983_),
    .Y(_0213_),
    .B1(_0979_));
 sg13g2_nor2_1 _4792_ (.A(net421),
    .B(net883),
    .Y(_0984_));
 sg13g2_nand2_1 _4793_ (.Y(_0985_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_xnor2_1 _4794_ (.Y(_0986_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_a21oi_1 _4795_ (.A1(\vgademo.soundtrack.tri_osc_i[3] ),
    .A2(net397),
    .Y(_0987_),
    .B1(_0981_));
 sg13g2_xnor2_1 _4796_ (.Y(_0988_),
    .A(_0986_),
    .B(_0987_));
 sg13g2_a21oi_1 _4797_ (.A1(net884),
    .A2(_0988_),
    .Y(_0214_),
    .B1(_0984_));
 sg13g2_nor2_1 _4798_ (.A(net413),
    .B(net883),
    .Y(_0989_));
 sg13g2_o21ai_1 _4799_ (.B1(_0985_),
    .Y(_0990_),
    .A1(_0986_),
    .A2(_0987_));
 sg13g2_nand2_1 _4800_ (.Y(_0991_),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_xor2_1 _4801_ (.B(net413),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(_0992_));
 sg13g2_xnor2_1 _4802_ (.Y(_0993_),
    .A(_0990_),
    .B(_0992_));
 sg13g2_a21oi_1 _4803_ (.A1(net883),
    .A2(_0993_),
    .Y(_0215_),
    .B1(_0989_));
 sg13g2_nor2_1 _4804_ (.A(_3139_),
    .B(_3196_),
    .Y(_0994_));
 sg13g2_xnor2_1 _4805_ (.Y(_0995_),
    .A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_o21ai_1 _4806_ (.B1(_0990_),
    .Y(_0996_),
    .A1(\vgademo.soundtrack.tri_osc_i[5] ),
    .A2(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_nand3_1 _4807_ (.B(_0995_),
    .C(_0996_),
    .A(_0991_),
    .Y(_0997_));
 sg13g2_a21oi_1 _4808_ (.A1(_0991_),
    .A2(_0996_),
    .Y(_0998_),
    .B1(_0995_));
 sg13g2_nand3b_1 _4809_ (.B(net883),
    .C(_0997_),
    .Y(_0999_),
    .A_N(_0998_));
 sg13g2_o21ai_1 _4810_ (.B1(_0999_),
    .Y(_0216_),
    .A1(_3196_),
    .A2(net883));
 sg13g2_nand2_1 _4811_ (.Y(_1000_),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .B(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_xor2_1 _4812_ (.B(\vgademo.soundtrack.tri_osc_p[7] ),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(_1001_));
 sg13g2_or3_1 _4813_ (.A(_0994_),
    .B(_0998_),
    .C(_1001_),
    .X(_1002_));
 sg13g2_o21ai_1 _4814_ (.B1(_1001_),
    .Y(_1003_),
    .A1(_0994_),
    .A2(_0998_));
 sg13g2_nand3_1 _4815_ (.B(_1002_),
    .C(_1003_),
    .A(net883),
    .Y(_1004_));
 sg13g2_o21ai_1 _4816_ (.B1(_1004_),
    .Y(_0217_),
    .A1(_3195_),
    .A2(net883));
 sg13g2_xnor2_1 _4817_ (.Y(_1005_),
    .A(\vgademo.soundtrack.tri_osc_i[8] ),
    .B(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_and3_1 _4818_ (.X(_1006_),
    .A(_1000_),
    .B(_1003_),
    .C(_1005_));
 sg13g2_a21oi_1 _4819_ (.A1(_1000_),
    .A2(_1003_),
    .Y(_1007_),
    .B1(_1005_));
 sg13g2_nor3_1 _4820_ (.A(net880),
    .B(_1006_),
    .C(_1007_),
    .Y(_1008_));
 sg13g2_a21o_1 _4821_ (.A2(net880),
    .A1(net453),
    .B1(_1008_),
    .X(_0218_));
 sg13g2_a21oi_2 _4822_ (.B1(_1007_),
    .Y(_1009_),
    .A2(\vgademo.soundtrack.tri_osc_p[8] ),
    .A1(\vgademo.soundtrack.tri_osc_i[8] ));
 sg13g2_nor3_2 _4823_ (.A(net371),
    .B(net880),
    .C(_1009_),
    .Y(_1010_));
 sg13g2_nand3_1 _4824_ (.B(net885),
    .C(_1009_),
    .A(net371),
    .Y(_1011_));
 sg13g2_o21ai_1 _4825_ (.B1(_1011_),
    .Y(_1012_),
    .A1(\vgademo.soundtrack.tri_osc_p[9] ),
    .A2(net885));
 sg13g2_nor2_1 _4826_ (.A(net372),
    .B(_1012_),
    .Y(_0219_));
 sg13g2_and2_1 _4827_ (.A(net281),
    .B(_1010_),
    .X(_1013_));
 sg13g2_xor2_1 _4828_ (.B(_1010_),
    .A(net281),
    .X(_0220_));
 sg13g2_xor2_1 _4829_ (.B(_1013_),
    .A(net358),
    .X(_0221_));
 sg13g2_nand3_1 _4830_ (.B(net358),
    .C(_1013_),
    .A(net431),
    .Y(_1014_));
 sg13g2_a21o_1 _4831_ (.A2(_1013_),
    .A1(net358),
    .B1(net431),
    .X(_1015_));
 sg13g2_and2_1 _4832_ (.A(_1014_),
    .B(_1015_),
    .X(_0222_));
 sg13g2_nand4_1 _4833_ (.B(net431),
    .C(net358),
    .A(net305),
    .Y(_1016_),
    .D(_1013_));
 sg13g2_xnor2_1 _4834_ (.Y(_0223_),
    .A(net305),
    .B(_1014_));
 sg13g2_xnor2_1 _4835_ (.Y(_0224_),
    .A(net354),
    .B(_1016_));
 sg13g2_o21ai_1 _4836_ (.B1(net1016),
    .Y(_1017_),
    .A1(_3194_),
    .A2(_1016_));
 sg13g2_o21ai_1 _4837_ (.B1(_1017_),
    .Y(_0225_),
    .A1(_0547_),
    .A2(_1016_));
 sg13g2_or2_1 _4838_ (.X(_1018_),
    .B(net999),
    .A(net996));
 sg13g2_nor2_1 _4839_ (.A(net1001),
    .B(net998),
    .Y(_1019_));
 sg13g2_or3_2 _4840_ (.A(net996),
    .B(net1001),
    .C(net998),
    .X(_1020_));
 sg13g2_nand2_1 _4841_ (.Y(_1021_),
    .A(net992),
    .B(_1020_));
 sg13g2_a21o_1 _4842_ (.A2(_1020_),
    .A1(net992),
    .B1(net991),
    .X(_1022_));
 sg13g2_nor2_1 _4843_ (.A(_3125_),
    .B(net955),
    .Y(_1023_));
 sg13g2_nand2_1 _4844_ (.Y(_1024_),
    .A(net986),
    .B(net987));
 sg13g2_nor3_2 _4845_ (.A(net982),
    .B(net980),
    .C(net983),
    .Y(_1025_));
 sg13g2_nand4_1 _4846_ (.B(net985),
    .C(net987),
    .A(net1003),
    .Y(_1026_),
    .D(_0066_));
 sg13g2_nand2b_1 _4847_ (.Y(_1027_),
    .B(net993),
    .A_N(net990));
 sg13g2_nand2_1 _4848_ (.Y(_1028_),
    .A(net1003),
    .B(_3130_));
 sg13g2_nor3_2 _4849_ (.A(net982),
    .B(\vgademo.a_scrolly[11] ),
    .C(_3131_),
    .Y(_1029_));
 sg13g2_nor4_1 _4850_ (.A(_3123_),
    .B(_1020_),
    .C(_1024_),
    .D(_1027_),
    .Y(_1030_));
 sg13g2_a22oi_1 _4851_ (.Y(_1031_),
    .B1(_1029_),
    .B2(_1030_),
    .A2(_1023_),
    .A1(_1022_));
 sg13g2_and2_1 _4852_ (.A(_1025_),
    .B(_1031_),
    .X(_1032_));
 sg13g2_nor2_2 _4853_ (.A(net990),
    .B(net993),
    .Y(_1033_));
 sg13g2_or2_1 _4854_ (.X(_1034_),
    .B(net993),
    .A(net991));
 sg13g2_nor4_2 _4855_ (.A(net990),
    .B(net992),
    .C(net995),
    .Y(_1035_),
    .D(net998));
 sg13g2_nor2b_1 _4856_ (.A(net1002),
    .B_N(net987),
    .Y(_1036_));
 sg13g2_nand3b_1 _4857_ (.B(net985),
    .C(\vgademo.a_scrolly[11] ),
    .Y(_1037_),
    .A_N(_0065_));
 sg13g2_a21oi_1 _4858_ (.A1(_1035_),
    .A2(_1036_),
    .Y(_1038_),
    .B1(_1037_));
 sg13g2_nand2b_1 _4859_ (.Y(_1039_),
    .B(net983),
    .A_N(net981));
 sg13g2_nor4_2 _4860_ (.A(_1020_),
    .B(_1026_),
    .C(_1034_),
    .Y(_1040_),
    .D(_1039_));
 sg13g2_nor4_2 _4861_ (.A(net981),
    .B(net980),
    .C(_1038_),
    .Y(_1041_),
    .D(_1040_));
 sg13g2_or4_1 _4862_ (.A(net981),
    .B(net980),
    .C(_1038_),
    .D(_1040_),
    .X(_1042_));
 sg13g2_and2_1 _4863_ (.A(net1001),
    .B(net997),
    .X(_1043_));
 sg13g2_nand2_2 _4864_ (.Y(_1044_),
    .A(net1005),
    .B(net1002));
 sg13g2_nand3_1 _4865_ (.B(net1001),
    .C(net997),
    .A(net1003),
    .Y(_1045_));
 sg13g2_nand2_1 _4866_ (.Y(_1046_),
    .A(_3129_),
    .B(_1045_));
 sg13g2_nand2b_1 _4867_ (.Y(_1047_),
    .B(net986),
    .A_N(net987));
 sg13g2_nor2_1 _4868_ (.A(_1027_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_a221oi_1 _4869_ (.B2(_1048_),
    .C1(_1023_),
    .B1(_1046_),
    .A1(net984),
    .Y(_1049_),
    .A2(net990));
 sg13g2_o21ai_1 _4870_ (.B1(_0067_),
    .Y(_1050_),
    .A1(_1039_),
    .A2(_1049_));
 sg13g2_and2_1 _4871_ (.A(_3131_),
    .B(_1050_),
    .X(_1051_));
 sg13g2_nand2_2 _4872_ (.Y(_1052_),
    .A(net981),
    .B(net980));
 sg13g2_nor2_1 _4873_ (.A(_1034_),
    .B(_1047_),
    .Y(_1053_));
 sg13g2_nand4_1 _4874_ (.B(net955),
    .C(_3129_),
    .A(net984),
    .Y(_1054_),
    .D(_1033_));
 sg13g2_nand2_1 _4875_ (.Y(_1055_),
    .A(net985),
    .B(_1054_));
 sg13g2_a221oi_1 _4876_ (.B2(net984),
    .C1(net983),
    .B1(_1054_),
    .A1(_1046_),
    .Y(_1056_),
    .A2(_1053_));
 sg13g2_or2_1 _4877_ (.X(_1057_),
    .B(_1056_),
    .A(_1052_));
 sg13g2_nand3_1 _4878_ (.B(_1050_),
    .C(_1057_),
    .A(_3131_),
    .Y(_1058_));
 sg13g2_a221oi_1 _4879_ (.B2(_1058_),
    .C1(_3132_),
    .B1(net943),
    .A1(_1025_),
    .Y(_1059_),
    .A2(_1031_));
 sg13g2_nand2b_1 _4880_ (.Y(_1060_),
    .B(\vgademo.bayer_j[0] ),
    .A_N(_1059_));
 sg13g2_xnor2_1 _4881_ (.Y(_1061_),
    .A(\vgademo.bayer_j[0] ),
    .B(_1059_));
 sg13g2_nand2b_1 _4882_ (.Y(_1062_),
    .B(_1061_),
    .A_N(\vgademo.audio_kick_frames[0] ));
 sg13g2_xnor2_1 _4883_ (.Y(_1063_),
    .A(\vgademo.audio_kick_frames[0] ),
    .B(_1061_));
 sg13g2_mux2_1 _4884_ (.A0(net427),
    .A1(_1063_),
    .S(net945),
    .X(_0226_));
 sg13g2_a22oi_1 _4885_ (.Y(_1064_),
    .B1(_1041_),
    .B2(_0069_),
    .A2(_1031_),
    .A1(_1025_));
 sg13g2_o21ai_1 _4886_ (.B1(_1064_),
    .Y(_1065_),
    .A1(_3130_),
    .A2(_1041_));
 sg13g2_a21oi_2 _4887_ (.B1(_1065_),
    .Y(_1066_),
    .A2(_1058_),
    .A1(net943));
 sg13g2_xnor2_1 _4888_ (.Y(_1067_),
    .A(\vgademo.bayer_j[1] ),
    .B(_1066_));
 sg13g2_xor2_1 _4889_ (.B(_1067_),
    .A(_0068_),
    .X(_1068_));
 sg13g2_nand2_1 _4890_ (.Y(_1069_),
    .A(_1060_),
    .B(_1062_));
 sg13g2_nand2_1 _4891_ (.Y(_1070_),
    .A(_1068_),
    .B(_1069_));
 sg13g2_xor2_1 _4892_ (.B(_1069_),
    .A(_1068_),
    .X(_1071_));
 sg13g2_and2_1 _4893_ (.A(net945),
    .B(_1071_),
    .X(_1072_));
 sg13g2_a21o_1 _4894_ (.A2(net944),
    .A1(net384),
    .B1(_1072_),
    .X(_0227_));
 sg13g2_nor2_1 _4895_ (.A(_0072_),
    .B(_1066_),
    .Y(_1073_));
 sg13g2_a21oi_1 _4896_ (.A1(_0068_),
    .A2(_1067_),
    .Y(_1074_),
    .B1(_1073_));
 sg13g2_nor2_2 _4897_ (.A(_1019_),
    .B(_1043_),
    .Y(_1075_));
 sg13g2_nand2_1 _4898_ (.Y(_1076_),
    .A(_1041_),
    .B(_1075_));
 sg13g2_nand2b_1 _4899_ (.Y(_1077_),
    .B(net942),
    .A_N(net999));
 sg13g2_a221oi_1 _4900_ (.B2(_1077_),
    .C1(_1032_),
    .B1(_1076_),
    .A1(net943),
    .Y(_1078_),
    .A2(_1058_));
 sg13g2_xnor2_1 _4901_ (.Y(_1079_),
    .A(_0071_),
    .B(_1078_));
 sg13g2_nor2b_1 _4902_ (.A(_1074_),
    .B_N(_1079_),
    .Y(_1080_));
 sg13g2_xor2_1 _4903_ (.B(_1079_),
    .A(_1074_),
    .X(_1081_));
 sg13g2_inv_1 _4904_ (.Y(_1082_),
    .A(_1081_));
 sg13g2_xnor2_1 _4905_ (.Y(_1083_),
    .A(_3108_),
    .B(_1081_));
 sg13g2_nor2_1 _4906_ (.A(_1070_),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_xor2_1 _4907_ (.B(_1083_),
    .A(_1070_),
    .X(_1085_));
 sg13g2_mux2_1 _4908_ (.A0(net289),
    .A1(_1085_),
    .S(net945),
    .X(_0228_));
 sg13g2_nor2_1 _4909_ (.A(net363),
    .B(net945),
    .Y(_1086_));
 sg13g2_and2_1 _4910_ (.A(_3111_),
    .B(_1078_),
    .X(_1087_));
 sg13g2_o21ai_1 _4911_ (.B1(net995),
    .Y(_1088_),
    .A1(net1001),
    .A2(net997));
 sg13g2_a21oi_1 _4912_ (.A1(_1020_),
    .A2(_1088_),
    .Y(_1089_),
    .B1(net942));
 sg13g2_a21o_1 _4913_ (.A2(net943),
    .A1(_0075_),
    .B1(_1089_),
    .X(_1090_));
 sg13g2_a221oi_1 _4914_ (.B2(_1058_),
    .C1(_1090_),
    .B1(net942),
    .A1(_1025_),
    .Y(_1091_),
    .A2(_1031_));
 sg13g2_nand2_1 _4915_ (.Y(_1092_),
    .A(_0074_),
    .B(_1091_));
 sg13g2_xor2_1 _4916_ (.B(_1091_),
    .A(_0074_),
    .X(_1093_));
 sg13g2_xnor2_1 _4917_ (.Y(_1094_),
    .A(_0074_),
    .B(_1091_));
 sg13g2_nand2b_1 _4918_ (.Y(_1095_),
    .B(_1094_),
    .A_N(_1087_));
 sg13g2_xnor2_1 _4919_ (.Y(_1096_),
    .A(_1087_),
    .B(_1094_));
 sg13g2_a21oi_1 _4920_ (.A1(_0060_),
    .A2(_1082_),
    .Y(_1097_),
    .B1(_1080_));
 sg13g2_nor2b_1 _4921_ (.A(_1097_),
    .B_N(_1096_),
    .Y(_1098_));
 sg13g2_xnor2_1 _4922_ (.Y(_1099_),
    .A(_1096_),
    .B(_1097_));
 sg13g2_xnor2_1 _4923_ (.Y(_1100_),
    .A(_1084_),
    .B(_1099_));
 sg13g2_a21oi_1 _4924_ (.A1(net945),
    .A2(_1100_),
    .Y(_0229_),
    .B1(_1086_));
 sg13g2_a21oi_1 _4925_ (.A1(_1084_),
    .A2(_1099_),
    .Y(_1101_),
    .B1(_1098_));
 sg13g2_nor2_1 _4926_ (.A(net992),
    .B(net995),
    .Y(_1102_));
 sg13g2_nor2_1 _4927_ (.A(_3128_),
    .B(_3129_),
    .Y(_1103_));
 sg13g2_nor2_1 _4928_ (.A(_1102_),
    .B(_1103_),
    .Y(_1104_));
 sg13g2_o21ai_1 _4929_ (.B1(_1104_),
    .Y(_1105_),
    .A1(_1052_),
    .A2(_1056_));
 sg13g2_nand4_1 _4930_ (.B(net942),
    .C(_1050_),
    .A(_3131_),
    .Y(_1106_),
    .D(_1105_));
 sg13g2_or2_1 _4931_ (.X(_1107_),
    .B(_1018_),
    .A(_3133_));
 sg13g2_xnor2_1 _4932_ (.Y(_1108_),
    .A(_0078_),
    .B(_1107_));
 sg13g2_a21oi_2 _4933_ (.B1(_1032_),
    .Y(_1109_),
    .A2(_1108_),
    .A1(_1041_));
 sg13g2_and2_1 _4934_ (.A(_1106_),
    .B(_1109_),
    .X(_1110_));
 sg13g2_nand2_1 _4935_ (.Y(_1111_),
    .A(_0077_),
    .B(_1110_));
 sg13g2_xnor2_1 _4936_ (.Y(_1112_),
    .A(_0077_),
    .B(_1110_));
 sg13g2_nand2_1 _4937_ (.Y(_1113_),
    .A(_1092_),
    .B(_1112_));
 sg13g2_xor2_1 _4938_ (.B(_1112_),
    .A(_1092_),
    .X(_1114_));
 sg13g2_nand2b_1 _4939_ (.Y(_1115_),
    .B(_1114_),
    .A_N(_1095_));
 sg13g2_xnor2_1 _4940_ (.Y(_1116_),
    .A(_1095_),
    .B(_1114_));
 sg13g2_inv_1 _4941_ (.Y(_1117_),
    .A(_1116_));
 sg13g2_xnor2_1 _4942_ (.Y(_1118_),
    .A(_1101_),
    .B(_1116_));
 sg13g2_mux2_1 _4943_ (.A0(net298),
    .A1(_1118_),
    .S(net946),
    .X(_0230_));
 sg13g2_nor2_1 _4944_ (.A(net370),
    .B(net946),
    .Y(_1119_));
 sg13g2_o21ai_1 _4945_ (.B1(_1115_),
    .Y(_1120_),
    .A1(_1101_),
    .A2(_1117_));
 sg13g2_inv_1 _4946_ (.Y(_1121_),
    .A(_1120_));
 sg13g2_xor2_1 _4947_ (.B(_1102_),
    .A(_0080_),
    .X(_1122_));
 sg13g2_o21ai_1 _4948_ (.B1(_1122_),
    .Y(_1123_),
    .A1(_1052_),
    .A2(_1056_));
 sg13g2_nand4_1 _4949_ (.B(net942),
    .C(_1050_),
    .A(_3131_),
    .Y(_1124_),
    .D(_1123_));
 sg13g2_nand2_1 _4950_ (.Y(_1125_),
    .A(net993),
    .B(_1107_));
 sg13g2_a21oi_1 _4951_ (.A1(_0080_),
    .A2(_1125_),
    .Y(_1126_),
    .B1(net943));
 sg13g2_o21ai_1 _4952_ (.B1(_1126_),
    .Y(_1127_),
    .A1(_0080_),
    .A2(_1125_));
 sg13g2_a21oi_2 _4953_ (.B1(_1032_),
    .Y(_1128_),
    .A2(_1127_),
    .A1(_1124_));
 sg13g2_nand2_1 _4954_ (.Y(_1129_),
    .A(net977),
    .B(_1128_));
 sg13g2_xnor2_1 _4955_ (.Y(_1130_),
    .A(net977),
    .B(_1128_));
 sg13g2_or2_1 _4956_ (.X(_1131_),
    .B(_1130_),
    .A(_1111_));
 sg13g2_xnor2_1 _4957_ (.Y(_1132_),
    .A(_1111_),
    .B(_1130_));
 sg13g2_nand2b_1 _4958_ (.Y(_1133_),
    .B(_1132_),
    .A_N(_1113_));
 sg13g2_xor2_1 _4959_ (.B(_1132_),
    .A(_1113_),
    .X(_1134_));
 sg13g2_xor2_1 _4960_ (.B(_1134_),
    .A(_1120_),
    .X(_1135_));
 sg13g2_a21oi_1 _4961_ (.A1(net946),
    .A2(_1135_),
    .Y(_0231_),
    .B1(_1119_));
 sg13g2_nor2_1 _4962_ (.A(net301),
    .B(net946),
    .Y(_1136_));
 sg13g2_o21ai_1 _4963_ (.B1(_1133_),
    .Y(_1137_),
    .A1(_1121_),
    .A2(_1134_));
 sg13g2_nand2b_1 _4964_ (.Y(_1138_),
    .B(_0063_),
    .A_N(_1128_));
 sg13g2_nand2_1 _4965_ (.Y(_1139_),
    .A(_0075_),
    .B(_1033_));
 sg13g2_nand3_1 _4966_ (.B(_0075_),
    .C(_1033_),
    .A(net955),
    .Y(_1140_));
 sg13g2_xnor2_1 _4967_ (.Y(_1141_),
    .A(net955),
    .B(_1139_));
 sg13g2_o21ai_1 _4968_ (.B1(_1141_),
    .Y(_1142_),
    .A1(_1052_),
    .A2(_1056_));
 sg13g2_nand4_1 _4969_ (.B(net942),
    .C(_1050_),
    .A(_3131_),
    .Y(_1143_),
    .D(_1142_));
 sg13g2_nand3_1 _4970_ (.B(net993),
    .C(_1107_),
    .A(\vgademo.a_scrolly[8] ),
    .Y(_1144_));
 sg13g2_xnor2_1 _4971_ (.Y(_1145_),
    .A(net955),
    .B(_1144_));
 sg13g2_nand2_1 _4972_ (.Y(_1146_),
    .A(_1041_),
    .B(_1145_));
 sg13g2_a21o_1 _4973_ (.A2(_1146_),
    .A1(_1143_),
    .B1(_1032_),
    .X(_1147_));
 sg13g2_xor2_1 _4974_ (.B(_1147_),
    .A(net975),
    .X(_1148_));
 sg13g2_nand2_1 _4975_ (.Y(_1149_),
    .A(_1138_),
    .B(_1148_));
 sg13g2_xor2_1 _4976_ (.B(_1148_),
    .A(_1138_),
    .X(_1150_));
 sg13g2_xnor2_1 _4977_ (.Y(_1151_),
    .A(_1131_),
    .B(_1150_));
 sg13g2_nor2b_1 _4978_ (.A(_1151_),
    .B_N(_1137_),
    .Y(_1152_));
 sg13g2_xor2_1 _4979_ (.B(_1151_),
    .A(_1137_),
    .X(_1153_));
 sg13g2_a21oi_1 _4980_ (.A1(net946),
    .A2(_1153_),
    .Y(_0232_),
    .B1(_1136_));
 sg13g2_a21o_1 _4981_ (.A2(_1150_),
    .A1(_1131_),
    .B1(_1152_),
    .X(_1154_));
 sg13g2_xor2_1 _4982_ (.B(_1140_),
    .A(_0015_),
    .X(_1155_));
 sg13g2_o21ai_1 _4983_ (.B1(_1155_),
    .Y(_1156_),
    .A1(_1052_),
    .A2(_1056_));
 sg13g2_nand3_1 _4984_ (.B(_1050_),
    .C(_1156_),
    .A(_3131_),
    .Y(_1157_));
 sg13g2_a21oi_1 _4985_ (.A1(_0065_),
    .A2(_1144_),
    .Y(_1158_),
    .B1(net985));
 sg13g2_and3_1 _4986_ (.X(_1159_),
    .A(net984),
    .B(_0065_),
    .C(_1144_));
 sg13g2_nor3_1 _4987_ (.A(net942),
    .B(_1158_),
    .C(_1159_),
    .Y(_1160_));
 sg13g2_a221oi_1 _4988_ (.B2(_1157_),
    .C1(_1160_),
    .B1(net942),
    .A1(_1025_),
    .Y(_1161_),
    .A2(_1031_));
 sg13g2_nand2b_1 _4989_ (.Y(_1162_),
    .B(_0014_),
    .A_N(_1161_));
 sg13g2_xnor2_1 _4990_ (.Y(_1163_),
    .A(_0014_),
    .B(_1161_));
 sg13g2_and2_1 _4991_ (.A(_0016_),
    .B(_1147_),
    .X(_1164_));
 sg13g2_nor2_1 _4992_ (.A(_1163_),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_xnor2_1 _4993_ (.Y(_1166_),
    .A(_1163_),
    .B(_1164_));
 sg13g2_nor2_1 _4994_ (.A(_1149_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_xor2_1 _4995_ (.B(_1166_),
    .A(_1149_),
    .X(_1168_));
 sg13g2_xor2_1 _4996_ (.B(_1168_),
    .A(_1154_),
    .X(_1169_));
 sg13g2_mux2_1 _4997_ (.A0(net285),
    .A1(_1169_),
    .S(_0645_),
    .X(_0233_));
 sg13g2_a21oi_1 _4998_ (.A1(_1154_),
    .A2(_1168_),
    .Y(_1170_),
    .B1(_1167_));
 sg13g2_a21oi_1 _4999_ (.A1(net955),
    .A2(_1144_),
    .Y(_1171_),
    .B1(_3125_));
 sg13g2_nand2_1 _5000_ (.Y(_1172_),
    .A(net983),
    .B(_1171_));
 sg13g2_xnor2_1 _5001_ (.Y(_1173_),
    .A(_0019_),
    .B(_1055_));
 sg13g2_nor3_1 _5002_ (.A(_1041_),
    .B(_1058_),
    .C(_1173_),
    .Y(_1174_));
 sg13g2_a21oi_2 _5003_ (.B1(_1174_),
    .Y(_1175_),
    .A2(_1172_),
    .A1(_1041_));
 sg13g2_xnor2_1 _5004_ (.Y(_1176_),
    .A(_3135_),
    .B(_1175_));
 sg13g2_xnor2_1 _5005_ (.Y(_1177_),
    .A(_1162_),
    .B(_1176_));
 sg13g2_xnor2_1 _5006_ (.Y(_1178_),
    .A(_1165_),
    .B(_1177_));
 sg13g2_xnor2_1 _5007_ (.Y(_1179_),
    .A(_1170_),
    .B(_1178_));
 sg13g2_and2_1 _5008_ (.A(_0645_),
    .B(_1179_),
    .X(_1180_));
 sg13g2_a21o_1 _5009_ (.A2(net944),
    .A1(net307),
    .B1(_1180_),
    .X(_0234_));
 sg13g2_nor2_1 _5010_ (.A(net1003),
    .B(net1001),
    .Y(_1181_));
 sg13g2_nand2_1 _5011_ (.Y(_1182_),
    .A(_3123_),
    .B(_3130_));
 sg13g2_nor2_1 _5012_ (.A(net984),
    .B(net988),
    .Y(_1183_));
 sg13g2_nand2_1 _5013_ (.Y(_1184_),
    .A(_3125_),
    .B(net955));
 sg13g2_nor2_1 _5014_ (.A(_3129_),
    .B(_1181_),
    .Y(_1185_));
 sg13g2_nand2_2 _5015_ (.Y(_1186_),
    .A(net996),
    .B(net999));
 sg13g2_nor2b_1 _5016_ (.A(_1185_),
    .B_N(_1029_),
    .Y(_1187_));
 sg13g2_nand4_1 _5017_ (.B(_1183_),
    .C(_1186_),
    .A(_1033_),
    .Y(_1188_),
    .D(_1187_));
 sg13g2_nor3_1 _5018_ (.A(\vgademo.audio_songpos[6] ),
    .B(net1045),
    .C(_3263_),
    .Y(_1189_));
 sg13g2_nand4_1 _5019_ (.B(net954),
    .C(_1188_),
    .A(_3268_),
    .Y(_1190_),
    .D(_1189_));
 sg13g2_nand2_1 _5020_ (.Y(_1191_),
    .A(net925),
    .B(_1190_));
 sg13g2_a21oi_1 _5021_ (.A1(net925),
    .A2(_1190_),
    .Y(_1192_),
    .B1(net1005));
 sg13g2_a21oi_1 _5022_ (.A1(net1005),
    .A2(net925),
    .Y(_0235_),
    .B1(_1192_));
 sg13g2_nand2_1 _5023_ (.Y(_1193_),
    .A(net1002),
    .B(net917));
 sg13g2_nand2_1 _5024_ (.Y(_1194_),
    .A(_1044_),
    .B(_1182_));
 sg13g2_o21ai_1 _5025_ (.B1(_1193_),
    .Y(_0236_),
    .A1(net890),
    .A2(_1194_));
 sg13g2_nand2_1 _5026_ (.Y(_1195_),
    .A(net1000),
    .B(net921));
 sg13g2_xor2_1 _5027_ (.B(_1044_),
    .A(net999),
    .X(_1196_));
 sg13g2_o21ai_1 _5028_ (.B1(_1195_),
    .Y(_0237_),
    .A1(_1191_),
    .A2(_1196_));
 sg13g2_nand2_1 _5029_ (.Y(_1197_),
    .A(net995),
    .B(net917));
 sg13g2_xnor2_1 _5030_ (.Y(_1198_),
    .A(net588),
    .B(_1045_));
 sg13g2_o21ai_1 _5031_ (.B1(_1197_),
    .Y(_0238_),
    .A1(net890),
    .A2(_1198_));
 sg13g2_nand2_1 _5032_ (.Y(_1199_),
    .A(net994),
    .B(net917));
 sg13g2_xor2_1 _5033_ (.B(_1186_),
    .A(_0078_),
    .X(_1200_));
 sg13g2_nand2_1 _5034_ (.Y(_1201_),
    .A(_0078_),
    .B(_1044_));
 sg13g2_o21ai_1 _5035_ (.B1(_1201_),
    .Y(_1202_),
    .A1(_1044_),
    .A2(_1200_));
 sg13g2_o21ai_1 _5036_ (.B1(_1199_),
    .Y(_0239_),
    .A1(_1191_),
    .A2(_1202_));
 sg13g2_nand2_1 _5037_ (.Y(_1203_),
    .A(net318),
    .B(net917));
 sg13g2_nor3_1 _5038_ (.A(_0078_),
    .B(_1044_),
    .C(_1186_),
    .Y(_1204_));
 sg13g2_xor2_1 _5039_ (.B(_1204_),
    .A(_0080_),
    .X(_1205_));
 sg13g2_o21ai_1 _5040_ (.B1(_1203_),
    .Y(_0240_),
    .A1(net890),
    .A2(_1205_));
 sg13g2_nand2_1 _5041_ (.Y(_1206_),
    .A(net987),
    .B(net921));
 sg13g2_nand4_1 _5042_ (.B(net990),
    .C(_1043_),
    .A(net1003),
    .Y(_1207_),
    .D(_1103_));
 sg13g2_nor2_1 _5043_ (.A(_0065_),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_xnor2_1 _5044_ (.Y(_1209_),
    .A(net525),
    .B(_1207_));
 sg13g2_o21ai_1 _5045_ (.B1(_1206_),
    .Y(_0241_),
    .A1(net890),
    .A2(_1209_));
 sg13g2_nand2_1 _5046_ (.Y(_1210_),
    .A(net986),
    .B(net917));
 sg13g2_xor2_1 _5047_ (.B(_1208_),
    .A(net442),
    .X(_1211_));
 sg13g2_o21ai_1 _5048_ (.B1(_1210_),
    .Y(_0242_),
    .A1(net890),
    .A2(net443));
 sg13g2_nand2_1 _5049_ (.Y(_1212_),
    .A(net983),
    .B(net917));
 sg13g2_nor2_2 _5050_ (.A(_1024_),
    .B(_1207_),
    .Y(_1213_));
 sg13g2_nand2b_1 _5051_ (.Y(_1214_),
    .B(_1213_),
    .A_N(net448));
 sg13g2_xor2_1 _5052_ (.B(_1213_),
    .A(net448),
    .X(_1215_));
 sg13g2_o21ai_1 _5053_ (.B1(_1212_),
    .Y(_0243_),
    .A1(net890),
    .A2(_1215_));
 sg13g2_nand2_1 _5054_ (.Y(_1216_),
    .A(net981),
    .B(net917));
 sg13g2_xnor2_1 _5055_ (.Y(_1217_),
    .A(_0067_),
    .B(_1214_));
 sg13g2_o21ai_1 _5056_ (.B1(_1216_),
    .Y(_0244_),
    .A1(net890),
    .A2(net449));
 sg13g2_nand2_1 _5057_ (.Y(_1218_),
    .A(net980),
    .B(net917));
 sg13g2_nand3_1 _5058_ (.B(net551),
    .C(_1213_),
    .A(net981),
    .Y(_1219_));
 sg13g2_xnor2_1 _5059_ (.Y(_1220_),
    .A(net568),
    .B(_1219_));
 sg13g2_o21ai_1 _5060_ (.B1(_1218_),
    .Y(_0245_),
    .A1(net890),
    .A2(_1220_));
 sg13g2_nand2_2 _5061_ (.Y(_1221_),
    .A(_3211_),
    .B(_0589_));
 sg13g2_a21oi_1 _5062_ (.A1(_3211_),
    .A2(_0589_),
    .Y(_1222_),
    .B1(net979));
 sg13g2_nand2_1 _5063_ (.Y(_1223_),
    .A(net979),
    .B(_3211_));
 sg13g2_nor2b_1 _5064_ (.A(_1222_),
    .B_N(_1223_),
    .Y(_0246_));
 sg13g2_xnor2_1 _5065_ (.Y(_0247_),
    .A(net589),
    .B(_1223_));
 sg13g2_nand2_1 _5066_ (.Y(_1224_),
    .A(\vgademo.v_count[2] ),
    .B(net949));
 sg13g2_nand2_2 _5067_ (.Y(_1225_),
    .A(\vgademo.bayer_j[1] ),
    .B(net979));
 sg13g2_nor2_1 _5068_ (.A(net470),
    .B(_1225_),
    .Y(_1226_));
 sg13g2_xnor2_1 _5069_ (.Y(_1227_),
    .A(net470),
    .B(_1225_));
 sg13g2_o21ai_1 _5070_ (.B1(_1224_),
    .Y(_0248_),
    .A1(_1221_),
    .A2(_1227_));
 sg13g2_nand2_1 _5071_ (.Y(_1228_),
    .A(net473),
    .B(net949));
 sg13g2_xor2_1 _5072_ (.B(_1226_),
    .A(_0074_),
    .X(_1229_));
 sg13g2_o21ai_1 _5073_ (.B1(_1228_),
    .Y(_0249_),
    .A1(_1221_),
    .A2(_1229_));
 sg13g2_nand2_1 _5074_ (.Y(_1230_),
    .A(net302),
    .B(net949));
 sg13g2_nor2_1 _5075_ (.A(_3236_),
    .B(_1225_),
    .Y(_1231_));
 sg13g2_nor3_1 _5076_ (.A(_0077_),
    .B(_3236_),
    .C(_1225_),
    .Y(_1232_));
 sg13g2_xor2_1 _5077_ (.B(_1231_),
    .A(_0077_),
    .X(_1233_));
 sg13g2_o21ai_1 _5078_ (.B1(_1230_),
    .Y(_0250_),
    .A1(_1221_),
    .A2(_1233_));
 sg13g2_nand2_1 _5079_ (.Y(_1234_),
    .A(net977),
    .B(net949));
 sg13g2_xor2_1 _5080_ (.B(_1232_),
    .A(net489),
    .X(_1235_));
 sg13g2_o21ai_1 _5081_ (.B1(_1234_),
    .Y(_0251_),
    .A1(_1221_),
    .A2(_1235_));
 sg13g2_nand2_1 _5082_ (.Y(_1236_),
    .A(net975),
    .B(net948));
 sg13g2_nand3_1 _5083_ (.B(net976),
    .C(_1231_),
    .A(net302),
    .Y(_1237_));
 sg13g2_nor2_1 _5084_ (.A(_0016_),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_xnor2_1 _5085_ (.Y(_1239_),
    .A(_0016_),
    .B(_1237_));
 sg13g2_o21ai_1 _5086_ (.B1(_1236_),
    .Y(_0252_),
    .A1(_1221_),
    .A2(_1239_));
 sg13g2_nand2_1 _5087_ (.Y(_1240_),
    .A(net287),
    .B(net948));
 sg13g2_xor2_1 _5088_ (.B(_1238_),
    .A(_0014_),
    .X(_1241_));
 sg13g2_o21ai_1 _5089_ (.B1(_1240_),
    .Y(_0253_),
    .A1(_1221_),
    .A2(_1241_));
 sg13g2_nand2_1 _5090_ (.Y(_1242_),
    .A(\vgademo.v_count[8] ),
    .B(net948));
 sg13g2_o21ai_1 _5091_ (.B1(net522),
    .Y(_1243_),
    .A1(_3234_),
    .A2(_1237_));
 sg13g2_nor3_2 _5092_ (.A(net522),
    .B(_3234_),
    .C(_1237_),
    .Y(_1244_));
 sg13g2_nand2b_1 _5093_ (.Y(_1245_),
    .B(net523),
    .A_N(_1221_));
 sg13g2_o21ai_1 _5094_ (.B1(_1242_),
    .Y(_0254_),
    .A1(_1244_),
    .A2(_1245_));
 sg13g2_nand2_1 _5095_ (.Y(_1246_),
    .A(net973),
    .B(net948));
 sg13g2_xor2_1 _5096_ (.B(_1244_),
    .A(net437),
    .X(_1247_));
 sg13g2_o21ai_1 _5097_ (.B1(_1246_),
    .Y(_0255_),
    .A1(_1221_),
    .A2(net438));
 sg13g2_o21ai_1 _5098_ (.B1(_0037_),
    .Y(_1248_),
    .A1(net957),
    .A2(\vgademo.scanline_audio_sample[5] ));
 sg13g2_xor2_1 _5099_ (.B(\vgademo.scanline_audio_sample[6] ),
    .A(net1008),
    .X(_1249_));
 sg13g2_nor2_1 _5100_ (.A(_1248_),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_nand2_1 _5101_ (.Y(_1251_),
    .A(net957),
    .B(\vgademo.scanline_audio_sample[5] ));
 sg13g2_o21ai_1 _5102_ (.B1(_1251_),
    .Y(_1252_),
    .A1(net1009),
    .A2(_3201_));
 sg13g2_a21oi_1 _5103_ (.A1(net1009),
    .A2(_3201_),
    .Y(_1253_),
    .B1(_1252_));
 sg13g2_and2_1 _5104_ (.A(_1250_),
    .B(_1253_),
    .X(_1254_));
 sg13g2_nand2_1 _5105_ (.Y(_1255_),
    .A(_3117_),
    .B(\vgademo.scanline_audio_sample[2] ));
 sg13g2_xor2_1 _5106_ (.B(\vgademo.scanline_audio_sample[2] ),
    .A(net1012),
    .X(_1256_));
 sg13g2_nor2b_1 _5107_ (.A(\vgademo.scanline_audio_sample[3] ),
    .B_N(net1010),
    .Y(_1257_));
 sg13g2_nand2b_1 _5108_ (.Y(_1258_),
    .B(\vgademo.scanline_audio_sample[3] ),
    .A_N(net1010));
 sg13g2_nor2b_1 _5109_ (.A(_1257_),
    .B_N(_1258_),
    .Y(_1259_));
 sg13g2_nand2_1 _5110_ (.Y(_1260_),
    .A(_1254_),
    .B(_1259_));
 sg13g2_nor2_1 _5111_ (.A(_1256_),
    .B(_1260_),
    .Y(_1261_));
 sg13g2_nor2b_1 _5112_ (.A(net1014),
    .B_N(\vgademo.scanline_audio_sample[1] ),
    .Y(_1262_));
 sg13g2_nand2_1 _5113_ (.Y(_1263_),
    .A(_3114_),
    .B(\vgademo.scanline_audio_sample[1] ));
 sg13g2_nor2_1 _5114_ (.A(_3115_),
    .B(\vgademo.scanline_audio_sample[0] ),
    .Y(_1264_));
 sg13g2_nor2_1 _5115_ (.A(_3114_),
    .B(\vgademo.scanline_audio_sample[1] ),
    .Y(_1265_));
 sg13g2_o21ai_1 _5116_ (.B1(_1263_),
    .Y(_1266_),
    .A1(_1264_),
    .A2(_1265_));
 sg13g2_nor2_1 _5117_ (.A(\vgademo.h_count[7] ),
    .B(net1008),
    .Y(_1267_));
 sg13g2_a22oi_1 _5118_ (.Y(_1268_),
    .B1(_1267_),
    .B2(\vgademo.scanline_audio_sample[6] ),
    .A2(_1252_),
    .A1(_1250_));
 sg13g2_a21oi_1 _5119_ (.A1(_1255_),
    .A2(_1258_),
    .Y(_1269_),
    .B1(_1257_));
 sg13g2_a22oi_1 _5120_ (.Y(_1270_),
    .B1(_1269_),
    .B2(_1254_),
    .A2(_1266_),
    .A1(_1261_));
 sg13g2_nor2b_1 _5121_ (.A(\vgademo.h_count[0] ),
    .B_N(\vgademo.scanline_audio_sample[0] ),
    .Y(_1271_));
 sg13g2_nor4_2 _5122_ (.A(_1262_),
    .B(_1264_),
    .C(_1265_),
    .Y(_1272_),
    .D(_1271_));
 sg13g2_nand2_1 _5123_ (.Y(_1273_),
    .A(net1006),
    .B(_0579_));
 sg13g2_a221oi_1 _5124_ (.B2(_1261_),
    .C1(_1273_),
    .B1(_1272_),
    .A1(_1268_),
    .Y(_1274_),
    .A2(_1270_));
 sg13g2_inv_2 _5125_ (.Y(_1275_),
    .A(_1274_));
 sg13g2_nor2_1 _5126_ (.A(\vgademo.scanline_audio_sample[4] ),
    .B(\vgademo.scanline_audio_sample[3] ),
    .Y(_1276_));
 sg13g2_nand2_1 _5127_ (.Y(_1277_),
    .A(_0043_),
    .B(_1276_));
 sg13g2_xor2_1 _5128_ (.B(_1277_),
    .A(\vgademo.scanline_audio_sample[6] ),
    .X(_1278_));
 sg13g2_xnor2_1 _5129_ (.Y(_1279_),
    .A(_0036_),
    .B(_1278_));
 sg13g2_nand2_1 _5130_ (.Y(_1280_),
    .A(_0037_),
    .B(_1279_));
 sg13g2_xnor2_1 _5131_ (.Y(_1281_),
    .A(_0043_),
    .B(_1276_));
 sg13g2_xnor2_1 _5132_ (.Y(_1282_),
    .A(_0035_),
    .B(_1281_));
 sg13g2_xnor2_1 _5133_ (.Y(_1283_),
    .A(\vgademo.scanline_audio_sample[4] ),
    .B(\vgademo.scanline_audio_sample[3] ));
 sg13g2_nand2_1 _5134_ (.Y(_1284_),
    .A(_0044_),
    .B(_1283_));
 sg13g2_xnor2_1 _5135_ (.Y(_1285_),
    .A(_0044_),
    .B(_1283_));
 sg13g2_nor3_1 _5136_ (.A(_1280_),
    .B(_1282_),
    .C(_1285_),
    .Y(_1286_));
 sg13g2_nor2_1 _5137_ (.A(_1256_),
    .B(_1259_),
    .Y(_1287_));
 sg13g2_nor2_1 _5138_ (.A(net1010),
    .B(\vgademo.scanline_audio_sample[3] ),
    .Y(_1288_));
 sg13g2_a21oi_1 _5139_ (.A1(_1266_),
    .A2(_1287_),
    .Y(_1289_),
    .B1(_1288_));
 sg13g2_o21ai_1 _5140_ (.B1(_1289_),
    .Y(_1290_),
    .A1(_1255_),
    .A2(_1259_));
 sg13g2_nor2b_1 _5141_ (.A(_1278_),
    .B_N(_1267_),
    .Y(_1291_));
 sg13g2_nand2_1 _5142_ (.Y(_1292_),
    .A(net957),
    .B(_1281_));
 sg13g2_o21ai_1 _5143_ (.B1(_1292_),
    .Y(_1293_),
    .A1(_1282_),
    .A2(_1284_));
 sg13g2_nor2b_1 _5144_ (.A(_1280_),
    .B_N(_1293_),
    .Y(_1294_));
 sg13g2_a21o_1 _5145_ (.A2(_1290_),
    .A1(_1286_),
    .B1(_1294_),
    .X(_1295_));
 sg13g2_nand3_1 _5146_ (.B(_1286_),
    .C(_1287_),
    .A(_1272_),
    .Y(_1296_));
 sg13g2_o21ai_1 _5147_ (.B1(_1296_),
    .Y(_1297_),
    .A1(_1291_),
    .A2(_1295_));
 sg13g2_nor2_2 _5148_ (.A(_1275_),
    .B(_1297_),
    .Y(_1298_));
 sg13g2_nor2_2 _5149_ (.A(\vgademo.v_count[8] ),
    .B(net973),
    .Y(_1299_));
 sg13g2_nand2b_1 _5150_ (.Y(_1300_),
    .B(_1299_),
    .A_N(_1175_));
 sg13g2_inv_1 _5151_ (.Y(_1301_),
    .A(_1300_));
 sg13g2_nand2b_1 _5152_ (.Y(_1302_),
    .B(_1163_),
    .A_N(_1148_));
 sg13g2_nor3_1 _5153_ (.A(_1112_),
    .B(_1130_),
    .C(_1302_),
    .Y(_1303_));
 sg13g2_xnor2_1 _5154_ (.Y(_1304_),
    .A(\vgademo.v_count[2] ),
    .B(_1078_));
 sg13g2_and2_1 _5155_ (.A(_1093_),
    .B(_1304_),
    .X(_1305_));
 sg13g2_nand2_1 _5156_ (.Y(_1306_),
    .A(_1093_),
    .B(_1304_));
 sg13g2_a22oi_1 _5157_ (.Y(_1307_),
    .B1(_1067_),
    .B2(_1060_),
    .A2(_1066_),
    .A1(_0072_));
 sg13g2_a22oi_1 _5158_ (.Y(_1308_),
    .B1(_1093_),
    .B2(_1087_),
    .A2(_1091_),
    .A1(_3110_));
 sg13g2_o21ai_1 _5159_ (.B1(_1308_),
    .Y(_1309_),
    .A1(_1306_),
    .A2(_1307_));
 sg13g2_nor2_1 _5160_ (.A(net974),
    .B(_1161_),
    .Y(_1310_));
 sg13g2_a21oi_1 _5161_ (.A1(_1163_),
    .A2(_1164_),
    .Y(_1311_),
    .B1(_1310_));
 sg13g2_nand3_1 _5162_ (.B(_1106_),
    .C(_1109_),
    .A(_3112_),
    .Y(_1312_));
 sg13g2_o21ai_1 _5163_ (.B1(_1312_),
    .Y(_1313_),
    .A1(net977),
    .A2(_1128_));
 sg13g2_nand2_1 _5164_ (.Y(_1314_),
    .A(_1129_),
    .B(_1313_));
 sg13g2_o21ai_1 _5165_ (.B1(_1311_),
    .Y(_1315_),
    .A1(_1302_),
    .A2(_1314_));
 sg13g2_a21o_1 _5166_ (.A2(_1309_),
    .A1(_1303_),
    .B1(_1315_),
    .X(_1316_));
 sg13g2_nor2_1 _5167_ (.A(net973),
    .B(_1176_),
    .Y(_1317_));
 sg13g2_a21o_2 _5168_ (.A2(_1317_),
    .A1(_1316_),
    .B1(_1301_),
    .X(_1318_));
 sg13g2_and2_1 _5169_ (.A(_1061_),
    .B(_1317_),
    .X(_1319_));
 sg13g2_nand4_1 _5170_ (.B(_1303_),
    .C(_1305_),
    .A(_1067_),
    .Y(_1320_),
    .D(_1319_));
 sg13g2_nand2_1 _5171_ (.Y(_1321_),
    .A(_1318_),
    .B(_1320_));
 sg13g2_inv_1 _5172_ (.Y(_1322_),
    .A(net872));
 sg13g2_mux2_1 _5173_ (.A0(_0071_),
    .A1(_0049_),
    .S(net876),
    .X(_1323_));
 sg13g2_nor2_1 _5174_ (.A(\vgademo.b_cos[7] ),
    .B(_1323_),
    .Y(_1324_));
 sg13g2_xnor2_1 _5175_ (.Y(_1325_),
    .A(_3156_),
    .B(_1323_));
 sg13g2_nor2b_1 _5176_ (.A(net979),
    .B_N(\vgademo.b_cos[5] ),
    .Y(_1326_));
 sg13g2_nor2_1 _5177_ (.A(\vgademo.b_cos[6] ),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_a21oi_1 _5178_ (.A1(\vgademo.b_cos[6] ),
    .A2(_1326_),
    .Y(_1328_),
    .B1(_0072_));
 sg13g2_nor2_1 _5179_ (.A(_1327_),
    .B(_1328_),
    .Y(_1329_));
 sg13g2_nor2b_2 _5180_ (.A(\vgademo.plane_du[2] ),
    .B_N(\vgademo.b_cos[5] ),
    .Y(_1330_));
 sg13g2_nand2_1 _5181_ (.Y(_1331_),
    .A(net971),
    .B(_1330_));
 sg13g2_nor2_1 _5182_ (.A(net971),
    .B(_1330_),
    .Y(_1332_));
 sg13g2_o21ai_1 _5183_ (.B1(_1331_),
    .Y(_1333_),
    .A1(_3202_),
    .A2(_1332_));
 sg13g2_mux2_1 _5184_ (.A0(_1329_),
    .A1(_1333_),
    .S(net876),
    .X(_1334_));
 sg13g2_inv_1 _5185_ (.Y(_1335_),
    .A(_1334_));
 sg13g2_a21oi_1 _5186_ (.A1(_1325_),
    .A2(_1335_),
    .Y(_1336_),
    .B1(_1324_));
 sg13g2_mux2_1 _5187_ (.A0(_0074_),
    .A1(_0051_),
    .S(net876),
    .X(_1337_));
 sg13g2_nor2_1 _5188_ (.A(\vgademo.b_cos[8] ),
    .B(_1337_),
    .Y(_1338_));
 sg13g2_xnor2_1 _5189_ (.Y(_1339_),
    .A(_3157_),
    .B(_1337_));
 sg13g2_nor2b_1 _5190_ (.A(_1336_),
    .B_N(_1339_),
    .Y(_1340_));
 sg13g2_xnor2_1 _5191_ (.Y(_1341_),
    .A(_1336_),
    .B(_1339_));
 sg13g2_inv_1 _5192_ (.Y(_1342_),
    .A(_1341_));
 sg13g2_nand2_1 _5193_ (.Y(_1343_),
    .A(net991),
    .B(_3128_));
 sg13g2_nor4_2 _5194_ (.A(net984),
    .B(net956),
    .C(net996),
    .Y(_1344_),
    .D(_1343_));
 sg13g2_nand2_2 _5195_ (.Y(_1345_),
    .A(net999),
    .B(_1182_));
 sg13g2_a22oi_1 _5196_ (.Y(_1346_),
    .B1(_1344_),
    .B2(_1345_),
    .A2(_0080_),
    .A1(_3125_));
 sg13g2_nand4_1 _5197_ (.B(_1029_),
    .C(_1181_),
    .A(net998),
    .Y(_1347_),
    .D(_1344_));
 sg13g2_nand2_1 _5198_ (.Y(_1348_),
    .A(_1025_),
    .B(_1347_));
 sg13g2_a21oi_2 _5199_ (.B1(_1348_),
    .Y(_1349_),
    .A2(_1346_),
    .A1(_1184_));
 sg13g2_a21oi_1 _5200_ (.A1(net988),
    .A2(_1022_),
    .Y(_1350_),
    .B1(net984));
 sg13g2_nand2_1 _5201_ (.Y(_1351_),
    .A(net980),
    .B(net983));
 sg13g2_o21ai_1 _5202_ (.B1(_1052_),
    .Y(_1352_),
    .A1(_1350_),
    .A2(_1351_));
 sg13g2_a21o_2 _5203_ (.A2(_1352_),
    .A1(_1051_),
    .B1(_1349_),
    .X(_1353_));
 sg13g2_inv_1 _5204_ (.Y(_1354_),
    .A(_1353_));
 sg13g2_nor2_1 _5205_ (.A(_1047_),
    .B(_1343_),
    .Y(_1355_));
 sg13g2_nand4_1 _5206_ (.B(net995),
    .C(_1019_),
    .A(net1003),
    .Y(_1356_),
    .D(_1355_));
 sg13g2_a221oi_1 _5207_ (.B2(_1355_),
    .C1(_3125_),
    .B1(_1088_),
    .A1(net955),
    .Y(_1357_),
    .A2(_3127_));
 sg13g2_nand2_1 _5208_ (.Y(_1358_),
    .A(_1025_),
    .B(_1356_));
 sg13g2_nor2_2 _5209_ (.A(_1357_),
    .B(_1358_),
    .Y(_1359_));
 sg13g2_nand2_1 _5210_ (.Y(_1360_),
    .A(_1018_),
    .B(_1186_));
 sg13g2_xor2_1 _5211_ (.B(_1345_),
    .A(_0075_),
    .X(_1361_));
 sg13g2_a221oi_1 _5212_ (.B2(_1352_),
    .C1(_1353_),
    .B1(_1361_),
    .A1(_1359_),
    .Y(_1362_),
    .A2(_1360_));
 sg13g2_nor3_1 _5213_ (.A(net1014),
    .B(net1010),
    .C(net1012),
    .Y(_1363_));
 sg13g2_and2_1 _5214_ (.A(_3119_),
    .B(_1363_),
    .X(_1364_));
 sg13g2_nor2_1 _5215_ (.A(net957),
    .B(_1364_),
    .Y(_1365_));
 sg13g2_nand2_1 _5216_ (.Y(_1366_),
    .A(net1008),
    .B(_1365_));
 sg13g2_inv_1 _5217_ (.Y(_1367_),
    .A(_1366_));
 sg13g2_xnor2_1 _5218_ (.Y(_1368_),
    .A(_3120_),
    .B(_1366_));
 sg13g2_nor2_1 _5219_ (.A(net875),
    .B(_1368_),
    .Y(_1369_));
 sg13g2_a21oi_2 _5220_ (.B1(_1369_),
    .Y(_1370_),
    .A2(net875),
    .A1(_0046_));
 sg13g2_nand2_2 _5221_ (.Y(_1371_),
    .A(_1362_),
    .B(_1370_));
 sg13g2_xor2_1 _5222_ (.B(_1181_),
    .A(net997),
    .X(_1372_));
 sg13g2_a221oi_1 _5223_ (.B2(_1352_),
    .C1(_1353_),
    .B1(_1372_),
    .A1(net999),
    .Y(_1373_),
    .A2(_1359_));
 sg13g2_xnor2_1 _5224_ (.Y(_1374_),
    .A(_0036_),
    .B(_1365_));
 sg13g2_nand2_1 _5225_ (.Y(_1375_),
    .A(_0030_),
    .B(net875));
 sg13g2_o21ai_1 _5226_ (.B1(_1375_),
    .Y(_1376_),
    .A1(net875),
    .A2(_1374_));
 sg13g2_nor2b_1 _5227_ (.A(_1376_),
    .B_N(_1373_),
    .Y(_1377_));
 sg13g2_nand2b_1 _5228_ (.Y(_1378_),
    .B(_1373_),
    .A_N(_1376_));
 sg13g2_nor2b_2 _5229_ (.A(_1051_),
    .B_N(_1352_),
    .Y(_1379_));
 sg13g2_a22oi_1 _5230_ (.Y(_1380_),
    .B1(_1379_),
    .B2(_1194_),
    .A2(_1359_),
    .A1(_3133_));
 sg13g2_or2_2 _5231_ (.X(_1381_),
    .B(_1380_),
    .A(_1349_));
 sg13g2_xnor2_1 _5232_ (.Y(_1382_),
    .A(net957),
    .B(_1364_));
 sg13g2_mux2_2 _5233_ (.A0(_1382_),
    .A1(_0047_),
    .S(net875),
    .X(_1383_));
 sg13g2_nor2_1 _5234_ (.A(_1381_),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_or2_1 _5235_ (.X(_1385_),
    .B(_1383_),
    .A(_1381_));
 sg13g2_a221oi_1 _5236_ (.B2(_0064_),
    .C1(_1353_),
    .B1(_1359_),
    .A1(net1005),
    .Y(_1386_),
    .A2(_1352_));
 sg13g2_xnor2_1 _5237_ (.Y(_1387_),
    .A(_0044_),
    .B(_1363_));
 sg13g2_a21oi_1 _5238_ (.A1(_1318_),
    .A2(_1320_),
    .Y(_1388_),
    .B1(_0029_));
 sg13g2_and3_1 _5239_ (.X(_1389_),
    .A(_1318_),
    .B(_1320_),
    .C(_1387_));
 sg13g2_o21ai_1 _5240_ (.B1(_1386_),
    .Y(_1390_),
    .A1(_1388_),
    .A2(_1389_));
 sg13g2_or3_1 _5241_ (.A(_1386_),
    .B(_1388_),
    .C(_1389_),
    .X(_1391_));
 sg13g2_a21o_1 _5242_ (.A2(_1320_),
    .A1(_1318_),
    .B1(_0048_),
    .X(_1392_));
 sg13g2_xnor2_1 _5243_ (.Y(_1393_),
    .A(_0034_),
    .B(_3243_));
 sg13g2_nand3_1 _5244_ (.B(_1320_),
    .C(_1393_),
    .A(_1318_),
    .Y(_1394_));
 sg13g2_and2_1 _5245_ (.A(_1392_),
    .B(_1394_),
    .X(_1395_));
 sg13g2_xnor2_1 _5246_ (.Y(_1396_),
    .A(net1015),
    .B(net1013));
 sg13g2_a21o_1 _5247_ (.A2(_1320_),
    .A1(_1318_),
    .B1(_0028_),
    .X(_1397_));
 sg13g2_nand3_1 _5248_ (.B(_1320_),
    .C(_1396_),
    .A(_1318_),
    .Y(_1398_));
 sg13g2_nand4_1 _5249_ (.B(_1394_),
    .C(_1397_),
    .A(_1392_),
    .Y(_1399_),
    .D(_1398_));
 sg13g2_and4_1 _5250_ (.A(_1354_),
    .B(_1390_),
    .C(_1391_),
    .D(_1399_),
    .X(_1400_));
 sg13g2_nand4_1 _5251_ (.B(_1390_),
    .C(_1391_),
    .A(_1354_),
    .Y(_1401_),
    .D(_1399_));
 sg13g2_xnor2_1 _5252_ (.Y(_1402_),
    .A(_1381_),
    .B(_1383_));
 sg13g2_a21oi_2 _5253_ (.B1(_1402_),
    .Y(_1403_),
    .A2(_1401_),
    .A1(_1390_));
 sg13g2_a21o_2 _5254_ (.A2(_1401_),
    .A1(_1390_),
    .B1(_1402_),
    .X(_1404_));
 sg13g2_xnor2_1 _5255_ (.Y(_1405_),
    .A(_1373_),
    .B(_1376_));
 sg13g2_xor2_1 _5256_ (.B(_1376_),
    .A(_1373_),
    .X(_1406_));
 sg13g2_a21oi_2 _5257_ (.B1(_1406_),
    .Y(_1407_),
    .A2(_1404_),
    .A1(_1385_));
 sg13g2_o21ai_1 _5258_ (.B1(_1405_),
    .Y(_1408_),
    .A1(_1384_),
    .A2(_1403_));
 sg13g2_xor2_1 _5259_ (.B(_1370_),
    .A(_1362_),
    .X(_1409_));
 sg13g2_xnor2_1 _5260_ (.Y(_1410_),
    .A(_1362_),
    .B(_1370_));
 sg13g2_o21ai_1 _5261_ (.B1(_1409_),
    .Y(_1411_),
    .A1(_1377_),
    .A2(net860));
 sg13g2_nand3_1 _5262_ (.B(_1028_),
    .C(_1075_),
    .A(_0075_),
    .Y(_1412_));
 sg13g2_xnor2_1 _5263_ (.Y(_1413_),
    .A(net992),
    .B(_1020_));
 sg13g2_nor2b_1 _5264_ (.A(_1412_),
    .B_N(_1413_),
    .Y(_1414_));
 sg13g2_xnor2_1 _5265_ (.Y(_1415_),
    .A(_1412_),
    .B(_1413_));
 sg13g2_a221oi_1 _5266_ (.B2(_1352_),
    .C1(_1353_),
    .B1(_1415_),
    .A1(_1200_),
    .Y(_1416_),
    .A2(_1359_));
 sg13g2_nand2_1 _5267_ (.Y(_1417_),
    .A(_0037_),
    .B(_1366_));
 sg13g2_xor2_1 _5268_ (.B(_1417_),
    .A(_0038_),
    .X(_1418_));
 sg13g2_nand2_1 _5269_ (.Y(_1419_),
    .A(_0031_),
    .B(net874));
 sg13g2_o21ai_1 _5270_ (.B1(_1419_),
    .Y(_1420_),
    .A1(net874),
    .A2(_1418_));
 sg13g2_nand2b_1 _5271_ (.Y(_1421_),
    .B(_1416_),
    .A_N(_1420_));
 sg13g2_inv_1 _5272_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_xnor2_1 _5273_ (.Y(_1423_),
    .A(_1416_),
    .B(_1420_));
 sg13g2_xor2_1 _5274_ (.B(_1420_),
    .A(_1416_),
    .X(_1424_));
 sg13g2_a21oi_1 _5275_ (.A1(_1371_),
    .A2(net854),
    .Y(_1425_),
    .B1(_1424_));
 sg13g2_a21o_1 _5276_ (.A2(net854),
    .A1(_1371_),
    .B1(_1424_),
    .X(_1426_));
 sg13g2_and3_2 _5277_ (.X(_1427_),
    .A(_1371_),
    .B(net854),
    .C(_1424_));
 sg13g2_nand3_1 _5278_ (.B(net854),
    .C(_1424_),
    .A(_1371_),
    .Y(_1428_));
 sg13g2_a21oi_2 _5279_ (.B1(_1423_),
    .Y(_1429_),
    .A2(net854),
    .A1(_1371_));
 sg13g2_and3_2 _5280_ (.X(_1430_),
    .A(_1371_),
    .B(net854),
    .C(_1423_));
 sg13g2_nor2_1 _5281_ (.A(net848),
    .B(_1427_),
    .Y(_1431_));
 sg13g2_nand2_2 _5282_ (.Y(_1432_),
    .A(net845),
    .B(net842));
 sg13g2_xnor2_1 _5283_ (.Y(_1433_),
    .A(_1325_),
    .B(_1334_));
 sg13g2_xnor2_1 _5284_ (.Y(_1434_),
    .A(_1325_),
    .B(_1335_));
 sg13g2_a21oi_2 _5285_ (.B1(net864),
    .Y(_1435_),
    .A2(net842),
    .A1(net845));
 sg13g2_o21ai_1 _5286_ (.B1(net865),
    .Y(_1436_),
    .A1(net847),
    .A2(net844));
 sg13g2_nor3_1 _5287_ (.A(_1384_),
    .B(_1403_),
    .C(_1405_),
    .Y(_1437_));
 sg13g2_nand3_1 _5288_ (.B(_1404_),
    .C(_1406_),
    .A(_1385_),
    .Y(_1438_));
 sg13g2_nand3_1 _5289_ (.B(_1404_),
    .C(_1405_),
    .A(_1385_),
    .Y(_1439_));
 sg13g2_o21ai_1 _5290_ (.B1(_1406_),
    .Y(_1440_),
    .A1(_1384_),
    .A2(_1403_));
 sg13g2_nor2_2 _5291_ (.A(_1407_),
    .B(net858),
    .Y(_1441_));
 sg13g2_nand2_2 _5292_ (.Y(_1442_),
    .A(_1408_),
    .B(_1438_));
 sg13g2_a22oi_1 _5293_ (.Y(_1443_),
    .B1(_1399_),
    .B2(_1354_),
    .A2(_1391_),
    .A1(_1390_));
 sg13g2_nor2_2 _5294_ (.A(_1400_),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_or2_1 _5295_ (.X(_1445_),
    .B(_1443_),
    .A(_1400_));
 sg13g2_and3_1 _5296_ (.X(_1446_),
    .A(_1390_),
    .B(_1401_),
    .C(_1402_));
 sg13g2_nand3_1 _5297_ (.B(_1401_),
    .C(_1402_),
    .A(_1390_),
    .Y(_1447_));
 sg13g2_nor2_1 _5298_ (.A(_1403_),
    .B(_1446_),
    .Y(_1448_));
 sg13g2_nand2_1 _5299_ (.Y(_1449_),
    .A(_1404_),
    .B(_1447_));
 sg13g2_a21oi_2 _5300_ (.B1(_1444_),
    .Y(_1450_),
    .A2(_1447_),
    .A1(_1404_));
 sg13g2_o21ai_1 _5301_ (.B1(net862),
    .Y(_1451_),
    .A1(_1403_),
    .A2(_1446_));
 sg13g2_nor3_2 _5302_ (.A(_1407_),
    .B(net858),
    .C(_1450_),
    .Y(_1452_));
 sg13g2_nand3_1 _5303_ (.B(_1397_),
    .C(_1398_),
    .A(_1354_),
    .Y(_1453_));
 sg13g2_xor2_1 _5304_ (.B(_1453_),
    .A(_1395_),
    .X(_1454_));
 sg13g2_xnor2_1 _5305_ (.Y(_1455_),
    .A(_1395_),
    .B(_1453_));
 sg13g2_nand2_2 _5306_ (.Y(_1456_),
    .A(_1445_),
    .B(_1455_));
 sg13g2_a22oi_1 _5307_ (.Y(_1457_),
    .B1(_1448_),
    .B2(_1456_),
    .A2(_1438_),
    .A1(_1408_));
 sg13g2_a21o_1 _5308_ (.A2(_1456_),
    .A1(net857),
    .B1(_1441_),
    .X(_1458_));
 sg13g2_nor2_2 _5309_ (.A(_1452_),
    .B(_1457_),
    .Y(_1459_));
 sg13g2_or2_1 _5310_ (.X(_1460_),
    .B(_1457_),
    .A(_1452_));
 sg13g2_nand3_1 _5311_ (.B(net859),
    .C(_1410_),
    .A(_1378_),
    .Y(_1461_));
 sg13g2_o21ai_1 _5312_ (.B1(_1410_),
    .Y(_1462_),
    .A1(_1377_),
    .A2(net860));
 sg13g2_nand3_1 _5313_ (.B(net859),
    .C(_1409_),
    .A(_1378_),
    .Y(_1463_));
 sg13g2_nand2_1 _5314_ (.Y(_1464_),
    .A(_1462_),
    .B(_1463_));
 sg13g2_nand2_1 _5315_ (.Y(_1465_),
    .A(net853),
    .B(net852));
 sg13g2_nor3_2 _5316_ (.A(net847),
    .B(net844),
    .C(net840),
    .Y(_1466_));
 sg13g2_nor4_2 _5317_ (.A(net848),
    .B(_1427_),
    .C(_1459_),
    .Y(_1467_),
    .D(net840));
 sg13g2_nand2_1 _5318_ (.Y(_1468_),
    .A(_1460_),
    .B(_1466_));
 sg13g2_nor3_2 _5319_ (.A(_1400_),
    .B(_1443_),
    .C(_1455_),
    .Y(_1469_));
 sg13g2_nand2_2 _5320_ (.Y(_1470_),
    .A(_1444_),
    .B(_1454_));
 sg13g2_xnor2_1 _5321_ (.Y(_1471_),
    .A(_1445_),
    .B(_1454_));
 sg13g2_nor2b_1 _5322_ (.A(_1471_),
    .B_N(_1452_),
    .Y(_1472_));
 sg13g2_or4_2 _5323_ (.A(net860),
    .B(net858),
    .C(_1450_),
    .D(_1471_),
    .X(_1473_));
 sg13g2_nor2_2 _5324_ (.A(net862),
    .B(net857),
    .Y(_1474_));
 sg13g2_nand2_1 _5325_ (.Y(_1475_),
    .A(_1444_),
    .B(_1449_));
 sg13g2_nand2_1 _5326_ (.Y(_1476_),
    .A(_1442_),
    .B(_1474_));
 sg13g2_a21oi_1 _5327_ (.A1(_1473_),
    .A2(_1476_),
    .Y(_1477_),
    .B1(_1465_));
 sg13g2_a221oi_1 _5328_ (.B2(_1476_),
    .C1(net839),
    .B1(_1473_),
    .A1(net845),
    .Y(_1478_),
    .A2(net842));
 sg13g2_a21oi_2 _5329_ (.B1(net840),
    .Y(_1479_),
    .A2(net842),
    .A1(net846));
 sg13g2_nor3_2 _5330_ (.A(_1407_),
    .B(_1437_),
    .C(net856),
    .Y(_1480_));
 sg13g2_nand2_1 _5331_ (.Y(_1481_),
    .A(_1444_),
    .B(_1480_));
 sg13g2_nor4_2 _5332_ (.A(net860),
    .B(net858),
    .C(net856),
    .Y(_1482_),
    .D(_1470_));
 sg13g2_nand2_1 _5333_ (.Y(_1483_),
    .A(_1469_),
    .B(_1480_));
 sg13g2_nor3_1 _5334_ (.A(_1441_),
    .B(_1454_),
    .C(_1475_),
    .Y(_1484_));
 sg13g2_nand3_1 _5335_ (.B(_1455_),
    .C(_1474_),
    .A(_1442_),
    .Y(_1485_));
 sg13g2_nand2_1 _5336_ (.Y(_1486_),
    .A(_1483_),
    .B(_1485_));
 sg13g2_a21oi_1 _5337_ (.A1(_1479_),
    .A2(_1486_),
    .Y(_1487_),
    .B1(_1478_));
 sg13g2_a21oi_1 _5338_ (.A1(_1468_),
    .A2(_1487_),
    .Y(_1488_),
    .B1(_1435_));
 sg13g2_a21oi_1 _5339_ (.A1(_1481_),
    .A2(_1485_),
    .Y(_1489_),
    .B1(net840));
 sg13g2_o21ai_1 _5340_ (.B1(_1435_),
    .Y(_1490_),
    .A1(_1477_),
    .A2(_1489_));
 sg13g2_o21ai_1 _5341_ (.B1(_1490_),
    .Y(_1491_),
    .A1(_1432_),
    .A2(_1473_));
 sg13g2_o21ai_1 _5342_ (.B1(net861),
    .Y(_1492_),
    .A1(_1488_),
    .A2(_1491_));
 sg13g2_nand4_1 _5343_ (.B(_1440_),
    .C(net856),
    .A(_1439_),
    .Y(_1493_),
    .D(_1470_));
 sg13g2_nand3_1 _5344_ (.B(_1461_),
    .C(_1493_),
    .A(net854),
    .Y(_1494_));
 sg13g2_nand4_1 _5345_ (.B(_1461_),
    .C(_1473_),
    .A(net853),
    .Y(_1495_),
    .D(_1493_));
 sg13g2_and3_1 _5346_ (.X(_1496_),
    .A(net845),
    .B(net843),
    .C(_1495_));
 sg13g2_o21ai_1 _5347_ (.B1(_1496_),
    .Y(_1497_),
    .A1(_1460_),
    .A2(net840));
 sg13g2_o21ai_1 _5348_ (.B1(_1497_),
    .Y(_1498_),
    .A1(net864),
    .A2(_1487_));
 sg13g2_xor2_1 _5349_ (.B(_1021_),
    .A(_0080_),
    .X(_1499_));
 sg13g2_nand2_1 _5350_ (.Y(_1500_),
    .A(_1414_),
    .B(_1499_));
 sg13g2_or2_1 _5351_ (.X(_1501_),
    .B(_1499_),
    .A(_1414_));
 sg13g2_nand3_1 _5352_ (.B(_1500_),
    .C(_1501_),
    .A(_1379_),
    .Y(_1502_));
 sg13g2_nand3_1 _5353_ (.B(_1018_),
    .C(_1186_),
    .A(_0078_),
    .Y(_1503_));
 sg13g2_or2_1 _5354_ (.X(_1504_),
    .B(_1503_),
    .A(_3127_));
 sg13g2_o21ai_1 _5355_ (.B1(net991),
    .Y(_1505_),
    .A1(net993),
    .A2(_1018_));
 sg13g2_nand3b_1 _5356_ (.B(_1503_),
    .C(_1505_),
    .Y(_1506_),
    .A_N(_1035_));
 sg13g2_nand3_1 _5357_ (.B(_1504_),
    .C(_1506_),
    .A(_1359_),
    .Y(_1507_));
 sg13g2_a21o_1 _5358_ (.A2(_1507_),
    .A1(_1502_),
    .B1(_1349_),
    .X(_1508_));
 sg13g2_nor3_1 _5359_ (.A(\vgademo.h_count[7] ),
    .B(net1007),
    .C(_1367_),
    .Y(_1509_));
 sg13g2_nor2_1 _5360_ (.A(_3121_),
    .B(_1509_),
    .Y(_1510_));
 sg13g2_inv_1 _5361_ (.Y(_1511_),
    .A(_1510_));
 sg13g2_xnor2_1 _5362_ (.Y(_1512_),
    .A(\vgademo.h_count[9] ),
    .B(_1509_));
 sg13g2_nand2_1 _5363_ (.Y(_1513_),
    .A(_0045_),
    .B(net874));
 sg13g2_o21ai_1 _5364_ (.B1(_1513_),
    .Y(_1514_),
    .A1(net874),
    .A2(_1512_));
 sg13g2_nor2_1 _5365_ (.A(_1508_),
    .B(_1514_),
    .Y(_1515_));
 sg13g2_xor2_1 _5366_ (.B(_1514_),
    .A(_1508_),
    .X(_1516_));
 sg13g2_inv_1 _5367_ (.Y(_1517_),
    .A(_1516_));
 sg13g2_a21oi_2 _5368_ (.B1(_1517_),
    .Y(_1518_),
    .A2(net846),
    .A1(_1421_));
 sg13g2_o21ai_1 _5369_ (.B1(_1516_),
    .Y(_1519_),
    .A1(_1422_),
    .A2(net847));
 sg13g2_nor3_2 _5370_ (.A(_1422_),
    .B(net847),
    .C(_1516_),
    .Y(_1520_));
 sg13g2_nand3_1 _5371_ (.B(net846),
    .C(_1517_),
    .A(_1421_),
    .Y(_1521_));
 sg13g2_nor2_2 _5372_ (.A(_1518_),
    .B(_1520_),
    .Y(_1522_));
 sg13g2_nand2_2 _5373_ (.Y(_1523_),
    .A(_1519_),
    .B(_1521_));
 sg13g2_nor2_2 _5374_ (.A(net861),
    .B(_1433_),
    .Y(_1524_));
 sg13g2_nand2_1 _5375_ (.Y(_1525_),
    .A(_1342_),
    .B(net864));
 sg13g2_o21ai_1 _5376_ (.B1(net862),
    .Y(_1526_),
    .A1(net860),
    .A2(net858));
 sg13g2_nand3_1 _5377_ (.B(_1438_),
    .C(_1471_),
    .A(net859),
    .Y(_1527_));
 sg13g2_nand4_1 _5378_ (.B(net852),
    .C(_1526_),
    .A(net853),
    .Y(_1528_),
    .D(_1527_));
 sg13g2_a21oi_2 _5379_ (.B1(_1528_),
    .Y(_1529_),
    .A2(net843),
    .A1(_1426_));
 sg13g2_a21oi_2 _5380_ (.B1(_1451_),
    .Y(_1530_),
    .A2(_1438_),
    .A1(net859));
 sg13g2_o21ai_1 _5381_ (.B1(_1450_),
    .Y(_1531_),
    .A1(net860),
    .A2(net858));
 sg13g2_nand4_1 _5382_ (.B(_1438_),
    .C(net857),
    .A(net859),
    .Y(_1532_),
    .D(_1470_));
 sg13g2_and2_1 _5383_ (.A(_1531_),
    .B(_1532_),
    .X(_1533_));
 sg13g2_a221oi_1 _5384_ (.B2(_1480_),
    .C1(_1530_),
    .B1(_1470_),
    .A1(net853),
    .Y(_1534_),
    .A2(net852));
 sg13g2_a221oi_1 _5385_ (.B2(_1479_),
    .C1(_1529_),
    .B1(_1533_),
    .A1(_1431_),
    .Y(_1535_),
    .A2(_1495_));
 sg13g2_o21ai_1 _5386_ (.B1(_1522_),
    .Y(_1536_),
    .A1(_1525_),
    .A2(_1535_));
 sg13g2_a21oi_1 _5387_ (.A1(net855),
    .A2(_1498_),
    .Y(_1537_),
    .B1(_1536_));
 sg13g2_nor2_1 _5388_ (.A(_1338_),
    .B(_1340_),
    .Y(_1538_));
 sg13g2_mux2_1 _5389_ (.A0(_0077_),
    .A1(_0052_),
    .S(net875),
    .X(_1539_));
 sg13g2_xnor2_1 _5390_ (.Y(_1540_),
    .A(_3158_),
    .B(_1539_));
 sg13g2_o21ai_1 _5391_ (.B1(_1540_),
    .Y(_1541_),
    .A1(_1338_),
    .A2(_1340_));
 sg13g2_xnor2_1 _5392_ (.Y(_1542_),
    .A(_1538_),
    .B(_1540_));
 sg13g2_inv_2 _5393_ (.Y(_1543_),
    .A(_1542_));
 sg13g2_nor4_1 _5394_ (.A(_1432_),
    .B(net856),
    .C(net840),
    .D(_1470_),
    .Y(_1544_));
 sg13g2_nor3_2 _5395_ (.A(net848),
    .B(net844),
    .C(net839),
    .Y(_1545_));
 sg13g2_nand3_1 _5396_ (.B(net842),
    .C(net840),
    .A(net845),
    .Y(_1546_));
 sg13g2_nand2b_1 _5397_ (.Y(_1547_),
    .B(_1480_),
    .A_N(_1471_));
 sg13g2_a21oi_1 _5398_ (.A1(_1485_),
    .A2(_1547_),
    .Y(_1548_),
    .B1(_1546_));
 sg13g2_or2_1 _5399_ (.X(_1549_),
    .B(_1548_),
    .A(_1544_));
 sg13g2_and2_1 _5400_ (.A(_1456_),
    .B(_1480_),
    .X(_1550_));
 sg13g2_nand2_2 _5401_ (.Y(_1551_),
    .A(net857),
    .B(_1471_));
 sg13g2_o21ai_1 _5402_ (.B1(_1531_),
    .Y(_1552_),
    .A1(_1442_),
    .A2(_1551_));
 sg13g2_nor4_2 _5403_ (.A(net848),
    .B(net844),
    .C(net839),
    .Y(_1553_),
    .D(_1552_));
 sg13g2_a21oi_1 _5404_ (.A1(_1442_),
    .A2(_1551_),
    .Y(_1554_),
    .B1(_1452_));
 sg13g2_a21o_1 _5405_ (.A2(_1551_),
    .A1(_1442_),
    .B1(_1452_),
    .X(_1555_));
 sg13g2_nor4_1 _5406_ (.A(net847),
    .B(_1427_),
    .C(net841),
    .D(_1554_),
    .Y(_1556_));
 sg13g2_o21ai_1 _5407_ (.B1(_1524_),
    .Y(_1557_),
    .A1(_1553_),
    .A2(_1556_));
 sg13g2_a21oi_1 _5408_ (.A1(net845),
    .A2(net842),
    .Y(_1558_),
    .B1(_1554_));
 sg13g2_a221oi_1 _5409_ (.B2(_1432_),
    .C1(_1522_),
    .B1(_1555_),
    .A1(_1525_),
    .Y(_1559_),
    .A2(_1549_));
 sg13g2_a221oi_1 _5410_ (.B2(_1559_),
    .C1(_1542_),
    .B1(_1557_),
    .A1(_1492_),
    .Y(_1560_),
    .A2(_1537_));
 sg13g2_mux2_1 _5411_ (.A0(_0063_),
    .A1(_0053_),
    .S(net875),
    .X(_1561_));
 sg13g2_xnor2_1 _5412_ (.Y(_1562_),
    .A(net970),
    .B(_1561_));
 sg13g2_o21ai_1 _5413_ (.B1(_1541_),
    .Y(_1563_),
    .A1(\vgademo.b_cos[9] ),
    .A2(_1539_));
 sg13g2_nand2_1 _5414_ (.Y(_1564_),
    .A(_1562_),
    .B(_1563_));
 sg13g2_xor2_1 _5415_ (.B(_1563_),
    .A(_1562_),
    .X(_1565_));
 sg13g2_and2_1 _5416_ (.A(_1452_),
    .B(_1551_),
    .X(_1566_));
 sg13g2_nor2b_1 _5417_ (.A(_1479_),
    .B_N(_1566_),
    .Y(_1567_));
 sg13g2_nor2_1 _5418_ (.A(_1441_),
    .B(_1450_),
    .Y(_1568_));
 sg13g2_o21ai_1 _5419_ (.B1(_1451_),
    .Y(_1569_),
    .A1(net860),
    .A2(net858));
 sg13g2_a22oi_1 _5420_ (.Y(_1570_),
    .B1(_1462_),
    .B2(_1463_),
    .A2(_1456_),
    .A1(net857));
 sg13g2_nand2_1 _5421_ (.Y(_1571_),
    .A(_1568_),
    .B(_1570_));
 sg13g2_o21ai_1 _5422_ (.B1(net839),
    .Y(_1572_),
    .A1(_1484_),
    .A2(_1550_));
 sg13g2_a21oi_1 _5423_ (.A1(_1571_),
    .A2(_1572_),
    .Y(_1573_),
    .B1(_1431_));
 sg13g2_nor4_1 _5424_ (.A(net865),
    .B(_1467_),
    .C(_1567_),
    .D(_1573_),
    .Y(_1574_));
 sg13g2_a22oi_1 _5425_ (.Y(_1575_),
    .B1(_1531_),
    .B2(_1532_),
    .A2(_1463_),
    .A1(_1462_));
 sg13g2_nor3_2 _5426_ (.A(net847),
    .B(net844),
    .C(_1575_),
    .Y(_1576_));
 sg13g2_a221oi_1 _5427_ (.B2(_1442_),
    .C1(_1452_),
    .B1(_1551_),
    .A1(_1411_),
    .Y(_1577_),
    .A2(_1461_));
 sg13g2_nor4_1 _5428_ (.A(net847),
    .B(net844),
    .C(_1575_),
    .D(_1577_),
    .Y(_1578_));
 sg13g2_nor3_2 _5429_ (.A(net847),
    .B(net844),
    .C(net863),
    .Y(_1579_));
 sg13g2_nand4_1 _5430_ (.B(net852),
    .C(_1493_),
    .A(_1411_),
    .Y(_1580_),
    .D(_1532_));
 sg13g2_nor2_1 _5431_ (.A(net862),
    .B(_1454_),
    .Y(_1581_));
 sg13g2_a221oi_1 _5432_ (.B2(_1456_),
    .C1(_1581_),
    .B1(net857),
    .A1(net859),
    .Y(_1582_),
    .A2(_1438_));
 sg13g2_a21o_1 _5433_ (.A2(net852),
    .A1(net853),
    .B1(_1582_),
    .X(_1583_));
 sg13g2_nand3_1 _5434_ (.B(_1580_),
    .C(_1583_),
    .A(net865),
    .Y(_1584_));
 sg13g2_nor2b_1 _5435_ (.A(_1579_),
    .B_N(_1584_),
    .Y(_1585_));
 sg13g2_o21ai_1 _5436_ (.B1(net855),
    .Y(_1586_),
    .A1(_1578_),
    .A2(_1585_));
 sg13g2_nand3_1 _5437_ (.B(net862),
    .C(_1447_),
    .A(_1404_),
    .Y(_1587_));
 sg13g2_nand4_1 _5438_ (.B(_1438_),
    .C(net862),
    .A(net859),
    .Y(_1588_),
    .D(net857));
 sg13g2_nand4_1 _5439_ (.B(net852),
    .C(_1493_),
    .A(net853),
    .Y(_1589_),
    .D(_1588_));
 sg13g2_a22oi_1 _5440_ (.Y(_1590_),
    .B1(_1583_),
    .B2(_1589_),
    .A2(net843),
    .A1(net846));
 sg13g2_or3_1 _5441_ (.A(net865),
    .B(_1578_),
    .C(_1590_),
    .X(_1591_));
 sg13g2_o21ai_1 _5442_ (.B1(_1469_),
    .Y(_1592_),
    .A1(_1403_),
    .A2(_1446_));
 sg13g2_nand4_1 _5443_ (.B(_1438_),
    .C(_1587_),
    .A(net859),
    .Y(_1593_),
    .D(_1592_));
 sg13g2_o21ai_1 _5444_ (.B1(net857),
    .Y(_1594_),
    .A1(net860),
    .A2(net858));
 sg13g2_a22oi_1 _5445_ (.Y(_1595_),
    .B1(_1593_),
    .B2(_1594_),
    .A2(_1463_),
    .A1(_1462_));
 sg13g2_nor4_1 _5446_ (.A(_1429_),
    .B(_1430_),
    .C(net863),
    .D(_1595_),
    .Y(_1596_));
 sg13g2_nand4_1 _5447_ (.B(net852),
    .C(_1569_),
    .A(net853),
    .Y(_1597_),
    .D(_1593_));
 sg13g2_nand2b_1 _5448_ (.Y(_1598_),
    .B(_1597_),
    .A_N(_1577_));
 sg13g2_a221oi_1 _5449_ (.B2(_1579_),
    .C1(net855),
    .B1(_1598_),
    .A1(_1583_),
    .Y(_1599_),
    .A2(_1596_));
 sg13g2_a21oi_1 _5450_ (.A1(_1591_),
    .A2(_1599_),
    .Y(_1600_),
    .B1(_1523_));
 sg13g2_o21ai_1 _5451_ (.B1(_1600_),
    .Y(_1601_),
    .A1(_1574_),
    .A2(_1586_));
 sg13g2_nor2_1 _5452_ (.A(net841),
    .B(_1552_),
    .Y(_1602_));
 sg13g2_a22oi_1 _5453_ (.Y(_1603_),
    .B1(_1480_),
    .B2(_1471_),
    .A2(_1474_),
    .A1(_1441_));
 sg13g2_nand3b_1 _5454_ (.B(_1603_),
    .C(_1545_),
    .Y(_1604_),
    .A_N(_1582_));
 sg13g2_nand3_1 _5455_ (.B(_1525_),
    .C(_1602_),
    .A(_1431_),
    .Y(_1605_));
 sg13g2_and2_1 _5456_ (.A(_1604_),
    .B(_1605_),
    .X(_1606_));
 sg13g2_a221oi_1 _5457_ (.B2(_1432_),
    .C1(_1522_),
    .B1(_1555_),
    .A1(_1524_),
    .Y(_1607_),
    .A2(_1544_));
 sg13g2_a21oi_1 _5458_ (.A1(_1606_),
    .A2(_1607_),
    .Y(_1608_),
    .B1(_1543_));
 sg13g2_a21o_1 _5459_ (.A2(_1608_),
    .A1(_1601_),
    .B1(_1565_),
    .X(_1609_));
 sg13g2_o21ai_1 _5460_ (.B1(_1564_),
    .Y(_1610_),
    .A1(_3159_),
    .A2(_1561_));
 sg13g2_nand2_2 _5461_ (.Y(_1611_),
    .A(net970),
    .B(_3160_));
 sg13g2_xor2_1 _5462_ (.B(\vgademo.b_cos[11] ),
    .A(\vgademo.b_cos[10] ),
    .X(_1612_));
 sg13g2_mux2_1 _5463_ (.A0(net975),
    .A1(net963),
    .S(net875),
    .X(_1613_));
 sg13g2_xnor2_1 _5464_ (.Y(_1614_),
    .A(_1612_),
    .B(_1613_));
 sg13g2_xor2_1 _5465_ (.B(_1614_),
    .A(_1610_),
    .X(_1615_));
 sg13g2_a221oi_1 _5466_ (.B2(net863),
    .C1(net856),
    .B1(_1455_),
    .A1(_1439_),
    .Y(_1616_),
    .A2(_1440_));
 sg13g2_nor4_2 _5467_ (.A(_1429_),
    .B(_1430_),
    .C(net863),
    .Y(_1617_),
    .D(_1493_));
 sg13g2_o21ai_1 _5468_ (.B1(net861),
    .Y(_1618_),
    .A1(_1616_),
    .A2(_1617_));
 sg13g2_nand2_2 _5469_ (.Y(_1619_),
    .A(net861),
    .B(_1433_));
 sg13g2_and3_1 _5470_ (.X(_1620_),
    .A(_1455_),
    .B(_1530_),
    .C(_1619_));
 sg13g2_a22oi_1 _5471_ (.Y(_1621_),
    .B1(_1620_),
    .B2(_1432_),
    .A2(_1480_),
    .A1(_1444_));
 sg13g2_a21oi_1 _5472_ (.A1(_1618_),
    .A2(_1621_),
    .Y(_1622_),
    .B1(net839));
 sg13g2_a21o_1 _5473_ (.A2(_1479_),
    .A1(_1458_),
    .B1(_1467_),
    .X(_1623_));
 sg13g2_o21ai_1 _5474_ (.B1(_1522_),
    .Y(_1624_),
    .A1(_1622_),
    .A2(_1623_));
 sg13g2_nand2_1 _5475_ (.Y(_1625_),
    .A(_1466_),
    .B(_1482_));
 sg13g2_a21oi_1 _5476_ (.A1(net845),
    .A2(net842),
    .Y(_1626_),
    .B1(_1459_));
 sg13g2_nor2b_1 _5477_ (.A(_1457_),
    .B_N(_1532_),
    .Y(_1627_));
 sg13g2_and2_1 _5478_ (.A(_1475_),
    .B(_1627_),
    .X(_1628_));
 sg13g2_nand2_1 _5479_ (.Y(_1629_),
    .A(_1545_),
    .B(_1628_));
 sg13g2_a21oi_1 _5480_ (.A1(_1545_),
    .A2(_1628_),
    .Y(_1630_),
    .B1(_1626_));
 sg13g2_a21oi_1 _5481_ (.A1(_1625_),
    .A2(_1630_),
    .Y(_1631_),
    .B1(_1522_));
 sg13g2_nor2b_1 _5482_ (.A(_1631_),
    .B_N(_1565_),
    .Y(_1632_));
 sg13g2_a21oi_1 _5483_ (.A1(_1624_),
    .A2(_1632_),
    .Y(_1633_),
    .B1(_1615_));
 sg13g2_o21ai_1 _5484_ (.B1(_1633_),
    .Y(_1634_),
    .A1(_1560_),
    .A2(_1609_));
 sg13g2_nor4_1 _5485_ (.A(_1433_),
    .B(_1467_),
    .C(_1553_),
    .D(_1626_),
    .Y(_1635_));
 sg13g2_nor4_1 _5486_ (.A(net863),
    .B(_1553_),
    .C(_1556_),
    .D(_1558_),
    .Y(_1636_));
 sg13g2_o21ai_1 _5487_ (.B1(_1341_),
    .Y(_1637_),
    .A1(_1635_),
    .A2(_1636_));
 sg13g2_mux2_1 _5488_ (.A0(_1459_),
    .A1(_1547_),
    .S(_1545_),
    .X(_1638_));
 sg13g2_a21oi_1 _5489_ (.A1(net855),
    .A2(_1638_),
    .Y(_1639_),
    .B1(_1522_));
 sg13g2_nor4_2 _5490_ (.A(_1429_),
    .B(_1430_),
    .C(net841),
    .Y(_1640_),
    .D(_1473_));
 sg13g2_o21ai_1 _5491_ (.B1(net863),
    .Y(_1641_),
    .A1(_1529_),
    .A2(_1640_));
 sg13g2_a21o_1 _5492_ (.A2(_1588_),
    .A1(_1458_),
    .B1(_1494_),
    .X(_1642_));
 sg13g2_a21oi_1 _5493_ (.A1(_1579_),
    .A2(_1642_),
    .Y(_1643_),
    .B1(net861));
 sg13g2_nand2_1 _5494_ (.Y(_1644_),
    .A(net839),
    .B(_1566_));
 sg13g2_a21o_1 _5495_ (.A2(_1644_),
    .A1(_1528_),
    .B1(_1436_),
    .X(_1645_));
 sg13g2_nor3_1 _5496_ (.A(net848),
    .B(net844),
    .C(net865),
    .Y(_1646_));
 sg13g2_nand3_1 _5497_ (.B(net843),
    .C(net863),
    .A(net846),
    .Y(_1647_));
 sg13g2_a21oi_1 _5498_ (.A1(_1470_),
    .A2(_1475_),
    .Y(_1648_),
    .B1(_1442_));
 sg13g2_o21ai_1 _5499_ (.B1(_1646_),
    .Y(_1649_),
    .A1(_1494_),
    .A2(_1648_));
 sg13g2_nand4_1 _5500_ (.B(_1643_),
    .C(_1645_),
    .A(_1641_),
    .Y(_1650_),
    .D(_1649_));
 sg13g2_nor2_1 _5501_ (.A(net839),
    .B(_1566_),
    .Y(_1651_));
 sg13g2_nand3b_1 _5502_ (.B(net841),
    .C(_1493_),
    .Y(_1652_),
    .A_N(_1566_));
 sg13g2_nor4_1 _5503_ (.A(_1429_),
    .B(_1430_),
    .C(net841),
    .D(_1552_),
    .Y(_1653_));
 sg13g2_a221oi_1 _5504_ (.B2(_1579_),
    .C1(net855),
    .B1(_1652_),
    .A1(_1432_),
    .Y(_1654_),
    .A2(_1602_));
 sg13g2_or2_1 _5505_ (.X(_1655_),
    .B(_1627_),
    .A(_1494_));
 sg13g2_a21oi_1 _5506_ (.A1(_1646_),
    .A2(_1655_),
    .Y(_1656_),
    .B1(_1529_));
 sg13g2_a21oi_1 _5507_ (.A1(_1654_),
    .A2(_1656_),
    .Y(_1657_),
    .B1(_1523_));
 sg13g2_a221oi_1 _5508_ (.B2(_1657_),
    .C1(_1543_),
    .B1(_1650_),
    .A1(_1637_),
    .Y(_1658_),
    .A2(_1639_));
 sg13g2_o21ai_1 _5509_ (.B1(net864),
    .Y(_1659_),
    .A1(_1546_),
    .A2(_1603_));
 sg13g2_a21oi_1 _5510_ (.A1(_1523_),
    .A2(_1659_),
    .Y(_1660_),
    .B1(_1342_));
 sg13g2_nor2_1 _5511_ (.A(_1619_),
    .B(_1638_),
    .Y(_1661_));
 sg13g2_o21ai_1 _5512_ (.B1(net865),
    .Y(_1662_),
    .A1(_1529_),
    .A2(_1640_));
 sg13g2_a221oi_1 _5513_ (.B2(_1471_),
    .C1(net840),
    .B1(_1441_),
    .A1(net845),
    .Y(_1663_),
    .A2(net842));
 sg13g2_o21ai_1 _5514_ (.B1(net864),
    .Y(_1664_),
    .A1(_1478_),
    .A2(_1663_));
 sg13g2_nor3_1 _5515_ (.A(_1496_),
    .B(_1518_),
    .C(_1520_),
    .Y(_1665_));
 sg13g2_nand3_1 _5516_ (.B(_1664_),
    .C(_1665_),
    .A(_1662_),
    .Y(_1666_));
 sg13g2_o21ai_1 _5517_ (.B1(_1666_),
    .Y(_1667_),
    .A1(_1660_),
    .A2(_1661_));
 sg13g2_nor3_2 _5518_ (.A(_1466_),
    .B(_1518_),
    .C(_1520_),
    .Y(_1668_));
 sg13g2_nor2_1 _5519_ (.A(_1472_),
    .B(_1478_),
    .Y(_1669_));
 sg13g2_nand3_1 _5520_ (.B(_1545_),
    .C(_1603_),
    .A(_1458_),
    .Y(_1670_));
 sg13g2_a22oi_1 _5521_ (.Y(_1671_),
    .B1(_1546_),
    .B2(_1482_),
    .A2(_1521_),
    .A1(_1519_));
 sg13g2_a22oi_1 _5522_ (.Y(_1672_),
    .B1(_1670_),
    .B2(_1671_),
    .A2(_1669_),
    .A1(_1668_));
 sg13g2_a21oi_1 _5523_ (.A1(_1342_),
    .A2(_1672_),
    .Y(_1673_),
    .B1(_1542_));
 sg13g2_a21o_1 _5524_ (.A2(_1673_),
    .A1(_1667_),
    .B1(_1658_),
    .X(_1674_));
 sg13g2_nand4_1 _5525_ (.B(net841),
    .C(_1469_),
    .A(net856),
    .Y(_1675_),
    .D(_1569_));
 sg13g2_or3_1 _5526_ (.A(net865),
    .B(_1534_),
    .C(_1595_),
    .X(_1676_));
 sg13g2_a22oi_1 _5527_ (.Y(_1677_),
    .B1(_1676_),
    .B2(_1647_),
    .A2(_1675_),
    .A1(_1576_));
 sg13g2_a21oi_1 _5528_ (.A1(net846),
    .A2(net843),
    .Y(_1678_),
    .B1(_1589_));
 sg13g2_nor4_1 _5529_ (.A(net863),
    .B(_1576_),
    .C(_1653_),
    .D(_1678_),
    .Y(_1679_));
 sg13g2_or3_1 _5530_ (.A(net861),
    .B(_1677_),
    .C(_1679_),
    .X(_1680_));
 sg13g2_a21oi_1 _5531_ (.A1(net846),
    .A2(net843),
    .Y(_1681_),
    .B1(_1580_));
 sg13g2_or4_1 _5532_ (.A(net865),
    .B(_1576_),
    .C(_1653_),
    .D(_1681_),
    .X(_1682_));
 sg13g2_a21oi_1 _5533_ (.A1(_1568_),
    .A2(_1570_),
    .Y(_1683_),
    .B1(_1566_));
 sg13g2_a221oi_1 _5534_ (.B2(_1435_),
    .C1(net855),
    .B1(_1683_),
    .A1(_1579_),
    .Y(_1684_),
    .A2(_1651_));
 sg13g2_a21oi_1 _5535_ (.A1(_1682_),
    .A2(_1684_),
    .Y(_1685_),
    .B1(_1523_));
 sg13g2_mux2_1 _5536_ (.A0(_1604_),
    .A1(_1670_),
    .S(_1341_),
    .X(_1686_));
 sg13g2_nor3_1 _5537_ (.A(_1483_),
    .B(_1545_),
    .C(_1619_),
    .Y(_1687_));
 sg13g2_nor2_1 _5538_ (.A(_1545_),
    .B(_1552_),
    .Y(_1688_));
 sg13g2_a221oi_1 _5539_ (.B2(_1688_),
    .C1(_1687_),
    .B1(_1619_),
    .A1(_1519_),
    .Y(_1689_),
    .A2(_1521_));
 sg13g2_a221oi_1 _5540_ (.B2(_1689_),
    .C1(_1543_),
    .B1(_1686_),
    .A1(_1680_),
    .Y(_1690_),
    .A2(_1685_));
 sg13g2_a21oi_1 _5541_ (.A1(net853),
    .A2(net852),
    .Y(_1691_),
    .B1(net855));
 sg13g2_nand4_1 _5542_ (.B(_1462_),
    .C(_1463_),
    .A(net861),
    .Y(_1692_),
    .D(_1482_));
 sg13g2_o21ai_1 _5543_ (.B1(_1530_),
    .Y(_1693_),
    .A1(_1455_),
    .A2(_1524_));
 sg13g2_o21ai_1 _5544_ (.B1(_1692_),
    .Y(_1694_),
    .A1(net839),
    .A2(_1693_));
 sg13g2_nor3_1 _5545_ (.A(_1481_),
    .B(_1524_),
    .C(_1691_),
    .Y(_1695_));
 sg13g2_a221oi_1 _5546_ (.B2(_1432_),
    .C1(_1695_),
    .B1(_1694_),
    .A1(_1524_),
    .Y(_1696_),
    .A2(_1550_));
 sg13g2_a221oi_1 _5547_ (.B2(_1668_),
    .C1(_1542_),
    .B1(_1696_),
    .A1(_1629_),
    .Y(_1697_),
    .A2(_1671_));
 sg13g2_or2_1 _5548_ (.X(_1698_),
    .B(_1697_),
    .A(_1565_));
 sg13g2_o21ai_1 _5549_ (.B1(_1615_),
    .Y(_1699_),
    .A1(_1690_),
    .A2(_1698_));
 sg13g2_a21o_1 _5550_ (.A2(_1674_),
    .A1(_1565_),
    .B1(_1699_),
    .X(_1700_));
 sg13g2_nand2_1 _5551_ (.Y(_1701_),
    .A(_1505_),
    .B(_1506_));
 sg13g2_xnor2_1 _5552_ (.Y(_1702_),
    .A(net989),
    .B(_1701_));
 sg13g2_xnor2_1 _5553_ (.Y(_1703_),
    .A(net988),
    .B(_1022_));
 sg13g2_nand2_1 _5554_ (.Y(_1704_),
    .A(_1501_),
    .B(_1703_));
 sg13g2_xor2_1 _5555_ (.B(_1703_),
    .A(_1501_),
    .X(_1705_));
 sg13g2_a221oi_1 _5556_ (.B2(_1352_),
    .C1(_1353_),
    .B1(_1705_),
    .A1(_1359_),
    .Y(_1706_),
    .A2(_1702_));
 sg13g2_xnor2_1 _5557_ (.Y(_1707_),
    .A(\vgademo.h_count[10] ),
    .B(_1510_));
 sg13g2_nor2_1 _5558_ (.A(net874),
    .B(_1707_),
    .Y(_1708_));
 sg13g2_a21oi_2 _5559_ (.B1(_1708_),
    .Y(_1709_),
    .A2(net874),
    .A1(_0032_));
 sg13g2_nand2_1 _5560_ (.Y(_1710_),
    .A(_1706_),
    .B(_1709_));
 sg13g2_nor2_1 _5561_ (.A(_1515_),
    .B(_1518_),
    .Y(_1711_));
 sg13g2_a21oi_1 _5562_ (.A1(_1022_),
    .A2(_1023_),
    .Y(_1712_),
    .B1(_1350_));
 sg13g2_xnor2_1 _5563_ (.Y(_1713_),
    .A(_1704_),
    .B(_1712_));
 sg13g2_a21oi_1 _5564_ (.A1(_1379_),
    .A2(_1713_),
    .Y(_1714_),
    .B1(_1359_));
 sg13g2_a21oi_1 _5565_ (.A1(net988),
    .A2(_1701_),
    .Y(_1715_),
    .B1(net984));
 sg13g2_nor3_1 _5566_ (.A(_1357_),
    .B(_1358_),
    .C(_1715_),
    .Y(_1716_));
 sg13g2_nor3_2 _5567_ (.A(_1349_),
    .B(_1714_),
    .C(_1716_),
    .Y(_1717_));
 sg13g2_o21ai_1 _5568_ (.B1(net1006),
    .Y(_1718_),
    .A1(\vgademo.h_count[10] ),
    .A2(_1511_));
 sg13g2_nor2_1 _5569_ (.A(net874),
    .B(_1718_),
    .Y(_1719_));
 sg13g2_a21oi_1 _5570_ (.A1(\vgademo.plane_u[21] ),
    .A2(net874),
    .Y(_1720_),
    .B1(_1719_));
 sg13g2_xnor2_1 _5571_ (.Y(_1721_),
    .A(_1717_),
    .B(_1720_));
 sg13g2_o21ai_1 _5572_ (.B1(_1710_),
    .Y(_1722_),
    .A1(_1711_),
    .A2(_1721_));
 sg13g2_nor2_1 _5573_ (.A(_1706_),
    .B(_1709_),
    .Y(_1723_));
 sg13g2_nor2_1 _5574_ (.A(_1721_),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_nor2_1 _5575_ (.A(_1711_),
    .B(_1724_),
    .Y(_1725_));
 sg13g2_mux2_1 _5576_ (.A0(_1724_),
    .A1(_1725_),
    .S(_1722_),
    .X(_1726_));
 sg13g2_nor2_1 _5577_ (.A(_3158_),
    .B(_1611_),
    .Y(_1727_));
 sg13g2_or2_1 _5578_ (.X(_1728_),
    .B(_1611_),
    .A(_3158_));
 sg13g2_a22oi_1 _5579_ (.Y(_1729_),
    .B1(_1326_),
    .B2(net971),
    .A2(\vgademo.b_cos[7] ),
    .A1(_3111_));
 sg13g2_o21ai_1 _5580_ (.B1(_1729_),
    .Y(_1730_),
    .A1(\vgademo.bayer_j[1] ),
    .A2(_1327_));
 sg13g2_a22oi_1 _5581_ (.Y(_1731_),
    .B1(_3157_),
    .B2(\vgademo.v_count[3] ),
    .A2(_3156_),
    .A1(\vgademo.v_count[2] ));
 sg13g2_a22oi_1 _5582_ (.Y(_1732_),
    .B1(_1730_),
    .B2(_1731_),
    .A2(\vgademo.b_cos[8] ),
    .A1(_3110_));
 sg13g2_o21ai_1 _5583_ (.B1(_1732_),
    .Y(_1733_),
    .A1(net978),
    .A2(_3158_));
 sg13g2_a22oi_1 _5584_ (.Y(_1734_),
    .B1(\vgademo.b_cos[10] ),
    .B2(net976),
    .A2(_3158_),
    .A1(net978));
 sg13g2_xnor2_1 _5585_ (.Y(_1735_),
    .A(_0016_),
    .B(_1612_));
 sg13g2_o21ai_1 _5586_ (.B1(_1735_),
    .Y(_1736_),
    .A1(net976),
    .A2(net970));
 sg13g2_a21oi_1 _5587_ (.A1(_1733_),
    .A2(_1734_),
    .Y(_1737_),
    .B1(_1736_));
 sg13g2_a221oi_1 _5588_ (.B2(net975),
    .C1(_1737_),
    .B1(_1612_),
    .A1(net974),
    .Y(_1738_),
    .A2(_1611_));
 sg13g2_nor2_1 _5589_ (.A(net973),
    .B(_3135_),
    .Y(_1739_));
 sg13g2_o21ai_1 _5590_ (.B1(_1739_),
    .Y(_1740_),
    .A1(net974),
    .A2(_1611_));
 sg13g2_o21ai_1 _5591_ (.B1(_0021_),
    .Y(_1741_),
    .A1(_1738_),
    .A2(_1740_));
 sg13g2_a22oi_1 _5592_ (.Y(_1742_),
    .B1(_1741_),
    .B2(_1299_),
    .A2(_1727_),
    .A1(_3241_));
 sg13g2_xnor2_1 _5593_ (.Y(_1743_),
    .A(\vgademo.b_cos[9] ),
    .B(net970));
 sg13g2_xnor2_1 _5594_ (.Y(_1744_),
    .A(_0063_),
    .B(_1743_));
 sg13g2_o21ai_1 _5595_ (.B1(_1732_),
    .Y(_1745_),
    .A1(net978),
    .A2(\vgademo.b_cos[9] ));
 sg13g2_o21ai_1 _5596_ (.B1(_1745_),
    .Y(_1746_),
    .A1(_3112_),
    .A2(_3158_));
 sg13g2_a22oi_1 _5597_ (.Y(_1747_),
    .B1(_1744_),
    .B2(_1746_),
    .A2(_1743_),
    .A1(net976));
 sg13g2_mux2_2 _5598_ (.A0(\vgademo.b_cos[11] ),
    .A1(_1612_),
    .S(\vgademo.b_cos[9] ),
    .X(_1748_));
 sg13g2_xor2_1 _5599_ (.B(_1748_),
    .A(_0016_),
    .X(_1749_));
 sg13g2_a22oi_1 _5600_ (.Y(_1750_),
    .B1(_1748_),
    .B2(net975),
    .A2(_3135_),
    .A1(net974));
 sg13g2_o21ai_1 _5601_ (.B1(_1750_),
    .Y(_1751_),
    .A1(_1747_),
    .A2(_1749_));
 sg13g2_nand3_1 _5602_ (.B(_0018_),
    .C(_1728_),
    .A(net974),
    .Y(_1752_));
 sg13g2_o21ai_1 _5603_ (.B1(_1752_),
    .Y(_1753_),
    .A1(_0018_),
    .A2(_1728_));
 sg13g2_a21o_1 _5604_ (.A2(_1753_),
    .A1(_1751_),
    .B1(_1742_),
    .X(_1754_));
 sg13g2_inv_1 _5605_ (.Y(_1755_),
    .A(_1754_));
 sg13g2_and4_2 _5606_ (.A(_1634_),
    .B(_1700_),
    .C(_1726_),
    .D(_1755_),
    .X(_1756_));
 sg13g2_nand4_1 _5607_ (.B(_1700_),
    .C(_1726_),
    .A(_1634_),
    .Y(_1757_),
    .D(_1755_));
 sg13g2_nand2_1 _5608_ (.Y(_1758_),
    .A(\vgademo.plane_du[7] ),
    .B(_1743_));
 sg13g2_xor2_1 _5609_ (.B(_1743_),
    .A(_0053_),
    .X(_1759_));
 sg13g2_a22oi_1 _5610_ (.Y(_1760_),
    .B1(_1330_),
    .B2(net971),
    .A2(_3171_),
    .A1(\vgademo.b_cos[7] ));
 sg13g2_o21ai_1 _5611_ (.B1(_1760_),
    .Y(_1761_),
    .A1(\vgademo.plane_du[3] ),
    .A2(_1332_));
 sg13g2_a22oi_1 _5612_ (.Y(_1762_),
    .B1(\vgademo.plane_du[5] ),
    .B2(_3157_),
    .A2(\vgademo.plane_du[4] ),
    .A1(_3156_));
 sg13g2_a22oi_1 _5613_ (.Y(_1763_),
    .B1(_1761_),
    .B2(_1762_),
    .A2(_3173_),
    .A1(\vgademo.b_cos[8] ));
 sg13g2_and2_1 _5614_ (.A(\vgademo.plane_du[6] ),
    .B(_1763_),
    .X(_1764_));
 sg13g2_or2_1 _5615_ (.X(_1765_),
    .B(_1763_),
    .A(\vgademo.plane_du[6] ));
 sg13g2_o21ai_1 _5616_ (.B1(_1765_),
    .Y(_1766_),
    .A1(\vgademo.b_cos[9] ),
    .A2(_1764_));
 sg13g2_o21ai_1 _5617_ (.B1(_1758_),
    .Y(_1767_),
    .A1(_1759_),
    .A2(_1766_));
 sg13g2_xnor2_1 _5618_ (.Y(_1768_),
    .A(_0054_),
    .B(_1748_));
 sg13g2_a22oi_1 _5619_ (.Y(_1769_),
    .B1(_1767_),
    .B2(_1768_),
    .A2(_1748_),
    .A1(net963));
 sg13g2_nand2_1 _5620_ (.Y(_1770_),
    .A(net962),
    .B(_1728_));
 sg13g2_a221oi_1 _5621_ (.B2(_3158_),
    .C1(_1764_),
    .B1(_1765_),
    .A1(net970),
    .Y(_1771_),
    .A2(\vgademo.plane_du[7] ));
 sg13g2_xnor2_1 _5622_ (.Y(_1772_),
    .A(_0054_),
    .B(_1612_));
 sg13g2_o21ai_1 _5623_ (.B1(_1772_),
    .Y(_1773_),
    .A1(net970),
    .A2(\vgademo.plane_du[7] ));
 sg13g2_a22oi_1 _5624_ (.Y(_1774_),
    .B1(_1612_),
    .B2(net963),
    .A2(_1611_),
    .A1(net962));
 sg13g2_o21ai_1 _5625_ (.B1(_1774_),
    .Y(_1775_),
    .A1(_1771_),
    .A2(_1773_));
 sg13g2_nor2_1 _5626_ (.A(net962),
    .B(_1611_),
    .Y(_1776_));
 sg13g2_o21ai_1 _5627_ (.B1(_1775_),
    .Y(_1777_),
    .A1(_1769_),
    .A2(_1770_));
 sg13g2_nor2_2 _5628_ (.A(_1776_),
    .B(_1777_),
    .Y(_1778_));
 sg13g2_nand4_1 _5629_ (.B(_1700_),
    .C(_1726_),
    .A(_1634_),
    .Y(_1779_),
    .D(_1778_));
 sg13g2_xor2_1 _5630_ (.B(\vgademo.plane_du[7] ),
    .A(net996),
    .X(_1780_));
 sg13g2_xnor2_1 _5631_ (.Y(_1781_),
    .A(net999),
    .B(\vgademo.plane_du[6] ));
 sg13g2_nand2_1 _5632_ (.Y(_1782_),
    .A(net1002),
    .B(\vgademo.plane_du[5] ));
 sg13g2_nand2_1 _5633_ (.Y(_1783_),
    .A(_3130_),
    .B(_3173_));
 sg13g2_nor2_1 _5634_ (.A(_3123_),
    .B(_3171_),
    .Y(_1784_));
 sg13g2_nand3_1 _5635_ (.B(_1783_),
    .C(_1784_),
    .A(_1782_),
    .Y(_1785_));
 sg13g2_a21oi_1 _5636_ (.A1(_1782_),
    .A2(_1785_),
    .Y(_1786_),
    .B1(_1781_));
 sg13g2_a21oi_1 _5637_ (.A1(net1000),
    .A2(\vgademo.plane_du[6] ),
    .Y(_1787_),
    .B1(_1786_));
 sg13g2_nand2b_1 _5638_ (.Y(_1788_),
    .B(_1780_),
    .A_N(_1787_));
 sg13g2_xnor2_1 _5639_ (.Y(_1789_),
    .A(_1780_),
    .B(_1787_));
 sg13g2_nand2_1 _5640_ (.Y(_1790_),
    .A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ));
 sg13g2_xnor2_1 _5641_ (.Y(_1791_),
    .A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ));
 sg13g2_xnor2_1 _5642_ (.Y(_1792_),
    .A(\vgademo.a_cos[9] ),
    .B(\vgademo.plane_u[14] ));
 sg13g2_nand2_1 _5643_ (.Y(_1793_),
    .A(\vgademo.a_cos[8] ),
    .B(\vgademo.plane_u[13] ));
 sg13g2_xnor2_1 _5644_ (.Y(_1794_),
    .A(\vgademo.a_cos[8] ),
    .B(\vgademo.plane_u[13] ));
 sg13g2_nand2_1 _5645_ (.Y(_1795_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.plane_u[12] ));
 sg13g2_xnor2_1 _5646_ (.Y(_1796_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.plane_u[12] ));
 sg13g2_or2_1 _5647_ (.X(_1797_),
    .B(\vgademo.plane_u[10] ),
    .A(\vgademo.a_cos[5] ));
 sg13g2_nand3_1 _5648_ (.B(\vgademo.plane_u[9] ),
    .C(_1797_),
    .A(\vgademo.a_cos[4] ),
    .Y(_1798_));
 sg13g2_a22oi_1 _5649_ (.Y(_1799_),
    .B1(\vgademo.plane_u[11] ),
    .B2(\vgademo.a_cos[6] ),
    .A2(\vgademo.plane_u[10] ),
    .A1(\vgademo.a_cos[5] ));
 sg13g2_a22oi_1 _5650_ (.Y(_1800_),
    .B1(_1798_),
    .B2(_1799_),
    .A2(_3181_),
    .A1(_3153_));
 sg13g2_nand2b_1 _5651_ (.Y(_1801_),
    .B(_1800_),
    .A_N(_1796_));
 sg13g2_a21o_1 _5652_ (.A2(_1801_),
    .A1(_1795_),
    .B1(_1794_),
    .X(_1802_));
 sg13g2_a21oi_1 _5653_ (.A1(_1793_),
    .A2(_1802_),
    .Y(_1803_),
    .B1(_1792_));
 sg13g2_a21oi_2 _5654_ (.B1(_1803_),
    .Y(_1804_),
    .A2(\vgademo.plane_u[14] ),
    .A1(\vgademo.a_cos[9] ));
 sg13g2_o21ai_1 _5655_ (.B1(_1790_),
    .Y(_1805_),
    .A1(_1791_),
    .A2(_1804_));
 sg13g2_and2_1 _5656_ (.A(\vgademo.a_cos[11] ),
    .B(\vgademo.plane_u[16] ),
    .X(_1806_));
 sg13g2_xor2_1 _5657_ (.B(\vgademo.plane_u[16] ),
    .A(\vgademo.a_cos[11] ),
    .X(_1807_));
 sg13g2_xnor2_1 _5658_ (.Y(_1808_),
    .A(_1805_),
    .B(_1807_));
 sg13g2_inv_1 _5659_ (.Y(_1809_),
    .A(_1808_));
 sg13g2_xor2_1 _5660_ (.B(_1808_),
    .A(_1789_),
    .X(_1810_));
 sg13g2_o21ai_1 _5661_ (.B1(_1788_),
    .Y(_1811_),
    .A1(_3129_),
    .A2(_3176_));
 sg13g2_and2_1 _5662_ (.A(net994),
    .B(net963),
    .X(_1812_));
 sg13g2_xor2_1 _5663_ (.B(net963),
    .A(net993),
    .X(_1813_));
 sg13g2_xnor2_1 _5664_ (.Y(_1814_),
    .A(_1811_),
    .B(_1813_));
 sg13g2_nor2_1 _5665_ (.A(_1810_),
    .B(_1814_),
    .Y(_1815_));
 sg13g2_and2_1 _5666_ (.A(net991),
    .B(net962),
    .X(_1816_));
 sg13g2_xor2_1 _5667_ (.B(net962),
    .A(net991),
    .X(_1817_));
 sg13g2_a21o_1 _5668_ (.A2(_1813_),
    .A1(_1811_),
    .B1(_1812_),
    .X(_1818_));
 sg13g2_xnor2_1 _5669_ (.Y(_1819_),
    .A(_1817_),
    .B(_1818_));
 sg13g2_and2_1 _5670_ (.A(\vgademo.a_cos[12] ),
    .B(\vgademo.plane_u[17] ),
    .X(_1820_));
 sg13g2_a21o_1 _5671_ (.A2(_1807_),
    .A1(_1805_),
    .B1(_1806_),
    .X(_1821_));
 sg13g2_xor2_1 _5672_ (.B(\vgademo.plane_u[17] ),
    .A(\vgademo.a_cos[12] ),
    .X(_1822_));
 sg13g2_a21o_1 _5673_ (.A2(_1822_),
    .A1(_1821_),
    .B1(_1820_),
    .X(_1823_));
 sg13g2_xor2_1 _5674_ (.B(\vgademo.plane_u[18] ),
    .A(\vgademo.a_cos[13] ),
    .X(_1824_));
 sg13g2_xnor2_1 _5675_ (.Y(_1825_),
    .A(_1823_),
    .B(_1824_));
 sg13g2_nor2_1 _5676_ (.A(_1819_),
    .B(_1825_),
    .Y(_1826_));
 sg13g2_xor2_1 _5677_ (.B(_1825_),
    .A(_1819_),
    .X(_1827_));
 sg13g2_xnor2_1 _5678_ (.Y(_1828_),
    .A(_1821_),
    .B(_1822_));
 sg13g2_xor2_1 _5679_ (.B(_1828_),
    .A(_1814_),
    .X(_1829_));
 sg13g2_nand3_1 _5680_ (.B(_1809_),
    .C(_1829_),
    .A(_1789_),
    .Y(_1830_));
 sg13g2_o21ai_1 _5681_ (.B1(_1830_),
    .Y(_1831_),
    .A1(_1814_),
    .A2(_1828_));
 sg13g2_a21oi_1 _5682_ (.A1(_1827_),
    .A2(_1831_),
    .Y(_1832_),
    .B1(_1826_));
 sg13g2_a21o_1 _5683_ (.A2(\vgademo.plane_u[18] ),
    .A1(\vgademo.a_cos[13] ),
    .B1(_1823_),
    .X(_1833_));
 sg13g2_o21ai_1 _5684_ (.B1(_1833_),
    .Y(_1834_),
    .A1(\vgademo.a_cos[13] ),
    .A2(\vgademo.plane_u[18] ));
 sg13g2_a21oi_1 _5685_ (.A1(_1817_),
    .A2(_1818_),
    .Y(_1835_),
    .B1(_1816_));
 sg13g2_xor2_1 _5686_ (.B(\vgademo.a_cos[14] ),
    .A(net989),
    .X(_1836_));
 sg13g2_xor2_1 _5687_ (.B(\vgademo.plane_u[19] ),
    .A(\vgademo.plane_du[10] ),
    .X(_1837_));
 sg13g2_xnor2_1 _5688_ (.Y(_1838_),
    .A(_1836_),
    .B(_1837_));
 sg13g2_xnor2_1 _5689_ (.Y(_1839_),
    .A(_1835_),
    .B(_1838_));
 sg13g2_xnor2_1 _5690_ (.Y(_1840_),
    .A(_1834_),
    .B(_1839_));
 sg13g2_xnor2_1 _5691_ (.Y(_1841_),
    .A(_1832_),
    .B(_1840_));
 sg13g2_xnor2_1 _5692_ (.Y(_1842_),
    .A(_1827_),
    .B(_1831_));
 sg13g2_or3_1 _5693_ (.A(net1054),
    .B(net1057),
    .C(_1810_),
    .X(_1843_));
 sg13g2_a21o_1 _5694_ (.A2(_1809_),
    .A1(_1789_),
    .B1(_1829_),
    .X(_1844_));
 sg13g2_o21ai_1 _5695_ (.B1(net1054),
    .Y(_1845_),
    .A1(net1057),
    .A2(_1810_));
 sg13g2_nand3_1 _5696_ (.B(_1844_),
    .C(_1845_),
    .A(_1830_),
    .Y(_1846_));
 sg13g2_nor2_1 _5697_ (.A(net1051),
    .B(_1842_),
    .Y(_1847_));
 sg13g2_a22oi_1 _5698_ (.Y(_1848_),
    .B1(_1843_),
    .B2(_1846_),
    .A2(_1842_),
    .A1(net1051));
 sg13g2_nor2_1 _5699_ (.A(_1847_),
    .B(_1848_),
    .Y(_1849_));
 sg13g2_a21oi_1 _5700_ (.A1(net1048),
    .A2(_1841_),
    .Y(_1850_),
    .B1(_1849_));
 sg13g2_nor2_1 _5701_ (.A(net1048),
    .B(_1841_),
    .Y(_1851_));
 sg13g2_nor4_2 _5702_ (.A(_3107_),
    .B(_3122_),
    .C(_1850_),
    .Y(_1852_),
    .D(_1851_));
 sg13g2_xnor2_1 _5703_ (.Y(_1853_),
    .A(net1057),
    .B(_1829_));
 sg13g2_xnor2_1 _5704_ (.Y(_1854_),
    .A(net1054),
    .B(_1789_));
 sg13g2_xor2_1 _5705_ (.B(_1808_),
    .A(net1060),
    .X(_1855_));
 sg13g2_nand4_1 _5706_ (.B(_1853_),
    .C(_1854_),
    .A(\vgademo.audio_songpos[7] ),
    .Y(_1856_),
    .D(_1855_));
 sg13g2_a21oi_1 _5707_ (.A1(_3098_),
    .A2(_1827_),
    .Y(_1857_),
    .B1(_1856_));
 sg13g2_o21ai_1 _5708_ (.B1(_1857_),
    .Y(_1858_),
    .A1(_3098_),
    .A2(_1827_));
 sg13g2_inv_2 _5709_ (.Y(_1859_),
    .A(_1858_));
 sg13g2_nand2b_1 _5710_ (.Y(_1860_),
    .B(_1858_),
    .A_N(_1852_));
 sg13g2_inv_1 _5711_ (.Y(_1861_),
    .A(_1860_));
 sg13g2_nor2_2 _5712_ (.A(_1815_),
    .B(_1860_),
    .Y(_1862_));
 sg13g2_nor2_1 _5713_ (.A(net866),
    .B(_1862_),
    .Y(_1863_));
 sg13g2_nand2_1 _5714_ (.Y(_1864_),
    .A(net1066),
    .B(net990));
 sg13g2_nand2_1 _5715_ (.Y(_1865_),
    .A(net992),
    .B(net1064));
 sg13g2_nand2_1 _5716_ (.Y(_1866_),
    .A(net990),
    .B(net1064));
 sg13g2_nand2_1 _5717_ (.Y(_1867_),
    .A(net1066),
    .B(net992));
 sg13g2_xor2_1 _5718_ (.B(_1867_),
    .A(_1866_),
    .X(_1868_));
 sg13g2_nand2_1 _5719_ (.Y(_1869_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1868_));
 sg13g2_o21ai_1 _5720_ (.B1(_1869_),
    .Y(_1870_),
    .A1(_1866_),
    .A2(_1867_));
 sg13g2_nand2_1 _5721_ (.Y(_1871_),
    .A(net987),
    .B(net1064));
 sg13g2_xor2_1 _5722_ (.B(_1871_),
    .A(_1864_),
    .X(_1872_));
 sg13g2_nand2_1 _5723_ (.Y(_1873_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1872_));
 sg13g2_xnor2_1 _5724_ (.Y(_1874_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1872_));
 sg13g2_nand2b_1 _5725_ (.Y(_1875_),
    .B(_1870_),
    .A_N(_1874_));
 sg13g2_xor2_1 _5726_ (.B(_1874_),
    .A(_1870_),
    .X(_1876_));
 sg13g2_o21ai_1 _5727_ (.B1(_1875_),
    .Y(_1877_),
    .A1(_3125_),
    .A2(_1876_));
 sg13g2_o21ai_1 _5728_ (.B1(_1873_),
    .Y(_1878_),
    .A1(_1864_),
    .A2(_1871_));
 sg13g2_nand2_1 _5729_ (.Y(_1879_),
    .A(net1066),
    .B(net986));
 sg13g2_nor2_1 _5730_ (.A(_1871_),
    .B(_1879_),
    .Y(_1880_));
 sg13g2_a22oi_1 _5731_ (.Y(_1881_),
    .B1(net1063),
    .B2(net986),
    .A2(net987),
    .A1(net1065));
 sg13g2_nor2_1 _5732_ (.A(_1880_),
    .B(_1881_),
    .Y(_1882_));
 sg13g2_xnor2_1 _5733_ (.Y(_1883_),
    .A(\vgademo.linelfsr[11] ),
    .B(_1882_));
 sg13g2_nand2b_1 _5734_ (.Y(_1884_),
    .B(_1878_),
    .A_N(_1883_));
 sg13g2_xor2_1 _5735_ (.B(_1883_),
    .A(_1878_),
    .X(_1885_));
 sg13g2_xnor2_1 _5736_ (.Y(_1886_),
    .A(_3124_),
    .B(_1885_));
 sg13g2_nand2b_1 _5737_ (.Y(_1887_),
    .B(_1877_),
    .A_N(_1886_));
 sg13g2_nand2_1 _5738_ (.Y(_1888_),
    .A(net995),
    .B(net1063));
 sg13g2_nand2_1 _5739_ (.Y(_1889_),
    .A(net1065),
    .B(net995));
 sg13g2_xor2_1 _5740_ (.B(_1889_),
    .A(_1865_),
    .X(_1890_));
 sg13g2_nand2_1 _5741_ (.Y(_1891_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1890_));
 sg13g2_o21ai_1 _5742_ (.B1(_1891_),
    .Y(_1892_),
    .A1(_1865_),
    .A2(_1889_));
 sg13g2_xnor2_1 _5743_ (.Y(_1893_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1868_));
 sg13g2_nand2b_1 _5744_ (.Y(_1894_),
    .B(_1892_),
    .A_N(_1893_));
 sg13g2_xor2_1 _5745_ (.B(_1893_),
    .A(_1892_),
    .X(_1895_));
 sg13g2_o21ai_1 _5746_ (.B1(_1894_),
    .Y(_1896_),
    .A1(net956),
    .A2(_1895_));
 sg13g2_xnor2_1 _5747_ (.Y(_1897_),
    .A(_3125_),
    .B(_1876_));
 sg13g2_nor2b_1 _5748_ (.A(_1897_),
    .B_N(_1896_),
    .Y(_1898_));
 sg13g2_xor2_1 _5749_ (.B(_1897_),
    .A(_1896_),
    .X(_1899_));
 sg13g2_xnor2_1 _5750_ (.Y(_1900_),
    .A(net956),
    .B(_1895_));
 sg13g2_nand2_1 _5751_ (.Y(_1901_),
    .A(net997),
    .B(net1063));
 sg13g2_nand2_1 _5752_ (.Y(_1902_),
    .A(net1065),
    .B(net997));
 sg13g2_xor2_1 _5753_ (.B(_1902_),
    .A(_1888_),
    .X(_1903_));
 sg13g2_nand2_1 _5754_ (.Y(_1904_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1903_));
 sg13g2_o21ai_1 _5755_ (.B1(_1904_),
    .Y(_1905_),
    .A1(_1888_),
    .A2(_1902_));
 sg13g2_xnor2_1 _5756_ (.Y(_1906_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1890_));
 sg13g2_nand2b_1 _5757_ (.Y(_1907_),
    .B(_1905_),
    .A_N(_1906_));
 sg13g2_xor2_1 _5758_ (.B(_1906_),
    .A(_1905_),
    .X(_1908_));
 sg13g2_o21ai_1 _5759_ (.B1(_1907_),
    .Y(_1909_),
    .A1(_3127_),
    .A2(_1908_));
 sg13g2_nor2b_1 _5760_ (.A(_1909_),
    .B_N(_1900_),
    .Y(_1910_));
 sg13g2_nand2b_1 _5761_ (.Y(_1911_),
    .B(_1909_),
    .A_N(_1900_));
 sg13g2_nand2_1 _5762_ (.Y(_1912_),
    .A(net1065),
    .B(net1001));
 sg13g2_xor2_1 _5763_ (.B(_1912_),
    .A(_1901_),
    .X(_1913_));
 sg13g2_nand2_1 _5764_ (.Y(_1914_),
    .A(\vgademo.linelfsr[6] ),
    .B(_1913_));
 sg13g2_o21ai_1 _5765_ (.B1(_1914_),
    .Y(_1915_),
    .A1(_1901_),
    .A2(_1912_));
 sg13g2_xnor2_1 _5766_ (.Y(_1916_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1903_));
 sg13g2_nand2b_1 _5767_ (.Y(_1917_),
    .B(_1915_),
    .A_N(_1916_));
 sg13g2_xor2_1 _5768_ (.B(_1916_),
    .A(_1915_),
    .X(_1918_));
 sg13g2_o21ai_1 _5769_ (.B1(_1917_),
    .Y(_1919_),
    .A1(_3128_),
    .A2(_1918_));
 sg13g2_xnor2_1 _5770_ (.Y(_1920_),
    .A(_3127_),
    .B(_1908_));
 sg13g2_nor2b_1 _5771_ (.A(_1920_),
    .B_N(_1919_),
    .Y(_1921_));
 sg13g2_xnor2_1 _5772_ (.Y(_1922_),
    .A(_1919_),
    .B(_1920_));
 sg13g2_nor3_1 _5773_ (.A(_3123_),
    .B(_3190_),
    .C(_1912_),
    .Y(_1923_));
 sg13g2_a22oi_1 _5774_ (.Y(_1924_),
    .B1(net1001),
    .B2(net1063),
    .A2(net1003),
    .A1(net1065));
 sg13g2_nor3_1 _5775_ (.A(_3191_),
    .B(_1923_),
    .C(_1924_),
    .Y(_1925_));
 sg13g2_or2_1 _5776_ (.X(_1926_),
    .B(_1925_),
    .A(_1923_));
 sg13g2_xnor2_1 _5777_ (.Y(_1927_),
    .A(\vgademo.linelfsr[6] ),
    .B(_1913_));
 sg13g2_nand2b_1 _5778_ (.Y(_1928_),
    .B(_1926_),
    .A_N(_1927_));
 sg13g2_xor2_1 _5779_ (.B(_1927_),
    .A(_1926_),
    .X(_1929_));
 sg13g2_o21ai_1 _5780_ (.B1(_1928_),
    .Y(_1930_),
    .A1(_3129_),
    .A2(_1929_));
 sg13g2_xnor2_1 _5781_ (.Y(_1931_),
    .A(_3128_),
    .B(_1918_));
 sg13g2_nand2b_1 _5782_ (.Y(_1932_),
    .B(_1930_),
    .A_N(_1931_));
 sg13g2_nor2b_1 _5783_ (.A(_1930_),
    .B_N(_1931_),
    .Y(_1933_));
 sg13g2_nand3_1 _5784_ (.B(net1063),
    .C(\vgademo.linelfsr[4] ),
    .A(net1004),
    .Y(_1934_));
 sg13g2_a21o_1 _5785_ (.A2(net1063),
    .A1(net1004),
    .B1(\vgademo.linelfsr[4] ),
    .X(_1935_));
 sg13g2_nand2_1 _5786_ (.Y(_1936_),
    .A(_1934_),
    .B(_1935_));
 sg13g2_o21ai_1 _5787_ (.B1(_1934_),
    .Y(_1937_),
    .A1(_3130_),
    .A2(_1936_));
 sg13g2_o21ai_1 _5788_ (.B1(_3191_),
    .Y(_1938_),
    .A1(_1923_),
    .A2(_1924_));
 sg13g2_nand2b_1 _5789_ (.Y(_1939_),
    .B(_1938_),
    .A_N(_1925_));
 sg13g2_nor2b_1 _5790_ (.A(_1939_),
    .B_N(_1937_),
    .Y(_1940_));
 sg13g2_nand2b_1 _5791_ (.Y(_1941_),
    .B(_1939_),
    .A_N(_1937_));
 sg13g2_nand2b_1 _5792_ (.Y(_1942_),
    .B(_1941_),
    .A_N(_1940_));
 sg13g2_a21o_1 _5793_ (.A2(_1941_),
    .A1(net997),
    .B1(_1940_),
    .X(_1943_));
 sg13g2_xnor2_1 _5794_ (.Y(_1944_),
    .A(_3129_),
    .B(_1929_));
 sg13g2_nor2b_1 _5795_ (.A(_1944_),
    .B_N(_1943_),
    .Y(_1945_));
 sg13g2_xor2_1 _5796_ (.B(_1942_),
    .A(net997),
    .X(_1946_));
 sg13g2_xnor2_1 _5797_ (.Y(_1947_),
    .A(_3130_),
    .B(_1936_));
 sg13g2_nand2_1 _5798_ (.Y(_1948_),
    .A(\vgademo.linelfsr[3] ),
    .B(net1004));
 sg13g2_nor2_1 _5799_ (.A(_1947_),
    .B(_1948_),
    .Y(_1949_));
 sg13g2_nor2b_1 _5800_ (.A(_1946_),
    .B_N(_1949_),
    .Y(_1950_));
 sg13g2_xor2_1 _5801_ (.B(_1944_),
    .A(_1943_),
    .X(_1951_));
 sg13g2_inv_1 _5802_ (.Y(_1952_),
    .A(_1951_));
 sg13g2_a21oi_1 _5803_ (.A1(_1950_),
    .A2(_1952_),
    .Y(_1953_),
    .B1(_1945_));
 sg13g2_a21oi_1 _5804_ (.A1(_1932_),
    .A2(_1953_),
    .Y(_1954_),
    .B1(_1933_));
 sg13g2_a21oi_1 _5805_ (.A1(_1922_),
    .A2(_1954_),
    .Y(_1955_),
    .B1(_1921_));
 sg13g2_o21ai_1 _5806_ (.B1(_1911_),
    .Y(_1956_),
    .A1(_1910_),
    .A2(_1955_));
 sg13g2_nor2b_1 _5807_ (.A(_1899_),
    .B_N(_1956_),
    .Y(_1957_));
 sg13g2_nor2_1 _5808_ (.A(_1898_),
    .B(_1957_),
    .Y(_1958_));
 sg13g2_xor2_1 _5809_ (.B(_1886_),
    .A(_1877_),
    .X(_1959_));
 sg13g2_o21ai_1 _5810_ (.B1(_1887_),
    .Y(_1960_),
    .A1(_1958_),
    .A2(_1959_));
 sg13g2_o21ai_1 _5811_ (.B1(_1884_),
    .Y(_1961_),
    .A1(_3124_),
    .A2(_1885_));
 sg13g2_a21oi_1 _5812_ (.A1(\vgademo.linelfsr[11] ),
    .A2(_1882_),
    .Y(_1962_),
    .B1(_1880_));
 sg13g2_xnor2_1 _5813_ (.Y(_1963_),
    .A(\vgademo.linelfsr[12] ),
    .B(net982));
 sg13g2_nand2_1 _5814_ (.Y(_1964_),
    .A(net983),
    .B(net1063));
 sg13g2_xnor2_1 _5815_ (.Y(_1965_),
    .A(_1879_),
    .B(_1964_));
 sg13g2_xnor2_1 _5816_ (.Y(_1966_),
    .A(_1963_),
    .B(_1965_));
 sg13g2_xnor2_1 _5817_ (.Y(_1967_),
    .A(_1962_),
    .B(_1966_));
 sg13g2_xnor2_1 _5818_ (.Y(_1968_),
    .A(_1961_),
    .B(_1967_));
 sg13g2_xnor2_1 _5819_ (.Y(_1969_),
    .A(_1960_),
    .B(_1968_));
 sg13g2_inv_1 _5820_ (.Y(_1970_),
    .A(_1969_));
 sg13g2_xor2_1 _5821_ (.B(_1959_),
    .A(_1958_),
    .X(_1971_));
 sg13g2_inv_1 _5822_ (.Y(_1972_),
    .A(_1971_));
 sg13g2_xor2_1 _5823_ (.B(_1956_),
    .A(_1899_),
    .X(_1973_));
 sg13g2_xor2_1 _5824_ (.B(_1954_),
    .A(_1922_),
    .X(_1974_));
 sg13g2_inv_1 _5825_ (.Y(_1975_),
    .A(_1974_));
 sg13g2_xor2_1 _5826_ (.B(_1931_),
    .A(_1930_),
    .X(_1976_));
 sg13g2_xor2_1 _5827_ (.B(_1976_),
    .A(_1953_),
    .X(_1977_));
 sg13g2_xnor2_1 _5828_ (.Y(_1978_),
    .A(_1946_),
    .B(_1949_));
 sg13g2_xor2_1 _5829_ (.B(net1004),
    .A(\vgademo.linelfsr[3] ),
    .X(_1979_));
 sg13g2_xnor2_1 _5830_ (.Y(_1980_),
    .A(\vgademo.linelfsr[3] ),
    .B(net1004));
 sg13g2_nor2_2 _5831_ (.A(_1947_),
    .B(_1980_),
    .Y(_1981_));
 sg13g2_nand2_1 _5832_ (.Y(_1982_),
    .A(_1978_),
    .B(_1981_));
 sg13g2_xnor2_1 _5833_ (.Y(_1983_),
    .A(_1950_),
    .B(_1951_));
 sg13g2_nor2b_1 _5834_ (.A(_1982_),
    .B_N(_1983_),
    .Y(_1984_));
 sg13g2_nand3_1 _5835_ (.B(_1977_),
    .C(_1984_),
    .A(_1974_),
    .Y(_1985_));
 sg13g2_nand2b_1 _5836_ (.Y(_1986_),
    .B(_1911_),
    .A_N(_1910_));
 sg13g2_xnor2_1 _5837_ (.Y(_1987_),
    .A(_1955_),
    .B(_1986_));
 sg13g2_nor2_1 _5838_ (.A(_1985_),
    .B(_1987_),
    .Y(_1988_));
 sg13g2_nor2b_1 _5839_ (.A(_1973_),
    .B_N(_1988_),
    .Y(_1989_));
 sg13g2_xor2_1 _5840_ (.B(_1988_),
    .A(_1973_),
    .X(_1990_));
 sg13g2_xnor2_1 _5841_ (.Y(_1991_),
    .A(_1978_),
    .B(_1981_));
 sg13g2_xor2_1 _5842_ (.B(_1948_),
    .A(_1947_),
    .X(_1992_));
 sg13g2_nor2_1 _5843_ (.A(_1979_),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_nor3_1 _5844_ (.A(net1023),
    .B(_1981_),
    .C(_1993_),
    .Y(_1994_));
 sg13g2_o21ai_1 _5845_ (.B1(net1023),
    .Y(_1995_),
    .A1(_1981_),
    .A2(_1993_));
 sg13g2_nor2b_1 _5846_ (.A(_1994_),
    .B_N(_1995_),
    .Y(_1996_));
 sg13g2_xnor2_1 _5847_ (.Y(_1997_),
    .A(net1027),
    .B(_1979_));
 sg13g2_nand2b_1 _5848_ (.Y(_1998_),
    .B(\vgademo.linelfsr[2] ),
    .A_N(\vgademo.audio_snare_frames[1] ));
 sg13g2_nor2_1 _5849_ (.A(_1997_),
    .B(_1998_),
    .Y(_1999_));
 sg13g2_a21oi_1 _5850_ (.A1(_3147_),
    .A2(_1980_),
    .Y(_2000_),
    .B1(_1999_));
 sg13g2_nand2b_1 _5851_ (.Y(_2001_),
    .B(_1996_),
    .A_N(_2000_));
 sg13g2_nor2b_1 _5852_ (.A(_1994_),
    .B_N(_2001_),
    .Y(_2002_));
 sg13g2_or2_1 _5853_ (.X(_2003_),
    .B(_2002_),
    .A(_1991_));
 sg13g2_nor3_2 _5854_ (.A(_1951_),
    .B(_1976_),
    .C(_2003_),
    .Y(_2004_));
 sg13g2_a21o_1 _5855_ (.A2(_1984_),
    .A1(_1977_),
    .B1(_1974_),
    .X(_2005_));
 sg13g2_and2_1 _5856_ (.A(_1985_),
    .B(_2005_),
    .X(_2006_));
 sg13g2_nand2_1 _5857_ (.Y(_2007_),
    .A(_1922_),
    .B(_2004_));
 sg13g2_or2_1 _5858_ (.X(_2008_),
    .B(_2007_),
    .A(_1986_));
 sg13g2_nor2_1 _5859_ (.A(_1990_),
    .B(_2008_),
    .Y(_2009_));
 sg13g2_or2_1 _5860_ (.X(_2010_),
    .B(_2009_),
    .A(_1989_));
 sg13g2_nand2_1 _5861_ (.Y(_2011_),
    .A(_1971_),
    .B(_2010_));
 sg13g2_nor2_1 _5862_ (.A(_1970_),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_a21oi_1 _5863_ (.A1(_1971_),
    .A2(_1989_),
    .Y(_2013_),
    .B1(_1969_));
 sg13g2_nor2_1 _5864_ (.A(_2012_),
    .B(_2013_),
    .Y(_2014_));
 sg13g2_nand2_1 _5865_ (.Y(_2015_),
    .A(\vgademo.h_count[10] ),
    .B(_2014_));
 sg13g2_xnor2_1 _5866_ (.Y(_2016_),
    .A(_1971_),
    .B(_2010_));
 sg13g2_xnor2_1 _5867_ (.Y(_2017_),
    .A(_0039_),
    .B(_2016_));
 sg13g2_xor2_1 _5868_ (.B(_2008_),
    .A(_1990_),
    .X(_2018_));
 sg13g2_nand2_1 _5869_ (.Y(_2019_),
    .A(_0038_),
    .B(_2018_));
 sg13g2_nand2_1 _5870_ (.Y(_2020_),
    .A(_1982_),
    .B(_2003_));
 sg13g2_nand2_1 _5871_ (.Y(_2021_),
    .A(_1983_),
    .B(_2020_));
 sg13g2_xnor2_1 _5872_ (.Y(_2022_),
    .A(_0035_),
    .B(_1977_));
 sg13g2_xor2_1 _5873_ (.B(_2022_),
    .A(_2021_),
    .X(_2023_));
 sg13g2_xor2_1 _5874_ (.B(_2020_),
    .A(_1983_),
    .X(_2024_));
 sg13g2_xnor2_1 _5875_ (.Y(_2025_),
    .A(_1991_),
    .B(_2002_));
 sg13g2_xnor2_1 _5876_ (.Y(_2026_),
    .A(_1996_),
    .B(_2000_));
 sg13g2_nor2_1 _5877_ (.A(net1014),
    .B(_1997_),
    .Y(_2027_));
 sg13g2_nor2b_1 _5878_ (.A(\vgademo.linelfsr[2] ),
    .B_N(\vgademo.audio_snare_frames[1] ),
    .Y(_2028_));
 sg13g2_a21oi_1 _5879_ (.A1(\vgademo.h_count[0] ),
    .A2(_1998_),
    .Y(_2029_),
    .B1(_2028_));
 sg13g2_a21oi_1 _5880_ (.A1(net1014),
    .A2(_1997_),
    .Y(_2030_),
    .B1(_1999_));
 sg13g2_o21ai_1 _5881_ (.B1(_2030_),
    .Y(_2031_),
    .A1(_2027_),
    .A2(_2029_));
 sg13g2_a21oi_1 _5882_ (.A1(_0033_),
    .A2(_2031_),
    .Y(_2032_),
    .B1(net1012));
 sg13g2_nand3b_1 _5883_ (.B(_2026_),
    .C(_2031_),
    .Y(_2033_),
    .A_N(_0033_));
 sg13g2_o21ai_1 _5884_ (.B1(_2033_),
    .Y(_2034_),
    .A1(_2026_),
    .A2(_2032_));
 sg13g2_a21o_1 _5885_ (.A2(_2034_),
    .A1(_2025_),
    .B1(net1010),
    .X(_2035_));
 sg13g2_o21ai_1 _5886_ (.B1(_2035_),
    .Y(_2036_),
    .A1(_2025_),
    .A2(_2034_));
 sg13g2_o21ai_1 _5887_ (.B1(_2036_),
    .Y(_2037_),
    .A1(_0044_),
    .A2(_2024_));
 sg13g2_nand2_1 _5888_ (.Y(_2038_),
    .A(_0044_),
    .B(_2024_));
 sg13g2_nand3_1 _5889_ (.B(_2037_),
    .C(_2038_),
    .A(_2023_),
    .Y(_2039_));
 sg13g2_xnor2_1 _5890_ (.Y(_2040_),
    .A(_1977_),
    .B(_2021_));
 sg13g2_o21ai_1 _5891_ (.B1(_2039_),
    .Y(_2041_),
    .A1(net957),
    .A2(_2040_));
 sg13g2_xnor2_1 _5892_ (.Y(_2042_),
    .A(_2004_),
    .B(_2006_));
 sg13g2_xnor2_1 _5893_ (.Y(_2043_),
    .A(_0036_),
    .B(_2042_));
 sg13g2_a22oi_1 _5894_ (.Y(_2044_),
    .B1(_2043_),
    .B2(_2041_),
    .A2(_2042_),
    .A1(net1008));
 sg13g2_nand2_1 _5895_ (.Y(_2045_),
    .A(_1985_),
    .B(_2007_));
 sg13g2_xnor2_1 _5896_ (.Y(_2046_),
    .A(_1987_),
    .B(_2045_));
 sg13g2_a21oi_1 _5897_ (.A1(_3120_),
    .A2(_2046_),
    .Y(_2047_),
    .B1(_2044_));
 sg13g2_nor2_1 _5898_ (.A(_3120_),
    .B(_2046_),
    .Y(_2048_));
 sg13g2_o21ai_1 _5899_ (.B1(_2019_),
    .Y(_2049_),
    .A1(_2047_),
    .A2(_2048_));
 sg13g2_o21ai_1 _5900_ (.B1(_2049_),
    .Y(_2050_),
    .A1(_0038_),
    .A2(_2018_));
 sg13g2_a22oi_1 _5901_ (.Y(_2051_),
    .B1(_2017_),
    .B2(_2050_),
    .A2(_2016_),
    .A1(\vgademo.h_count[9] ));
 sg13g2_xor2_1 _5902_ (.B(_2014_),
    .A(net1006),
    .X(_2052_));
 sg13g2_o21ai_1 _5903_ (.B1(_2015_),
    .Y(_2053_),
    .A1(_2051_),
    .A2(_2052_));
 sg13g2_o21ai_1 _5904_ (.B1(_2053_),
    .Y(_2054_),
    .A1(_1969_),
    .A2(_2011_));
 sg13g2_nor2_1 _5905_ (.A(\vgademo.h_count[7] ),
    .B(_1987_),
    .Y(_2055_));
 sg13g2_nor2_1 _5906_ (.A(net957),
    .B(_1977_),
    .Y(_2056_));
 sg13g2_or2_1 _5907_ (.X(_2057_),
    .B(_1983_),
    .A(_0044_));
 sg13g2_nor2_1 _5908_ (.A(_3117_),
    .B(_1992_),
    .Y(_2058_));
 sg13g2_xnor2_1 _5909_ (.Y(_2059_),
    .A(_0033_),
    .B(_1992_));
 sg13g2_a22oi_1 _5910_ (.Y(_2060_),
    .B1(_1979_),
    .B2(_3114_),
    .A2(_3115_),
    .A1(\vgademo.linelfsr[2] ));
 sg13g2_a21oi_1 _5911_ (.A1(net1014),
    .A2(_1980_),
    .Y(_2061_),
    .B1(_2060_));
 sg13g2_nand2b_1 _5912_ (.Y(_2062_),
    .B(net1010),
    .A_N(_1978_));
 sg13g2_o21ai_1 _5913_ (.B1(_2062_),
    .Y(_2063_),
    .A1(_2059_),
    .A2(_2061_));
 sg13g2_nand2b_1 _5914_ (.Y(_2064_),
    .B(_1978_),
    .A_N(net1010));
 sg13g2_o21ai_1 _5915_ (.B1(_2064_),
    .Y(_2065_),
    .A1(_2058_),
    .A2(_2063_));
 sg13g2_a21o_1 _5916_ (.A2(_1983_),
    .A1(_0044_),
    .B1(_2065_),
    .X(_2066_));
 sg13g2_a21oi_1 _5917_ (.A1(_2057_),
    .A2(_2066_),
    .Y(_2067_),
    .B1(_2022_));
 sg13g2_xor2_1 _5918_ (.B(_1974_),
    .A(_0036_),
    .X(_2068_));
 sg13g2_o21ai_1 _5919_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_2056_),
    .A2(_2067_));
 sg13g2_a22oi_1 _5920_ (.Y(_2070_),
    .B1(_1987_),
    .B2(\vgademo.h_count[7] ),
    .A2(_1975_),
    .A1(net1008));
 sg13g2_a21oi_1 _5921_ (.A1(_2069_),
    .A2(_2070_),
    .Y(_2071_),
    .B1(_2055_));
 sg13g2_xnor2_1 _5922_ (.Y(_2072_),
    .A(_0038_),
    .B(_1973_));
 sg13g2_a22oi_1 _5923_ (.Y(_2073_),
    .B1(_2071_),
    .B2(_2072_),
    .A2(_1973_),
    .A1(net1007));
 sg13g2_a21oi_1 _5924_ (.A1(_3121_),
    .A2(_1971_),
    .Y(_2074_),
    .B1(_2073_));
 sg13g2_a21oi_1 _5925_ (.A1(\vgademo.h_count[9] ),
    .A2(_1972_),
    .Y(_2075_),
    .B1(_2074_));
 sg13g2_o21ai_1 _5926_ (.B1(_2075_),
    .Y(_2076_),
    .A1(net1006),
    .A2(_1970_));
 sg13g2_nand2_1 _5927_ (.Y(_2077_),
    .A(net1006),
    .B(_1970_));
 sg13g2_nor2_1 _5928_ (.A(\vgademo.v_count[8] ),
    .B(net989),
    .Y(_2078_));
 sg13g2_nor2_1 _5929_ (.A(net973),
    .B(net985),
    .Y(_2079_));
 sg13g2_xnor2_1 _5930_ (.Y(_2080_),
    .A(net973),
    .B(net985));
 sg13g2_nand2b_1 _5931_ (.Y(_2081_),
    .B(_2080_),
    .A_N(_2078_));
 sg13g2_nand2_1 _5932_ (.Y(_2082_),
    .A(net974),
    .B(\vgademo.a_scrolly[8] ));
 sg13g2_xor2_1 _5933_ (.B(net989),
    .A(\vgademo.v_count[8] ),
    .X(_2083_));
 sg13g2_or2_1 _5934_ (.X(_2084_),
    .B(_2083_),
    .A(_2082_));
 sg13g2_xnor2_1 _5935_ (.Y(_2085_),
    .A(net974),
    .B(net991));
 sg13g2_nor2_1 _5936_ (.A(net975),
    .B(net994),
    .Y(_2086_));
 sg13g2_nor2_1 _5937_ (.A(_2085_),
    .B(_2086_),
    .Y(_2087_));
 sg13g2_nor2_1 _5938_ (.A(net976),
    .B(net996),
    .Y(_2088_));
 sg13g2_xor2_1 _5939_ (.B(net994),
    .A(net975),
    .X(_2089_));
 sg13g2_nor2_1 _5940_ (.A(_2088_),
    .B(_2089_),
    .Y(_2090_));
 sg13g2_or2_1 _5941_ (.X(_2091_),
    .B(net1000),
    .A(net978));
 sg13g2_xnor2_1 _5942_ (.Y(_2092_),
    .A(net976),
    .B(net996));
 sg13g2_or2_1 _5943_ (.X(_2093_),
    .B(_2092_),
    .A(_2091_));
 sg13g2_xnor2_1 _5944_ (.Y(_2094_),
    .A(net978),
    .B(net999));
 sg13g2_o21ai_1 _5945_ (.B1(_2094_),
    .Y(_2095_),
    .A1(\vgademo.v_count[3] ),
    .A2(net1002));
 sg13g2_a21oi_1 _5946_ (.A1(\vgademo.v_count[3] ),
    .A2(net1002),
    .Y(_2096_),
    .B1(_2094_));
 sg13g2_a21o_1 _5947_ (.A2(_3123_),
    .A1(_3111_),
    .B1(_2096_),
    .X(_2097_));
 sg13g2_nand2_1 _5948_ (.Y(_2098_),
    .A(_2093_),
    .B(_2095_));
 sg13g2_nor2b_1 _5949_ (.A(_2095_),
    .B_N(_2093_),
    .Y(_2099_));
 sg13g2_a21oi_1 _5950_ (.A1(_2091_),
    .A2(_2092_),
    .Y(_2100_),
    .B1(_2099_));
 sg13g2_o21ai_1 _5951_ (.B1(_2100_),
    .Y(_2101_),
    .A1(_2097_),
    .A2(_2098_));
 sg13g2_nand2_1 _5952_ (.Y(_2102_),
    .A(_2088_),
    .B(_2089_));
 sg13g2_nand2b_1 _5953_ (.Y(_2103_),
    .B(_2102_),
    .A_N(_2090_));
 sg13g2_a21oi_1 _5954_ (.A1(_2101_),
    .A2(_2102_),
    .Y(_2104_),
    .B1(_2090_));
 sg13g2_xnor2_1 _5955_ (.Y(_2105_),
    .A(_2085_),
    .B(_2086_));
 sg13g2_nor2_1 _5956_ (.A(_2104_),
    .B(_2105_),
    .Y(_2106_));
 sg13g2_nor2_2 _5957_ (.A(_2087_),
    .B(_2106_),
    .Y(_2107_));
 sg13g2_xnor2_1 _5958_ (.Y(_2108_),
    .A(_2082_),
    .B(_2083_));
 sg13g2_o21ai_1 _5959_ (.B1(_2084_),
    .Y(_2109_),
    .A1(_2107_),
    .A2(_2108_));
 sg13g2_xor2_1 _5960_ (.B(_2080_),
    .A(_2078_),
    .X(_2110_));
 sg13g2_nand2b_1 _5961_ (.Y(_2111_),
    .B(_2109_),
    .A_N(_2110_));
 sg13g2_xnor2_1 _5962_ (.Y(_2112_),
    .A(_3124_),
    .B(_2079_));
 sg13g2_a21oi_2 _5963_ (.B1(_2112_),
    .Y(_2113_),
    .A2(_2111_),
    .A1(_2081_));
 sg13g2_nor2_1 _5964_ (.A(_0019_),
    .B(_2079_),
    .Y(_2114_));
 sg13g2_nor2_1 _5965_ (.A(_2113_),
    .B(_2114_),
    .Y(_2115_));
 sg13g2_nand2b_1 _5966_ (.Y(_2116_),
    .B(_2115_),
    .A_N(net981));
 sg13g2_nor4_2 _5967_ (.A(net981),
    .B(\vgademo.a_scrolly[13] ),
    .C(_2113_),
    .Y(_2117_),
    .D(_2114_));
 sg13g2_a21oi_2 _5968_ (.B1(_2117_),
    .Y(_2118_),
    .A2(_2116_),
    .A1(\vgademo.a_scrolly[13] ));
 sg13g2_a21o_1 _5969_ (.A2(_2116_),
    .A1(net980),
    .B1(_2117_),
    .X(_2119_));
 sg13g2_and3_1 _5970_ (.X(_2120_),
    .A(_2081_),
    .B(_2111_),
    .C(_2112_));
 sg13g2_xor2_1 _5971_ (.B(_2110_),
    .A(_2109_),
    .X(_2121_));
 sg13g2_xor2_1 _5972_ (.B(_2108_),
    .A(_2107_),
    .X(_2122_));
 sg13g2_xor2_1 _5973_ (.B(_2105_),
    .A(_2104_),
    .X(_2123_));
 sg13g2_xnor2_1 _5974_ (.Y(_2124_),
    .A(_2101_),
    .B(_2103_));
 sg13g2_nand3_1 _5975_ (.B(_2123_),
    .C(_2124_),
    .A(_2122_),
    .Y(_2125_));
 sg13g2_xor2_1 _5976_ (.B(_2115_),
    .A(_0067_),
    .X(_2126_));
 sg13g2_nand2_1 _5977_ (.Y(_2127_),
    .A(_2118_),
    .B(_2126_));
 sg13g2_nor2b_1 _5978_ (.A(net980),
    .B_N(_2116_),
    .Y(_2128_));
 sg13g2_xnor2_1 _5979_ (.Y(_2129_),
    .A(_0066_),
    .B(_2128_));
 sg13g2_inv_1 _5980_ (.Y(_2130_),
    .A(_2129_));
 sg13g2_nand2_1 _5981_ (.Y(_2131_),
    .A(_2118_),
    .B(_2121_));
 sg13g2_o21ai_1 _5982_ (.B1(_2118_),
    .Y(_2132_),
    .A1(_2113_),
    .A2(_2120_));
 sg13g2_o21ai_1 _5983_ (.B1(_2118_),
    .Y(_2133_),
    .A1(_2121_),
    .A2(_2125_));
 sg13g2_nand4_1 _5984_ (.B(_2129_),
    .C(_2132_),
    .A(_2127_),
    .Y(_2134_),
    .D(_2133_));
 sg13g2_nand4_1 _5985_ (.B(_2076_),
    .C(_2077_),
    .A(_2054_),
    .Y(_2135_),
    .D(_2134_));
 sg13g2_inv_1 _5986_ (.Y(_2136_),
    .A(_2135_));
 sg13g2_nor4_1 _5987_ (.A(net1004),
    .B(_1020_),
    .C(_1184_),
    .D(_1343_),
    .Y(_2137_));
 sg13g2_a21oi_1 _5988_ (.A1(_3127_),
    .A2(_1183_),
    .Y(_2138_),
    .B1(_2137_));
 sg13g2_a21oi_1 _5989_ (.A1(_0066_),
    .A2(_2137_),
    .Y(_2139_),
    .B1(_2138_));
 sg13g2_and2_2 _5990_ (.A(_1025_),
    .B(_2139_),
    .X(_2140_));
 sg13g2_nand2_1 _5991_ (.Y(_2141_),
    .A(_0078_),
    .B(_2140_));
 sg13g2_a21oi_2 _5992_ (.B1(net871),
    .Y(_2142_),
    .A2(_2141_),
    .A1(_2135_));
 sg13g2_nor2_2 _5993_ (.A(_2130_),
    .B(_2140_),
    .Y(_2143_));
 sg13g2_nor3_1 _5994_ (.A(net871),
    .B(_2130_),
    .C(_2140_),
    .Y(_2144_));
 sg13g2_a221oi_1 _5995_ (.B2(_2144_),
    .C1(_2142_),
    .B1(_2127_),
    .A1(net834),
    .Y(_2145_),
    .A2(_1863_));
 sg13g2_or2_1 _5996_ (.X(_2146_),
    .B(_2145_),
    .A(_1756_));
 sg13g2_nor2_1 _5997_ (.A(net856),
    .B(_1543_),
    .Y(_2147_));
 sg13g2_xnor2_1 _5998_ (.Y(_2148_),
    .A(net856),
    .B(_1542_));
 sg13g2_nor2_1 _5999_ (.A(net855),
    .B(net862),
    .Y(_2149_));
 sg13g2_a21oi_1 _6000_ (.A1(_2148_),
    .A2(_2149_),
    .Y(_2150_),
    .B1(_2147_));
 sg13g2_xnor2_1 _6001_ (.Y(_2151_),
    .A(_1442_),
    .B(_1565_));
 sg13g2_xnor2_1 _6002_ (.Y(_2152_),
    .A(_2150_),
    .B(_2151_));
 sg13g2_inv_1 _6003_ (.Y(_2153_),
    .A(_2152_));
 sg13g2_a21oi_2 _6004_ (.B1(net879),
    .Y(_2154_),
    .A2(_2153_),
    .A1(_1756_));
 sg13g2_o21ai_1 _6005_ (.B1(_1275_),
    .Y(_2155_),
    .A1(net836),
    .A2(_2152_));
 sg13g2_xnor2_1 _6006_ (.Y(_2156_),
    .A(net861),
    .B(net862));
 sg13g2_a21o_1 _6007_ (.A2(_2156_),
    .A1(_2148_),
    .B1(net879),
    .X(_2157_));
 sg13g2_nand2_2 _6008_ (.Y(_2158_),
    .A(_2155_),
    .B(_2157_));
 sg13g2_a21oi_2 _6009_ (.B1(_1298_),
    .Y(_2159_),
    .A2(_2158_),
    .A1(_2146_));
 sg13g2_a21o_1 _6010_ (.A2(_2158_),
    .A1(_2146_),
    .B1(_1298_),
    .X(_2160_));
 sg13g2_and3_2 _6011_ (.X(_2161_),
    .A(_1789_),
    .B(_1808_),
    .C(_1858_));
 sg13g2_a21o_2 _6012_ (.A2(_1859_),
    .A1(_0055_),
    .B1(_1852_),
    .X(_2162_));
 sg13g2_nor2_1 _6013_ (.A(_2161_),
    .B(_2162_),
    .Y(_2163_));
 sg13g2_nor2_1 _6014_ (.A(net866),
    .B(_2163_),
    .Y(_2164_));
 sg13g2_and2_1 _6015_ (.A(net834),
    .B(_2164_),
    .X(_2165_));
 sg13g2_a21oi_1 _6016_ (.A1(_0075_),
    .A2(_2140_),
    .Y(_2166_),
    .B1(_2136_));
 sg13g2_nand2_1 _6017_ (.Y(_2167_),
    .A(_2132_),
    .B(_2143_));
 sg13g2_a21oi_1 _6018_ (.A1(_2166_),
    .A2(_2167_),
    .Y(_2168_),
    .B1(net871));
 sg13g2_o21ai_1 _6019_ (.B1(net835),
    .Y(_2169_),
    .A1(_2165_),
    .A2(_2168_));
 sg13g2_nand2_2 _6020_ (.Y(_2170_),
    .A(_2158_),
    .B(_2169_));
 sg13g2_xor2_1 _6021_ (.B(\vgademo.a_scrolly[3] ),
    .A(\vgademo.h_count[0] ),
    .X(_2171_));
 sg13g2_xnor2_1 _6022_ (.Y(_2172_),
    .A(net979),
    .B(net953));
 sg13g2_xnor2_1 _6023_ (.Y(_2173_),
    .A(_3109_),
    .B(net953));
 sg13g2_nand3_1 _6024_ (.B(_2169_),
    .C(_2172_),
    .A(_2158_),
    .Y(_2174_));
 sg13g2_a21oi_1 _6025_ (.A1(_2170_),
    .A2(_2173_),
    .Y(_2175_),
    .B1(_2159_));
 sg13g2_a21o_1 _6026_ (.A2(_2174_),
    .A1(_2159_),
    .B1(_2175_),
    .X(_2176_));
 sg13g2_nand2_1 _6027_ (.Y(_2177_),
    .A(_1275_),
    .B(_2156_));
 sg13g2_xor2_1 _6028_ (.B(_2149_),
    .A(_2148_),
    .X(_2178_));
 sg13g2_nand2b_1 _6029_ (.Y(_2179_),
    .B(_1756_),
    .A_N(_2178_));
 sg13g2_and2_1 _6030_ (.A(_2154_),
    .B(_2179_),
    .X(_2180_));
 sg13g2_nor2_1 _6031_ (.A(_2152_),
    .B(_2178_),
    .Y(_2181_));
 sg13g2_a22oi_1 _6032_ (.Y(_2182_),
    .B1(_2181_),
    .B2(_1275_),
    .A2(_2179_),
    .A1(_2154_));
 sg13g2_nor3_2 _6033_ (.A(_1789_),
    .B(_1808_),
    .C(_1859_),
    .Y(_2183_));
 sg13g2_nor2_2 _6034_ (.A(_1810_),
    .B(_1859_),
    .Y(_2184_));
 sg13g2_inv_1 _6035_ (.Y(_2185_),
    .A(_2184_));
 sg13g2_and3_1 _6036_ (.X(_2186_),
    .A(_1781_),
    .B(_1782_),
    .C(_1785_));
 sg13g2_nor3_1 _6037_ (.A(_1786_),
    .B(_2185_),
    .C(_2186_),
    .Y(_2187_));
 sg13g2_a21o_2 _6038_ (.A2(_1859_),
    .A1(_0057_),
    .B1(_1852_),
    .X(_2188_));
 sg13g2_nor2_1 _6039_ (.A(_2187_),
    .B(_2188_),
    .Y(_2189_));
 sg13g2_mux2_1 _6040_ (.A0(_1862_),
    .A1(_2189_),
    .S(net834),
    .X(_2190_));
 sg13g2_nand2_1 _6041_ (.Y(_2191_),
    .A(_0056_),
    .B(_2140_));
 sg13g2_a21oi_2 _6042_ (.B1(net871),
    .Y(_2192_),
    .A2(_2191_),
    .A1(_2135_));
 sg13g2_a21oi_1 _6043_ (.A1(_2131_),
    .A2(_2144_),
    .Y(_2193_),
    .B1(_2192_));
 sg13g2_o21ai_1 _6044_ (.B1(_2193_),
    .Y(_2194_),
    .A1(net866),
    .A2(_2190_));
 sg13g2_a22oi_1 _6045_ (.Y(_2195_),
    .B1(_2194_),
    .B2(net835),
    .A2(_2182_),
    .A1(_2177_));
 sg13g2_nor2b_1 _6046_ (.A(_2195_),
    .B_N(net953),
    .Y(_2196_));
 sg13g2_xnor2_1 _6047_ (.Y(_2197_),
    .A(net953),
    .B(_2195_));
 sg13g2_a21oi_1 _6048_ (.A1(_2170_),
    .A2(_2197_),
    .Y(_2198_),
    .B1(_2196_));
 sg13g2_xnor2_1 _6049_ (.Y(_2199_),
    .A(_2170_),
    .B(_2172_));
 sg13g2_xnor2_1 _6050_ (.Y(_2200_),
    .A(_2159_),
    .B(_2199_));
 sg13g2_or2_1 _6051_ (.X(_2201_),
    .B(_2200_),
    .A(_2198_));
 sg13g2_nand2_1 _6052_ (.Y(_2202_),
    .A(net866),
    .B(_2135_));
 sg13g2_nand2_2 _6053_ (.Y(_2203_),
    .A(net835),
    .B(_2202_));
 sg13g2_a21oi_1 _6054_ (.A1(_0064_),
    .A2(_2140_),
    .Y(_2204_),
    .B1(_2202_));
 sg13g2_or2_1 _6055_ (.X(_2205_),
    .B(_2204_),
    .A(_1756_));
 sg13g2_o21ai_1 _6056_ (.B1(_2143_),
    .Y(_2206_),
    .A1(_2119_),
    .A2(_2123_));
 sg13g2_nand2b_1 _6057_ (.Y(_2207_),
    .B(net835),
    .A_N(_2206_));
 sg13g2_or2_1 _6058_ (.X(_2208_),
    .B(_2189_),
    .A(net834));
 sg13g2_nor2_1 _6059_ (.A(net1005),
    .B(\vgademo.plane_du[4] ),
    .Y(_2209_));
 sg13g2_or3_1 _6060_ (.A(_1784_),
    .B(_2185_),
    .C(_2209_),
    .X(_2210_));
 sg13g2_a21oi_2 _6061_ (.B1(_1852_),
    .Y(_2211_),
    .A2(_1859_),
    .A1(_0059_));
 sg13g2_nand2_1 _6062_ (.Y(_2212_),
    .A(_2210_),
    .B(_2211_));
 sg13g2_a21oi_1 _6063_ (.A1(net832),
    .A2(_2212_),
    .Y(_2213_),
    .B1(_1322_));
 sg13g2_a22oi_1 _6064_ (.Y(_2214_),
    .B1(_2208_),
    .B2(_2213_),
    .A2(_2207_),
    .A1(_2205_));
 sg13g2_nor2_1 _6065_ (.A(net878),
    .B(_2214_),
    .Y(_2215_));
 sg13g2_inv_1 _6066_ (.Y(_2216_),
    .A(_2215_));
 sg13g2_a21o_1 _6067_ (.A2(_1783_),
    .A1(_1782_),
    .B1(_1784_),
    .X(_2217_));
 sg13g2_nand3_1 _6068_ (.B(_2184_),
    .C(_2217_),
    .A(_1785_),
    .Y(_2218_));
 sg13g2_a21o_2 _6069_ (.A2(_1859_),
    .A1(_0062_),
    .B1(_1852_),
    .X(_2219_));
 sg13g2_nor2b_1 _6070_ (.A(_2219_),
    .B_N(_2218_),
    .Y(_2220_));
 sg13g2_a21oi_2 _6071_ (.B1(_1852_),
    .Y(_2221_),
    .A2(_1859_),
    .A1(_0058_));
 sg13g2_inv_1 _6072_ (.Y(_2222_),
    .A(_2221_));
 sg13g2_a21oi_1 _6073_ (.A1(\vgademo.plane_du[3] ),
    .A2(_2184_),
    .Y(_2223_),
    .B1(_2222_));
 sg13g2_mux2_1 _6074_ (.A0(_2220_),
    .A1(_2223_),
    .S(net832),
    .X(_2224_));
 sg13g2_o21ai_1 _6075_ (.B1(_2143_),
    .Y(_2225_),
    .A1(_2119_),
    .A2(_2124_));
 sg13g2_nand2b_1 _6076_ (.Y(_2226_),
    .B(net835),
    .A_N(_2225_));
 sg13g2_a22oi_1 _6077_ (.Y(_2227_),
    .B1(_2226_),
    .B2(_2203_),
    .A2(_2224_),
    .A1(net871));
 sg13g2_nor2_1 _6078_ (.A(net878),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_xor2_1 _6079_ (.B(net1005),
    .A(net1015),
    .X(_2229_));
 sg13g2_nor2b_1 _6080_ (.A(_2228_),
    .B_N(net951),
    .Y(_2230_));
 sg13g2_o21ai_1 _6081_ (.B1(net951),
    .Y(_2231_),
    .A1(net878),
    .A2(_2227_));
 sg13g2_nor3_1 _6082_ (.A(net878),
    .B(_2227_),
    .C(net951),
    .Y(_2232_));
 sg13g2_xnor2_1 _6083_ (.Y(_2233_),
    .A(_2228_),
    .B(net951));
 sg13g2_xnor2_1 _6084_ (.Y(_2234_),
    .A(_2216_),
    .B(_2233_));
 sg13g2_a21o_1 _6085_ (.A2(_2140_),
    .A1(_0069_),
    .B1(_2202_),
    .X(_2235_));
 sg13g2_nand2_1 _6086_ (.Y(_2236_),
    .A(net835),
    .B(_2235_));
 sg13g2_o21ai_1 _6087_ (.B1(_2143_),
    .Y(_2237_),
    .A1(_2119_),
    .A2(_2122_));
 sg13g2_inv_1 _6088_ (.Y(_2238_),
    .A(_2237_));
 sg13g2_o21ai_1 _6089_ (.B1(net835),
    .Y(_2239_),
    .A1(_2235_),
    .A2(_2238_));
 sg13g2_mux2_1 _6090_ (.A0(_2163_),
    .A1(_2220_),
    .S(net834),
    .X(_2240_));
 sg13g2_a21o_1 _6091_ (.A2(_2240_),
    .A1(net871),
    .B1(_2239_),
    .X(_2241_));
 sg13g2_nand2_1 _6092_ (.Y(_2242_),
    .A(_2154_),
    .B(_2241_));
 sg13g2_xor2_1 _6093_ (.B(net1005),
    .A(net1013),
    .X(_2243_));
 sg13g2_inv_1 _6094_ (.Y(_2244_),
    .A(_2243_));
 sg13g2_o21ai_1 _6095_ (.B1(_2243_),
    .Y(_2245_),
    .A1(net878),
    .A2(_2214_));
 sg13g2_nor3_1 _6096_ (.A(net878),
    .B(_2214_),
    .C(_2243_),
    .Y(_2246_));
 sg13g2_a21oi_1 _6097_ (.A1(_2160_),
    .A2(_2245_),
    .Y(_2247_),
    .B1(_2246_));
 sg13g2_nand2_1 _6098_ (.Y(_2248_),
    .A(_2242_),
    .B(_2247_));
 sg13g2_a21oi_1 _6099_ (.A1(_2216_),
    .A2(_2233_),
    .Y(_2249_),
    .B1(_2230_));
 sg13g2_o21ai_1 _6100_ (.B1(_2231_),
    .Y(_2250_),
    .A1(_2215_),
    .A2(_2232_));
 sg13g2_xnor2_1 _6101_ (.Y(_2251_),
    .A(\vgademo.bayer_j[1] ),
    .B(net952));
 sg13g2_xor2_1 _6102_ (.B(net952),
    .A(\vgademo.bayer_j[1] ),
    .X(_2252_));
 sg13g2_a21oi_1 _6103_ (.A1(_2154_),
    .A2(_2241_),
    .Y(_2253_),
    .B1(_2251_));
 sg13g2_and3_1 _6104_ (.X(_2254_),
    .A(_2154_),
    .B(_2241_),
    .C(_2251_));
 sg13g2_or3_1 _6105_ (.A(_2195_),
    .B(_2253_),
    .C(_2254_),
    .X(_2255_));
 sg13g2_o21ai_1 _6106_ (.B1(_2195_),
    .Y(_2256_),
    .A1(_2253_),
    .A2(_2254_));
 sg13g2_nand2_1 _6107_ (.Y(_2257_),
    .A(_2255_),
    .B(_2256_));
 sg13g2_nor2_1 _6108_ (.A(_2242_),
    .B(_2247_),
    .Y(_2258_));
 sg13g2_a221oi_1 _6109_ (.B2(_2257_),
    .C1(_2258_),
    .B1(_2249_),
    .A1(_2234_),
    .Y(_2259_),
    .A2(_2248_));
 sg13g2_nand3_1 _6110_ (.B(_2255_),
    .C(_2256_),
    .A(_2250_),
    .Y(_2260_));
 sg13g2_nor2b_1 _6111_ (.A(_2253_),
    .B_N(_2255_),
    .Y(_2261_));
 sg13g2_xnor2_1 _6112_ (.Y(_2262_),
    .A(_2170_),
    .B(_2197_));
 sg13g2_o21ai_1 _6113_ (.B1(_2260_),
    .Y(_2263_),
    .A1(_2261_),
    .A2(_2262_));
 sg13g2_a22oi_1 _6114_ (.Y(_2264_),
    .B1(_2261_),
    .B2(_2262_),
    .A2(_2200_),
    .A1(_2198_));
 sg13g2_o21ai_1 _6115_ (.B1(_2264_),
    .Y(_2265_),
    .A1(_2259_),
    .A2(_2263_));
 sg13g2_a21oi_1 _6116_ (.A1(_2201_),
    .A2(_2265_),
    .Y(_2266_),
    .B1(_2176_));
 sg13g2_and3_1 _6117_ (.X(_2267_),
    .A(_2176_),
    .B(_2201_),
    .C(_2265_));
 sg13g2_nor4_1 _6118_ (.A(net1010),
    .B(net1012),
    .C(\vgademo.h_count[5] ),
    .D(net1009),
    .Y(_2268_));
 sg13g2_o21ai_1 _6119_ (.B1(_0579_),
    .Y(_2269_),
    .A1(_3203_),
    .A2(_2268_));
 sg13g2_nand2b_2 _6120_ (.Y(_2270_),
    .B(_2269_),
    .A_N(net1006));
 sg13g2_nor2_1 _6121_ (.A(\vgademo.v_count[3] ),
    .B(\vgademo.v_count[2] ),
    .Y(_2271_));
 sg13g2_nand4_1 _6122_ (.B(_3240_),
    .C(_3241_),
    .A(_3237_),
    .Y(_2272_),
    .D(_2271_));
 sg13g2_a21oi_1 _6123_ (.A1(\vgademo.v_count[8] ),
    .A2(_3235_),
    .Y(_2273_),
    .B1(\vgademo.v_count[9] ));
 sg13g2_nand3_1 _6124_ (.B(_2272_),
    .C(_2273_),
    .A(_2270_),
    .Y(_2274_));
 sg13g2_nor3_1 _6125_ (.A(_2266_),
    .B(_2267_),
    .C(_2274_),
    .Y(_0256_));
 sg13g2_a21oi_1 _6126_ (.A1(_2159_),
    .A2(_2174_),
    .Y(_2275_),
    .B1(_2266_));
 sg13g2_nor2_1 _6127_ (.A(_2274_),
    .B(_2275_),
    .Y(_0257_));
 sg13g2_nand2_1 _6128_ (.Y(_2276_),
    .A(\vgademo.a_sin[6] ),
    .B(net922));
 sg13g2_xnor2_1 _6129_ (.Y(_0258_),
    .A(net237),
    .B(_2276_));
 sg13g2_nor2_1 _6130_ (.A(net308),
    .B(net924),
    .Y(_2277_));
 sg13g2_nor2b_1 _6131_ (.A(\vgademo.a_sin[7] ),
    .B_N(\vgademo.a_cos[1] ),
    .Y(_2278_));
 sg13g2_xor2_1 _6132_ (.B(net308),
    .A(\vgademo.a_sin[7] ),
    .X(_2279_));
 sg13g2_nor2b_1 _6133_ (.A(net237),
    .B_N(\vgademo.a_sin[6] ),
    .Y(_2280_));
 sg13g2_nor2_1 _6134_ (.A(_2279_),
    .B(_2280_),
    .Y(_2281_));
 sg13g2_xnor2_1 _6135_ (.Y(_2282_),
    .A(_2279_),
    .B(_2280_));
 sg13g2_a21oi_1 _6136_ (.A1(net924),
    .A2(_2282_),
    .Y(_0259_),
    .B1(_2277_));
 sg13g2_nand2_1 _6137_ (.Y(_2283_),
    .A(_3164_),
    .B(net320));
 sg13g2_xnor2_1 _6138_ (.Y(_2284_),
    .A(\vgademo.a_sin[8] ),
    .B(\vgademo.a_cos[2] ));
 sg13g2_nor3_1 _6139_ (.A(_2278_),
    .B(_2281_),
    .C(_2284_),
    .Y(_2285_));
 sg13g2_o21ai_1 _6140_ (.B1(_2284_),
    .Y(_2286_),
    .A1(_2278_),
    .A2(_2281_));
 sg13g2_nor2b_1 _6141_ (.A(_2285_),
    .B_N(_2286_),
    .Y(_2287_));
 sg13g2_mux2_1 _6142_ (.A0(net320),
    .A1(_2287_),
    .S(net923),
    .X(_0260_));
 sg13g2_nand2_1 _6143_ (.Y(_2288_),
    .A(\vgademo.a_cos[3] ),
    .B(_3165_));
 sg13g2_xor2_1 _6144_ (.B(\vgademo.a_sin[9] ),
    .A(\vgademo.a_cos[3] ),
    .X(_2289_));
 sg13g2_nand3_1 _6145_ (.B(_2286_),
    .C(_2289_),
    .A(_2283_),
    .Y(_2290_));
 sg13g2_a21o_1 _6146_ (.A2(_2286_),
    .A1(_2283_),
    .B1(_2289_),
    .X(_2291_));
 sg13g2_nand3_1 _6147_ (.B(_2290_),
    .C(_2291_),
    .A(net923),
    .Y(_2292_));
 sg13g2_o21ai_1 _6148_ (.B1(_2292_),
    .Y(_0261_),
    .A1(_3149_),
    .A2(net923));
 sg13g2_nand2_1 _6149_ (.Y(_2293_),
    .A(net469),
    .B(net920));
 sg13g2_xor2_1 _6150_ (.B(\vgademo.a_sin[10] ),
    .A(\vgademo.a_cos[4] ),
    .X(_2294_));
 sg13g2_nand3_1 _6151_ (.B(_2291_),
    .C(_2294_),
    .A(_2288_),
    .Y(_2295_));
 sg13g2_a21oi_1 _6152_ (.A1(_2288_),
    .A2(_2291_),
    .Y(_2296_),
    .B1(_2294_));
 sg13g2_nand2_1 _6153_ (.Y(_2297_),
    .A(net923),
    .B(_2295_));
 sg13g2_o21ai_1 _6154_ (.B1(_2293_),
    .Y(_0262_),
    .A1(_2296_),
    .A2(_2297_));
 sg13g2_a21o_1 _6155_ (.A2(_3166_),
    .A1(\vgademo.a_cos[4] ),
    .B1(_2296_),
    .X(_2298_));
 sg13g2_nor2b_1 _6156_ (.A(\vgademo.a_sin[11] ),
    .B_N(\vgademo.a_cos[5] ),
    .Y(_2299_));
 sg13g2_nand2b_1 _6157_ (.Y(_2300_),
    .B(\vgademo.a_sin[11] ),
    .A_N(\vgademo.a_cos[5] ));
 sg13g2_nand2b_1 _6158_ (.Y(_2301_),
    .B(_2300_),
    .A_N(_2299_));
 sg13g2_xnor2_1 _6159_ (.Y(_2302_),
    .A(_2298_),
    .B(_2301_));
 sg13g2_mux2_1 _6160_ (.A0(net436),
    .A1(_2302_),
    .S(_0593_),
    .X(_0263_));
 sg13g2_xor2_1 _6161_ (.B(\vgademo.a_sin[12] ),
    .A(\vgademo.a_cos[6] ),
    .X(_2303_));
 sg13g2_a21oi_2 _6162_ (.B1(_2299_),
    .Y(_2304_),
    .A2(_2300_),
    .A1(_2298_));
 sg13g2_nor2_1 _6163_ (.A(_2303_),
    .B(_2304_),
    .Y(_2305_));
 sg13g2_xor2_1 _6164_ (.B(_2304_),
    .A(_2303_),
    .X(_2306_));
 sg13g2_and2_1 _6165_ (.A(net924),
    .B(_2306_),
    .X(_2307_));
 sg13g2_a21o_1 _6166_ (.A2(net919),
    .A1(net499),
    .B1(_2307_),
    .X(_0264_));
 sg13g2_a21oi_1 _6167_ (.A1(\vgademo.a_cos[6] ),
    .A2(_3167_),
    .Y(_2308_),
    .B1(_2305_));
 sg13g2_xnor2_1 _6168_ (.Y(_2309_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.a_sin[13] ));
 sg13g2_nand2b_1 _6169_ (.Y(_2310_),
    .B(_2309_),
    .A_N(_2308_));
 sg13g2_xnor2_1 _6170_ (.Y(_2311_),
    .A(_2308_),
    .B(_2309_));
 sg13g2_nor2_1 _6171_ (.A(net919),
    .B(_2311_),
    .Y(_2312_));
 sg13g2_a21oi_1 _6172_ (.A1(_3155_),
    .A2(net918),
    .Y(_0265_),
    .B1(_2312_));
 sg13g2_xnor2_1 _6173_ (.Y(_2313_),
    .A(\vgademo.a_cos[8] ),
    .B(net972));
 sg13g2_o21ai_1 _6174_ (.B1(_2310_),
    .Y(_2314_),
    .A1(_3155_),
    .A2(\vgademo.a_sin[13] ));
 sg13g2_and2_1 _6175_ (.A(_2313_),
    .B(_2314_),
    .X(_2315_));
 sg13g2_xor2_1 _6176_ (.B(_2314_),
    .A(_2313_),
    .X(_2316_));
 sg13g2_mux2_1 _6177_ (.A0(net555),
    .A1(_2316_),
    .S(net922),
    .X(_0266_));
 sg13g2_nor2_1 _6178_ (.A(net511),
    .B(net922),
    .Y(_2317_));
 sg13g2_xnor2_1 _6179_ (.Y(_2318_),
    .A(\vgademo.a_cos[9] ),
    .B(net972));
 sg13g2_a21oi_1 _6180_ (.A1(\vgademo.a_cos[8] ),
    .A2(_3168_),
    .Y(_2319_),
    .B1(_2315_));
 sg13g2_xor2_1 _6181_ (.B(_2319_),
    .A(_2318_),
    .X(_2320_));
 sg13g2_a21oi_1 _6182_ (.A1(net922),
    .A2(_2320_),
    .Y(_0267_),
    .B1(_2317_));
 sg13g2_nor2_1 _6183_ (.A(\vgademo.a_cos[10] ),
    .B(_3168_),
    .Y(_2321_));
 sg13g2_nand2_1 _6184_ (.Y(_2322_),
    .A(\vgademo.a_cos[10] ),
    .B(_3168_));
 sg13g2_nor2b_1 _6185_ (.A(_2321_),
    .B_N(_2322_),
    .Y(_2323_));
 sg13g2_and2_1 _6186_ (.A(_2315_),
    .B(_2318_),
    .X(_2324_));
 sg13g2_o21ai_1 _6187_ (.B1(_3168_),
    .Y(_2325_),
    .A1(\vgademo.a_cos[8] ),
    .A2(\vgademo.a_cos[9] ));
 sg13g2_nor2b_1 _6188_ (.A(_2324_),
    .B_N(_2325_),
    .Y(_2326_));
 sg13g2_xnor2_1 _6189_ (.Y(_2327_),
    .A(_2323_),
    .B(_2326_));
 sg13g2_mux2_1 _6190_ (.A0(net487),
    .A1(_2327_),
    .S(net925),
    .X(_0268_));
 sg13g2_nor2_1 _6191_ (.A(net466),
    .B(net925),
    .Y(_2328_));
 sg13g2_xnor2_1 _6192_ (.Y(_2329_),
    .A(\vgademo.a_cos[11] ),
    .B(net972));
 sg13g2_o21ai_1 _6193_ (.B1(_2322_),
    .Y(_2330_),
    .A1(_2321_),
    .A2(_2326_));
 sg13g2_xnor2_1 _6194_ (.Y(_2331_),
    .A(_2329_),
    .B(_2330_));
 sg13g2_a21oi_1 _6195_ (.A1(net925),
    .A2(_2331_),
    .Y(_0269_),
    .B1(_2328_));
 sg13g2_nor2b_1 _6196_ (.A(net972),
    .B_N(\vgademo.a_cos[12] ),
    .Y(_2332_));
 sg13g2_nand2b_1 _6197_ (.Y(_2333_),
    .B(net972),
    .A_N(\vgademo.a_cos[12] ));
 sg13g2_nand2b_1 _6198_ (.Y(_2334_),
    .B(_2333_),
    .A_N(_2332_));
 sg13g2_nand3_1 _6199_ (.B(_2324_),
    .C(_2329_),
    .A(_2323_),
    .Y(_2335_));
 sg13g2_o21ai_1 _6200_ (.B1(_3168_),
    .Y(_2336_),
    .A1(\vgademo.a_cos[10] ),
    .A2(\vgademo.a_cos[11] ));
 sg13g2_nand3_1 _6201_ (.B(_2335_),
    .C(_2336_),
    .A(_2325_),
    .Y(_2337_));
 sg13g2_xnor2_1 _6202_ (.Y(_2338_),
    .A(_2334_),
    .B(_2337_));
 sg13g2_mux2_1 _6203_ (.A0(net368),
    .A1(_2338_),
    .S(_0590_),
    .X(_0270_));
 sg13g2_nor2_1 _6204_ (.A(net232),
    .B(net922),
    .Y(_2339_));
 sg13g2_a21oi_2 _6205_ (.B1(_2332_),
    .Y(_2340_),
    .A2(_2337_),
    .A1(_2333_));
 sg13g2_nand2_1 _6206_ (.Y(_2341_),
    .A(\vgademo.a_cos[13] ),
    .B(_3168_));
 sg13g2_nor2_1 _6207_ (.A(\vgademo.a_cos[13] ),
    .B(_3168_),
    .Y(_2342_));
 sg13g2_xnor2_1 _6208_ (.Y(_2343_),
    .A(\vgademo.a_cos[13] ),
    .B(net972));
 sg13g2_xnor2_1 _6209_ (.Y(_2344_),
    .A(_2340_),
    .B(_2343_));
 sg13g2_a21oi_1 _6210_ (.A1(net922),
    .A2(_2344_),
    .Y(_0271_),
    .B1(_2339_));
 sg13g2_nand2_1 _6211_ (.Y(_2345_),
    .A(net472),
    .B(net918));
 sg13g2_o21ai_1 _6212_ (.B1(_2341_),
    .Y(_2346_),
    .A1(_2340_),
    .A2(_2342_));
 sg13g2_xnor2_1 _6213_ (.Y(_2347_),
    .A(\vgademo.a_cos[14] ),
    .B(net972));
 sg13g2_xnor2_1 _6214_ (.Y(_2348_),
    .A(_2346_),
    .B(_2347_));
 sg13g2_inv_1 _6215_ (.Y(_2349_),
    .A(net838));
 sg13g2_o21ai_1 _6216_ (.B1(_2345_),
    .Y(_0272_),
    .A1(net918),
    .A2(net838));
 sg13g2_xor2_1 _6217_ (.B(_2307_),
    .A(net215),
    .X(_0273_));
 sg13g2_nand2_1 _6218_ (.Y(_2350_),
    .A(net215),
    .B(_2306_));
 sg13g2_xnor2_1 _6219_ (.Y(_2351_),
    .A(\vgademo.a_sin[1] ),
    .B(_2311_));
 sg13g2_nor2_1 _6220_ (.A(_2350_),
    .B(_2351_),
    .Y(_2352_));
 sg13g2_nand2_1 _6221_ (.Y(_2353_),
    .A(net296),
    .B(net918));
 sg13g2_a21o_1 _6222_ (.A2(_2351_),
    .A1(_2350_),
    .B1(net918),
    .X(_2354_));
 sg13g2_o21ai_1 _6223_ (.B1(_2353_),
    .Y(_0274_),
    .A1(_2352_),
    .A2(_2354_));
 sg13g2_and2_1 _6224_ (.A(\vgademo.a_sin[2] ),
    .B(_2316_),
    .X(_2355_));
 sg13g2_xnor2_1 _6225_ (.Y(_2356_),
    .A(net295),
    .B(_2316_));
 sg13g2_a21oi_1 _6226_ (.A1(\vgademo.a_sin[1] ),
    .A2(_2311_),
    .Y(_2357_),
    .B1(_2352_));
 sg13g2_nor2_1 _6227_ (.A(_2356_),
    .B(_2357_),
    .Y(_2358_));
 sg13g2_nand2_1 _6228_ (.Y(_2359_),
    .A(net295),
    .B(net920));
 sg13g2_a21o_1 _6229_ (.A2(_2357_),
    .A1(_2356_),
    .B1(net920),
    .X(_2360_));
 sg13g2_o21ai_1 _6230_ (.B1(_2359_),
    .Y(_0275_),
    .A1(_2358_),
    .A2(_2360_));
 sg13g2_or2_1 _6231_ (.X(_2361_),
    .B(_2320_),
    .A(_3161_));
 sg13g2_xnor2_1 _6232_ (.Y(_2362_),
    .A(\vgademo.a_sin[3] ),
    .B(_2320_));
 sg13g2_o21ai_1 _6233_ (.B1(_2362_),
    .Y(_2363_),
    .A1(_2355_),
    .A2(_2358_));
 sg13g2_or3_1 _6234_ (.A(_2355_),
    .B(_2358_),
    .C(_2362_),
    .X(_2364_));
 sg13g2_a21oi_1 _6235_ (.A1(_2363_),
    .A2(_2364_),
    .Y(_2365_),
    .B1(net920));
 sg13g2_a21oi_1 _6236_ (.A1(_3161_),
    .A2(net920),
    .Y(_0276_),
    .B1(_2365_));
 sg13g2_and2_1 _6237_ (.A(\vgademo.a_sin[4] ),
    .B(_2327_),
    .X(_2366_));
 sg13g2_xnor2_1 _6238_ (.Y(_2367_),
    .A(\vgademo.a_sin[4] ),
    .B(_2327_));
 sg13g2_a21oi_1 _6239_ (.A1(_2361_),
    .A2(_2363_),
    .Y(_2368_),
    .B1(_2367_));
 sg13g2_nand3_1 _6240_ (.B(_2363_),
    .C(_2367_),
    .A(_2361_),
    .Y(_2369_));
 sg13g2_nand2_1 _6241_ (.Y(_2370_),
    .A(net346),
    .B(net920));
 sg13g2_nand2_1 _6242_ (.Y(_2371_),
    .A(net922),
    .B(_2369_));
 sg13g2_o21ai_1 _6243_ (.B1(_2370_),
    .Y(_0277_),
    .A1(_2368_),
    .A2(_2371_));
 sg13g2_nand2b_1 _6244_ (.Y(_2372_),
    .B(net341),
    .A_N(_2331_));
 sg13g2_xnor2_1 _6245_ (.Y(_2373_),
    .A(\vgademo.a_sin[5] ),
    .B(_2331_));
 sg13g2_o21ai_1 _6246_ (.B1(_2373_),
    .Y(_2374_),
    .A1(_2366_),
    .A2(_2368_));
 sg13g2_or3_1 _6247_ (.A(_2366_),
    .B(_2368_),
    .C(_2373_),
    .X(_2375_));
 sg13g2_a21oi_1 _6248_ (.A1(_2374_),
    .A2(_2375_),
    .Y(_2376_),
    .B1(net920));
 sg13g2_a21oi_1 _6249_ (.A1(_3162_),
    .A2(net920),
    .Y(_0278_),
    .B1(_2376_));
 sg13g2_and2_1 _6250_ (.A(\vgademo.a_sin[6] ),
    .B(_2338_),
    .X(_2377_));
 sg13g2_xnor2_1 _6251_ (.Y(_2378_),
    .A(\vgademo.a_sin[6] ),
    .B(_2338_));
 sg13g2_a21oi_1 _6252_ (.A1(_2372_),
    .A2(_2374_),
    .Y(_2379_),
    .B1(_2378_));
 sg13g2_nand3_1 _6253_ (.B(_2374_),
    .C(_2378_),
    .A(_2372_),
    .Y(_2380_));
 sg13g2_nand2_1 _6254_ (.Y(_2381_),
    .A(net429),
    .B(net918));
 sg13g2_nand2_1 _6255_ (.Y(_2382_),
    .A(net922),
    .B(_2380_));
 sg13g2_o21ai_1 _6256_ (.B1(_2381_),
    .Y(_0279_),
    .A1(_2379_),
    .A2(_2382_));
 sg13g2_nand2_1 _6257_ (.Y(_2383_),
    .A(\vgademo.a_sin[7] ),
    .B(_2344_));
 sg13g2_xnor2_1 _6258_ (.Y(_2384_),
    .A(_3163_),
    .B(_2344_));
 sg13g2_o21ai_1 _6259_ (.B1(_2384_),
    .Y(_2385_),
    .A1(_2377_),
    .A2(_2379_));
 sg13g2_or3_1 _6260_ (.A(_2377_),
    .B(_2379_),
    .C(_2384_),
    .X(_2386_));
 sg13g2_a21oi_1 _6261_ (.A1(_2385_),
    .A2(_2386_),
    .Y(_2387_),
    .B1(net918));
 sg13g2_a21oi_1 _6262_ (.A1(_3163_),
    .A2(net918),
    .Y(_0280_),
    .B1(_2387_));
 sg13g2_xnor2_1 _6263_ (.Y(_2388_),
    .A(_3164_),
    .B(net837));
 sg13g2_a21oi_1 _6264_ (.A1(_2383_),
    .A2(_2385_),
    .Y(_2389_),
    .B1(_2388_));
 sg13g2_nand3_1 _6265_ (.B(_2385_),
    .C(_2388_),
    .A(_2383_),
    .Y(_2390_));
 sg13g2_nand3b_1 _6266_ (.B(_2390_),
    .C(net923),
    .Y(_2391_),
    .A_N(_2389_));
 sg13g2_o21ai_1 _6267_ (.B1(_2391_),
    .Y(_0281_),
    .A1(_3164_),
    .A2(net923));
 sg13g2_nand2_1 _6268_ (.Y(_2392_),
    .A(net450),
    .B(net919));
 sg13g2_xnor2_1 _6269_ (.Y(_2393_),
    .A(\vgademo.a_sin[9] ),
    .B(net838));
 sg13g2_a21oi_1 _6270_ (.A1(net596),
    .A2(_2349_),
    .Y(_2394_),
    .B1(_2389_));
 sg13g2_xor2_1 _6271_ (.B(_2394_),
    .A(_2393_),
    .X(_2395_));
 sg13g2_o21ai_1 _6272_ (.B1(_2392_),
    .Y(_0282_),
    .A1(net919),
    .A2(_2395_));
 sg13g2_xnor2_1 _6273_ (.Y(_2396_),
    .A(\vgademo.a_sin[10] ),
    .B(net837));
 sg13g2_a21oi_1 _6274_ (.A1(_3164_),
    .A2(_3165_),
    .Y(_2397_),
    .B1(net837));
 sg13g2_and2_1 _6275_ (.A(_2389_),
    .B(_2393_),
    .X(_2398_));
 sg13g2_o21ai_1 _6276_ (.B1(_2396_),
    .Y(_2399_),
    .A1(_2397_),
    .A2(_2398_));
 sg13g2_or3_1 _6277_ (.A(_2396_),
    .B(_2397_),
    .C(_2398_),
    .X(_2400_));
 sg13g2_a21oi_1 _6278_ (.A1(_2399_),
    .A2(_2400_),
    .Y(_2401_),
    .B1(net919));
 sg13g2_a21oi_1 _6279_ (.A1(_3166_),
    .A2(net919),
    .Y(_0283_),
    .B1(_2401_));
 sg13g2_xnor2_1 _6280_ (.Y(_2402_),
    .A(\vgademo.a_sin[11] ),
    .B(net837));
 sg13g2_o21ai_1 _6281_ (.B1(_2399_),
    .Y(_2403_),
    .A1(_3166_),
    .A2(net837));
 sg13g2_o21ai_1 _6282_ (.B1(net923),
    .Y(_2404_),
    .A1(_2402_),
    .A2(_2403_));
 sg13g2_a21oi_1 _6283_ (.A1(_2402_),
    .A2(_2403_),
    .Y(_2405_),
    .B1(_2404_));
 sg13g2_a21o_1 _6284_ (.A2(net919),
    .A1(net491),
    .B1(_2405_),
    .X(_0284_));
 sg13g2_nor2_1 _6285_ (.A(net478),
    .B(net923),
    .Y(_2406_));
 sg13g2_and2_1 _6286_ (.A(_2396_),
    .B(_2402_),
    .X(_2407_));
 sg13g2_o21ai_1 _6287_ (.B1(_2349_),
    .Y(_2408_),
    .A1(\vgademo.a_sin[10] ),
    .A2(\vgademo.a_sin[11] ));
 sg13g2_nand2b_1 _6288_ (.Y(_2409_),
    .B(_2408_),
    .A_N(_2397_));
 sg13g2_a21oi_2 _6289_ (.B1(_2409_),
    .Y(_2410_),
    .A2(_2407_),
    .A1(_2398_));
 sg13g2_xnor2_1 _6290_ (.Y(_2411_),
    .A(_3167_),
    .B(net837));
 sg13g2_xnor2_1 _6291_ (.Y(_2412_),
    .A(_2410_),
    .B(_2411_));
 sg13g2_a21oi_1 _6292_ (.A1(net924),
    .A2(_2412_),
    .Y(_0285_),
    .B1(_2406_));
 sg13g2_o21ai_1 _6293_ (.B1(_2410_),
    .Y(_2413_),
    .A1(\vgademo.a_sin[12] ),
    .A2(net837));
 sg13g2_a21o_1 _6294_ (.A2(net837),
    .A1(\vgademo.a_sin[12] ),
    .B1(_2410_),
    .X(_2414_));
 sg13g2_nand3_1 _6295_ (.B(_2413_),
    .C(_2414_),
    .A(_0593_),
    .Y(_2415_));
 sg13g2_xnor2_1 _6296_ (.Y(_0286_),
    .A(net458),
    .B(_2415_));
 sg13g2_xor2_1 _6297_ (.B(net838),
    .A(\vgademo.a_sin[13] ),
    .X(_2416_));
 sg13g2_nor2_1 _6298_ (.A(_2415_),
    .B(_2416_),
    .Y(_2417_));
 sg13g2_xnor2_1 _6299_ (.Y(_0287_),
    .A(_3168_),
    .B(_2417_));
 sg13g2_and4_1 _6300_ (.A(\vgademo.h_count[10] ),
    .B(net1075),
    .C(_0578_),
    .D(_0579_),
    .X(_2418_));
 sg13g2_mux2_1 _6301_ (.A0(net317),
    .A1(_0498_),
    .S(net912),
    .X(_0288_));
 sg13g2_mux2_1 _6302_ (.A0(net378),
    .A1(_0512_),
    .S(net912),
    .X(_0289_));
 sg13g2_mux2_1 _6303_ (.A0(net347),
    .A1(_0526_),
    .S(net912),
    .X(_0290_));
 sg13g2_mux2_1 _6304_ (.A0(net509),
    .A1(_0542_),
    .S(net912),
    .X(_0291_));
 sg13g2_mux2_1 _6305_ (.A0(net430),
    .A1(_0556_),
    .S(net912),
    .X(_0292_));
 sg13g2_mux2_1 _6306_ (.A0(net360),
    .A1(_0562_),
    .S(net912),
    .X(_0293_));
 sg13g2_mux2_1 _6307_ (.A0(net463),
    .A1(_0560_),
    .S(net912),
    .X(_0294_));
 sg13g2_o21ai_1 _6308_ (.B1(net293),
    .Y(_2419_),
    .A1(_3148_),
    .A2(net927));
 sg13g2_nor2_2 _6309_ (.A(net293),
    .B(_3148_),
    .Y(_2420_));
 sg13g2_nor2_1 _6310_ (.A(net938),
    .B(net927),
    .Y(_2421_));
 sg13g2_nand2_2 _6311_ (.Y(_2422_),
    .A(net932),
    .B(_0583_));
 sg13g2_a22oi_1 _6312_ (.Y(_2423_),
    .B1(_2420_),
    .B2(net904),
    .A2(net908),
    .A1(\vgademo.a_cos[3] ));
 sg13g2_o21ai_1 _6313_ (.B1(_2423_),
    .Y(_0295_),
    .A1(net907),
    .A2(_2419_));
 sg13g2_nand2b_1 _6314_ (.Y(_2424_),
    .B(net907),
    .A_N(\vgademo.a_cos[4] ));
 sg13g2_xnor2_1 _6315_ (.Y(_2425_),
    .A(net433),
    .B(\vgademo.b_sin[8] ));
 sg13g2_nor2b_1 _6316_ (.A(_2420_),
    .B_N(_2425_),
    .Y(_2426_));
 sg13g2_xor2_1 _6317_ (.B(_2425_),
    .A(_2420_),
    .X(_2427_));
 sg13g2_o21ai_1 _6318_ (.B1(_2424_),
    .Y(_2428_),
    .A1(net433),
    .A2(_0583_));
 sg13g2_a21oi_1 _6319_ (.A1(net904),
    .A2(_2427_),
    .Y(_0296_),
    .B1(_2428_));
 sg13g2_a21oi_1 _6320_ (.A1(net594),
    .A2(_3150_),
    .Y(_2429_),
    .B1(_2426_));
 sg13g2_xnor2_1 _6321_ (.Y(_2430_),
    .A(net422),
    .B(\vgademo.b_sin[9] ));
 sg13g2_nor2b_1 _6322_ (.A(_2429_),
    .B_N(_2430_),
    .Y(_2431_));
 sg13g2_xor2_1 _6323_ (.B(_2430_),
    .A(_2429_),
    .X(_2432_));
 sg13g2_nand2b_1 _6324_ (.Y(_2433_),
    .B(net907),
    .A_N(\vgademo.a_cos[5] ));
 sg13g2_o21ai_1 _6325_ (.B1(_2433_),
    .Y(_2434_),
    .A1(net422),
    .A2(_0583_));
 sg13g2_a21oi_1 _6326_ (.A1(net904),
    .A2(_2432_),
    .Y(_0297_),
    .B1(net423));
 sg13g2_xnor2_1 _6327_ (.Y(_2435_),
    .A(\vgademo.b_cos[3] ),
    .B(\vgademo.b_sin[10] ));
 sg13g2_a21oi_1 _6328_ (.A1(\vgademo.b_cos[2] ),
    .A2(_3151_),
    .Y(_2436_),
    .B1(_2431_));
 sg13g2_nor2b_1 _6329_ (.A(_2436_),
    .B_N(_2435_),
    .Y(_2437_));
 sg13g2_xor2_1 _6330_ (.B(_2436_),
    .A(_2435_),
    .X(_2438_));
 sg13g2_nor2_1 _6331_ (.A(net325),
    .B(net929),
    .Y(_2439_));
 sg13g2_a221oi_1 _6332_ (.B2(_2438_),
    .C1(_2439_),
    .B1(net904),
    .A1(_3153_),
    .Y(_0298_),
    .A2(net908));
 sg13g2_xnor2_1 _6333_ (.Y(_2440_),
    .A(\vgademo.b_cos[4] ),
    .B(net965));
 sg13g2_a21oi_1 _6334_ (.A1(net325),
    .A2(_3152_),
    .Y(_2441_),
    .B1(_2437_));
 sg13g2_nor2b_1 _6335_ (.A(_2441_),
    .B_N(_2440_),
    .Y(_2442_));
 sg13g2_xor2_1 _6336_ (.B(_2441_),
    .A(_2440_),
    .X(_2443_));
 sg13g2_nor2_1 _6337_ (.A(net402),
    .B(net929),
    .Y(_2444_));
 sg13g2_a221oi_1 _6338_ (.B2(_2443_),
    .C1(_2444_),
    .B1(net904),
    .A1(_3155_),
    .Y(_0299_),
    .A2(net907));
 sg13g2_xnor2_1 _6339_ (.Y(_2445_),
    .A(net964),
    .B(\vgademo.b_cos[5] ));
 sg13g2_a21oi_1 _6340_ (.A1(net402),
    .A2(_3154_),
    .Y(_2446_),
    .B1(_2442_));
 sg13g2_xor2_1 _6341_ (.B(_2446_),
    .A(_2445_),
    .X(_2447_));
 sg13g2_a22oi_1 _6342_ (.Y(_2448_),
    .B1(net906),
    .B2(net555),
    .A2(net926),
    .A1(\vgademo.b_cos[5] ));
 sg13g2_o21ai_1 _6343_ (.B1(net556),
    .Y(_0300_),
    .A1(_2422_),
    .A2(_2447_));
 sg13g2_xor2_1 _6344_ (.B(net971),
    .A(net964),
    .X(_2449_));
 sg13g2_o21ai_1 _6345_ (.B1(_3154_),
    .Y(_2450_),
    .A1(\vgademo.b_cos[4] ),
    .A2(\vgademo.b_cos[5] ));
 sg13g2_nand2_1 _6346_ (.Y(_2451_),
    .A(_2442_),
    .B(_2445_));
 sg13g2_a21oi_1 _6347_ (.A1(_2450_),
    .A2(_2451_),
    .Y(_2452_),
    .B1(_2449_));
 sg13g2_nand3_1 _6348_ (.B(_2450_),
    .C(_2451_),
    .A(_2449_),
    .Y(_2453_));
 sg13g2_nand2_1 _6349_ (.Y(_2454_),
    .A(net903),
    .B(_2453_));
 sg13g2_a22oi_1 _6350_ (.Y(_2455_),
    .B1(net905),
    .B2(net511),
    .A2(net926),
    .A1(net971));
 sg13g2_o21ai_1 _6351_ (.B1(_2455_),
    .Y(_0301_),
    .A1(_2452_),
    .A2(_2454_));
 sg13g2_xor2_1 _6352_ (.B(\vgademo.b_cos[7] ),
    .A(net964),
    .X(_2456_));
 sg13g2_a21oi_1 _6353_ (.A1(_3154_),
    .A2(net971),
    .Y(_2457_),
    .B1(_2452_));
 sg13g2_xor2_1 _6354_ (.B(_2457_),
    .A(_2456_),
    .X(_2458_));
 sg13g2_nand2_1 _6355_ (.Y(_2459_),
    .A(net487),
    .B(net905));
 sg13g2_a22oi_1 _6356_ (.Y(_2460_),
    .B1(net903),
    .B2(_2458_),
    .A2(net926),
    .A1(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6357_ (.Y(_0302_),
    .A(_2459_),
    .B(_2460_));
 sg13g2_xor2_1 _6358_ (.B(\vgademo.b_cos[8] ),
    .A(net964),
    .X(_2461_));
 sg13g2_nor3_1 _6359_ (.A(_2449_),
    .B(_2451_),
    .C(_2456_),
    .Y(_2462_));
 sg13g2_o21ai_1 _6360_ (.B1(_3154_),
    .Y(_2463_),
    .A1(net971),
    .A2(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6361_ (.Y(_2464_),
    .A(_2450_),
    .B(_2463_));
 sg13g2_nor2_1 _6362_ (.A(_2462_),
    .B(_2464_),
    .Y(_2465_));
 sg13g2_nor2_1 _6363_ (.A(_2461_),
    .B(_2465_),
    .Y(_2466_));
 sg13g2_xor2_1 _6364_ (.B(_2465_),
    .A(_2461_),
    .X(_2467_));
 sg13g2_nand2_1 _6365_ (.Y(_2468_),
    .A(net466),
    .B(net905));
 sg13g2_a22oi_1 _6366_ (.Y(_2469_),
    .B1(net903),
    .B2(_2467_),
    .A2(net926),
    .A1(\vgademo.b_cos[8] ));
 sg13g2_nand2_1 _6367_ (.Y(_0303_),
    .A(_2468_),
    .B(_2469_));
 sg13g2_xnor2_1 _6368_ (.Y(_2470_),
    .A(net964),
    .B(\vgademo.b_cos[9] ));
 sg13g2_a21oi_1 _6369_ (.A1(_3154_),
    .A2(\vgademo.b_cos[8] ),
    .Y(_2471_),
    .B1(_2466_));
 sg13g2_xnor2_1 _6370_ (.Y(_2472_),
    .A(_2470_),
    .B(_2471_));
 sg13g2_nand2_1 _6371_ (.Y(_2473_),
    .A(net368),
    .B(net905));
 sg13g2_a22oi_1 _6372_ (.Y(_2474_),
    .B1(net903),
    .B2(_2472_),
    .A2(net926),
    .A1(\vgademo.b_cos[9] ));
 sg13g2_nand2_1 _6373_ (.Y(_0304_),
    .A(_2473_),
    .B(_2474_));
 sg13g2_a22oi_1 _6374_ (.Y(_2475_),
    .B1(_2466_),
    .B2(_2470_),
    .A2(\vgademo.b_cos[8] ),
    .A1(_3154_));
 sg13g2_o21ai_1 _6375_ (.B1(_2475_),
    .Y(_2476_),
    .A1(net964),
    .A2(_3158_));
 sg13g2_nor2_1 _6376_ (.A(net964),
    .B(_3159_),
    .Y(_2477_));
 sg13g2_xnor2_1 _6377_ (.Y(_2478_),
    .A(net965),
    .B(net970));
 sg13g2_xor2_1 _6378_ (.B(_2478_),
    .A(_2476_),
    .X(_2479_));
 sg13g2_a22oi_1 _6379_ (.Y(_2480_),
    .B1(net903),
    .B2(_2479_),
    .A2(net905),
    .A1(net585));
 sg13g2_o21ai_1 _6380_ (.B1(_2480_),
    .Y(_0305_),
    .A1(_3159_),
    .A2(net929));
 sg13g2_a21oi_2 _6381_ (.B1(_2477_),
    .Y(_2481_),
    .A2(_2478_),
    .A1(_2476_));
 sg13g2_xnor2_1 _6382_ (.Y(_2482_),
    .A(net965),
    .B(\vgademo.b_cos[11] ));
 sg13g2_xnor2_1 _6383_ (.Y(_2483_),
    .A(_2481_),
    .B(_2482_));
 sg13g2_a22oi_1 _6384_ (.Y(_2484_),
    .B1(net903),
    .B2(net851),
    .A2(net906),
    .A1(net472));
 sg13g2_o21ai_1 _6385_ (.B1(_2484_),
    .Y(_0306_),
    .A1(_3160_),
    .A2(net929));
 sg13g2_mux2_1 _6386_ (.A0(net336),
    .A1(_0226_),
    .S(_0649_),
    .X(_0307_));
 sg13g2_xor2_1 _6387_ (.B(\vgademo.plane_dx_div.d[17] ),
    .A(\vgademo.plane_dx_div.d[16] ),
    .X(_2485_));
 sg13g2_nor2_1 _6388_ (.A(net967),
    .B(_2485_),
    .Y(_2486_));
 sg13g2_a21oi_1 _6389_ (.A1(net967),
    .A2(_0070_),
    .Y(_2487_),
    .B1(_2486_));
 sg13g2_nand2_1 _6390_ (.Y(_2488_),
    .A(\vgademo.plane_dx_div.r[16] ),
    .B(_2487_));
 sg13g2_xnor2_1 _6391_ (.Y(_2489_),
    .A(\vgademo.plane_dx_div.r[16] ),
    .B(_2487_));
 sg13g2_a22oi_1 _6392_ (.Y(_2490_),
    .B1(_2489_),
    .B2(_0647_),
    .A2(_1063_),
    .A1(net945));
 sg13g2_mux2_1 _6393_ (.A0(_2490_),
    .A1(_1063_),
    .S(_1072_),
    .X(_2491_));
 sg13g2_o21ai_1 _6394_ (.B1(_2491_),
    .Y(_2492_),
    .A1(net428),
    .A2(_0649_));
 sg13g2_inv_1 _6395_ (.Y(_0308_),
    .A(_2492_));
 sg13g2_nor2_1 _6396_ (.A(net327),
    .B(_0649_),
    .Y(_2493_));
 sg13g2_o21ai_1 _6397_ (.B1(\vgademo.plane_dx_div.d[18] ),
    .Y(_2494_),
    .A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ));
 sg13g2_or3_2 _6398_ (.A(\vgademo.plane_dx_div.d[16] ),
    .B(\vgademo.plane_dx_div.d[17] ),
    .C(\vgademo.plane_dx_div.d[18] ),
    .X(_2495_));
 sg13g2_a21oi_1 _6399_ (.A1(_2494_),
    .A2(_2495_),
    .Y(_2496_),
    .B1(net966));
 sg13g2_a21oi_1 _6400_ (.A1(net966),
    .A2(_0073_),
    .Y(_2497_),
    .B1(_2496_));
 sg13g2_nand2_1 _6401_ (.Y(_2498_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2497_));
 sg13g2_xnor2_1 _6402_ (.Y(_2499_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2497_));
 sg13g2_xnor2_1 _6403_ (.Y(_2500_),
    .A(_2488_),
    .B(_2499_));
 sg13g2_nand2_1 _6404_ (.Y(_2501_),
    .A(_1063_),
    .B(_1071_));
 sg13g2_nand2b_1 _6405_ (.Y(_2502_),
    .B(_2501_),
    .A_N(_1085_));
 sg13g2_xor2_1 _6406_ (.B(_2501_),
    .A(_1085_),
    .X(_2503_));
 sg13g2_a221oi_1 _6407_ (.B2(net945),
    .C1(_2493_),
    .B1(_2503_),
    .A1(net916),
    .Y(_0309_),
    .A2(_2500_));
 sg13g2_xor2_1 _6408_ (.B(_2495_),
    .A(\vgademo.plane_dx_div.d[19] ),
    .X(_2504_));
 sg13g2_nor2_1 _6409_ (.A(net966),
    .B(_2504_),
    .Y(_2505_));
 sg13g2_a21oi_1 _6410_ (.A1(net966),
    .A2(_0076_),
    .Y(_2506_),
    .B1(_2505_));
 sg13g2_and2_1 _6411_ (.A(\vgademo.plane_dx_div.r[18] ),
    .B(_2506_),
    .X(_2507_));
 sg13g2_xor2_1 _6412_ (.B(_2506_),
    .A(net327),
    .X(_2508_));
 sg13g2_o21ai_1 _6413_ (.B1(_2498_),
    .Y(_2509_),
    .A1(_2488_),
    .A2(_2499_));
 sg13g2_and2_1 _6414_ (.A(_2508_),
    .B(_2509_),
    .X(_2510_));
 sg13g2_xnor2_1 _6415_ (.Y(_2511_),
    .A(_2508_),
    .B(_2509_));
 sg13g2_nor2_1 _6416_ (.A(net334),
    .B(_0649_),
    .Y(_2512_));
 sg13g2_nand2b_1 _6417_ (.Y(_2513_),
    .B(_1100_),
    .A_N(_2502_));
 sg13g2_xor2_1 _6418_ (.B(_2502_),
    .A(_1100_),
    .X(_2514_));
 sg13g2_a221oi_1 _6419_ (.B2(net945),
    .C1(_2512_),
    .B1(_2514_),
    .A1(net916),
    .Y(_0310_),
    .A2(_2511_));
 sg13g2_o21ai_1 _6420_ (.B1(\vgademo.plane_dx_div.d[20] ),
    .Y(_2515_),
    .A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2495_));
 sg13g2_or3_2 _6421_ (.A(\vgademo.plane_dx_div.d[19] ),
    .B(\vgademo.plane_dx_div.d[20] ),
    .C(_2495_),
    .X(_2516_));
 sg13g2_a21oi_1 _6422_ (.A1(_2515_),
    .A2(_2516_),
    .Y(_2517_),
    .B1(net967));
 sg13g2_a21oi_1 _6423_ (.A1(net967),
    .A2(_0079_),
    .Y(_2518_),
    .B1(_2517_));
 sg13g2_nand2_1 _6424_ (.Y(_2519_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .B(_2518_));
 sg13g2_xor2_1 _6425_ (.B(_2518_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .X(_2520_));
 sg13g2_o21ai_1 _6426_ (.B1(_2520_),
    .Y(_2521_),
    .A1(_2507_),
    .A2(_2510_));
 sg13g2_or3_1 _6427_ (.A(_2507_),
    .B(_2510_),
    .C(_2520_),
    .X(_2522_));
 sg13g2_nand2_1 _6428_ (.Y(_2523_),
    .A(_2521_),
    .B(_2522_));
 sg13g2_nor2_1 _6429_ (.A(net312),
    .B(_0649_),
    .Y(_2524_));
 sg13g2_nor2_1 _6430_ (.A(_1118_),
    .B(_2513_),
    .Y(_2525_));
 sg13g2_xnor2_1 _6431_ (.Y(_2526_),
    .A(_1118_),
    .B(_2513_));
 sg13g2_a221oi_1 _6432_ (.B2(net946),
    .C1(_2524_),
    .B1(_2526_),
    .A1(net916),
    .Y(_0311_),
    .A2(_2523_));
 sg13g2_nand2_1 _6433_ (.Y(_2527_),
    .A(_1135_),
    .B(_2525_));
 sg13g2_xor2_1 _6434_ (.B(_2525_),
    .A(_1135_),
    .X(_2528_));
 sg13g2_xor2_1 _6435_ (.B(_2516_),
    .A(\vgademo.plane_dx_div.d[21] ),
    .X(_2529_));
 sg13g2_nor2_1 _6436_ (.A(net966),
    .B(_2529_),
    .Y(_2530_));
 sg13g2_a21oi_1 _6437_ (.A1(net966),
    .A2(_0081_),
    .Y(_2531_),
    .B1(_2530_));
 sg13g2_xnor2_1 _6438_ (.Y(_2532_),
    .A(\vgademo.plane_dx_div.r[20] ),
    .B(_2531_));
 sg13g2_a21oi_1 _6439_ (.A1(_2519_),
    .A2(_2521_),
    .Y(_2533_),
    .B1(_2532_));
 sg13g2_and3_1 _6440_ (.X(_2534_),
    .A(_2519_),
    .B(_2521_),
    .C(_2532_));
 sg13g2_o21ai_1 _6441_ (.B1(net916),
    .Y(_2535_),
    .A1(_2533_),
    .A2(_2534_));
 sg13g2_o21ai_1 _6442_ (.B1(_2535_),
    .Y(_2536_),
    .A1(net944),
    .A2(_2528_));
 sg13g2_a21oi_1 _6443_ (.A1(_3134_),
    .A2(_0648_),
    .Y(_0312_),
    .B1(_2536_));
 sg13g2_a21oi_1 _6444_ (.A1(\vgademo.plane_dx_div.r[20] ),
    .A2(_2531_),
    .Y(_2537_),
    .B1(_2533_));
 sg13g2_nand2b_1 _6445_ (.Y(_2538_),
    .B(net966),
    .A_N(_0013_));
 sg13g2_nor3_2 _6446_ (.A(\vgademo.plane_dx_div.d[21] ),
    .B(\vgademo.plane_dx_div.d[22] ),
    .C(_2516_),
    .Y(_2539_));
 sg13g2_o21ai_1 _6447_ (.B1(\vgademo.plane_dx_div.d[22] ),
    .Y(_2540_),
    .A1(\vgademo.plane_dx_div.d[21] ),
    .A2(_2516_));
 sg13g2_nor2b_1 _6448_ (.A(net966),
    .B_N(_2540_),
    .Y(_2541_));
 sg13g2_nand2b_1 _6449_ (.Y(_2542_),
    .B(_2541_),
    .A_N(_2539_));
 sg13g2_a21oi_1 _6450_ (.A1(_2538_),
    .A2(_2542_),
    .Y(_2543_),
    .B1(_3134_));
 sg13g2_and3_1 _6451_ (.X(_2544_),
    .A(_3134_),
    .B(_2538_),
    .C(_2542_));
 sg13g2_nor2_1 _6452_ (.A(_2543_),
    .B(_2544_),
    .Y(_2545_));
 sg13g2_xor2_1 _6453_ (.B(_2545_),
    .A(_2537_),
    .X(_2546_));
 sg13g2_nor2_1 _6454_ (.A(net321),
    .B(_0649_),
    .Y(_2547_));
 sg13g2_nand2b_1 _6455_ (.Y(_2548_),
    .B(_1153_),
    .A_N(_2527_));
 sg13g2_xor2_1 _6456_ (.B(_2527_),
    .A(_1153_),
    .X(_2549_));
 sg13g2_a221oi_1 _6457_ (.B2(net947),
    .C1(_2547_),
    .B1(_2549_),
    .A1(net916),
    .Y(_0313_),
    .A2(_2546_));
 sg13g2_nand2b_1 _6458_ (.Y(_2550_),
    .B(\vgademo.plane_dx_div.d[23] ),
    .A_N(_2539_));
 sg13g2_nand2b_1 _6459_ (.Y(_2551_),
    .B(_2539_),
    .A_N(\vgademo.plane_dx_div.d[23] ));
 sg13g2_a21oi_1 _6460_ (.A1(_2550_),
    .A2(_2551_),
    .Y(_2552_),
    .B1(net969));
 sg13g2_a21oi_1 _6461_ (.A1(net969),
    .A2(_0017_),
    .Y(_2553_),
    .B1(_2552_));
 sg13g2_and2_1 _6462_ (.A(\vgademo.plane_dx_div.r[22] ),
    .B(_2553_),
    .X(_2554_));
 sg13g2_xor2_1 _6463_ (.B(_2553_),
    .A(\vgademo.plane_dx_div.r[22] ),
    .X(_2555_));
 sg13g2_nor2b_1 _6464_ (.A(_2543_),
    .B_N(_2537_),
    .Y(_2556_));
 sg13g2_nor2_1 _6465_ (.A(_2544_),
    .B(_2556_),
    .Y(_2557_));
 sg13g2_and2_1 _6466_ (.A(_2555_),
    .B(_2557_),
    .X(_2558_));
 sg13g2_xor2_1 _6467_ (.B(_2557_),
    .A(_2555_),
    .X(_2559_));
 sg13g2_a21oi_1 _6468_ (.A1(_0646_),
    .A2(_2559_),
    .Y(_2560_),
    .B1(_0648_));
 sg13g2_nand2_1 _6469_ (.Y(_2561_),
    .A(_1169_),
    .B(_2548_));
 sg13g2_or2_1 _6470_ (.X(_2562_),
    .B(_2548_),
    .A(_1169_));
 sg13g2_nand3_1 _6471_ (.B(_2561_),
    .C(_2562_),
    .A(net947),
    .Y(_2563_));
 sg13g2_a22oi_1 _6472_ (.Y(_0314_),
    .B1(_2560_),
    .B2(_2563_),
    .A2(net914),
    .A1(_3137_));
 sg13g2_nand2_1 _6473_ (.Y(_2564_),
    .A(\vgademo.plane_dx_div.d[24] ),
    .B(_2551_));
 sg13g2_nor2_1 _6474_ (.A(\vgademo.plane_dx_div.d[24] ),
    .B(_2551_),
    .Y(_2565_));
 sg13g2_nor2_1 _6475_ (.A(net968),
    .B(_2565_),
    .Y(_2566_));
 sg13g2_a22oi_1 _6476_ (.Y(_2567_),
    .B1(_2564_),
    .B2(_2566_),
    .A2(_3136_),
    .A1(net968));
 sg13g2_xnor2_1 _6477_ (.Y(_2568_),
    .A(\vgademo.plane_dx_div.r[23] ),
    .B(_2567_));
 sg13g2_or3_1 _6478_ (.A(_2554_),
    .B(_2558_),
    .C(_2568_),
    .X(_2569_));
 sg13g2_o21ai_1 _6479_ (.B1(_2568_),
    .Y(_2570_),
    .A1(_2554_),
    .A2(_2558_));
 sg13g2_nand3_1 _6480_ (.B(_2569_),
    .C(_2570_),
    .A(net944),
    .Y(_2571_));
 sg13g2_nand2_1 _6481_ (.Y(_2572_),
    .A(_1179_),
    .B(_2562_));
 sg13g2_a21o_1 _6482_ (.A2(_2562_),
    .A1(net947),
    .B1(_1180_),
    .X(_2573_));
 sg13g2_a21oi_1 _6483_ (.A1(_2572_),
    .A2(_2573_),
    .Y(_2574_),
    .B1(net914));
 sg13g2_a22oi_1 _6484_ (.Y(_0315_),
    .B1(_2571_),
    .B2(_2574_),
    .A2(net914),
    .A1(_3138_));
 sg13g2_nand2_1 _6485_ (.Y(_2575_),
    .A(net968),
    .B(net914));
 sg13g2_o21ai_1 _6486_ (.B1(_2570_),
    .Y(_2576_),
    .A1(_3137_),
    .A2(_2567_));
 sg13g2_xnor2_1 _6487_ (.Y(_2577_),
    .A(\vgademo.plane_dx_div.r[24] ),
    .B(_2566_));
 sg13g2_xnor2_1 _6488_ (.Y(_2578_),
    .A(_2576_),
    .B(_2577_));
 sg13g2_a21oi_1 _6489_ (.A1(_0646_),
    .A2(_2578_),
    .Y(_2579_),
    .B1(_2573_));
 sg13g2_o21ai_1 _6490_ (.B1(_2575_),
    .Y(_0316_),
    .A1(net914),
    .A2(_2579_));
 sg13g2_or2_1 _6491_ (.X(_2580_),
    .B(_2188_),
    .A(_2161_));
 sg13g2_o21ai_1 _6492_ (.B1(_1861_),
    .Y(_2581_),
    .A1(_1810_),
    .A2(_1819_));
 sg13g2_mux2_1 _6493_ (.A0(_2581_),
    .A1(_2580_),
    .S(net834),
    .X(_2582_));
 sg13g2_a21o_1 _6494_ (.A2(_2582_),
    .A1(net872),
    .B1(_2192_),
    .X(_2583_));
 sg13g2_a21oi_2 _6495_ (.B1(_2182_),
    .Y(_2584_),
    .A2(_2583_),
    .A1(net835));
 sg13g2_nor2b_1 _6496_ (.A(_2584_),
    .B_N(net953),
    .Y(_2585_));
 sg13g2_a21o_2 _6497_ (.A2(_1858_),
    .A1(_1815_),
    .B1(_2162_),
    .X(_2586_));
 sg13g2_inv_1 _6498_ (.Y(_2587_),
    .A(_2586_));
 sg13g2_a21oi_1 _6499_ (.A1(net834),
    .A2(_2586_),
    .Y(_2588_),
    .B1(net866));
 sg13g2_a21o_1 _6500_ (.A2(_2166_),
    .A1(net866),
    .B1(_1756_),
    .X(_2589_));
 sg13g2_or2_1 _6501_ (.X(_2590_),
    .B(_2178_),
    .A(_2156_));
 sg13g2_nor2_1 _6502_ (.A(net836),
    .B(_2181_),
    .Y(_2591_));
 sg13g2_a21oi_1 _6503_ (.A1(_2590_),
    .A2(_2591_),
    .Y(_2592_),
    .B1(net879));
 sg13g2_o21ai_1 _6504_ (.B1(_2592_),
    .Y(_2593_),
    .A1(_2588_),
    .A2(_2589_));
 sg13g2_xnor2_1 _6505_ (.Y(_2594_),
    .A(net953),
    .B(_2584_));
 sg13g2_a21oi_1 _6506_ (.A1(_2593_),
    .A2(_2594_),
    .Y(_2595_),
    .B1(_2585_));
 sg13g2_nand3_1 _6507_ (.B(net832),
    .C(_2581_),
    .A(net872),
    .Y(_2596_));
 sg13g2_nor2_1 _6508_ (.A(_1756_),
    .B(_2142_),
    .Y(_2597_));
 sg13g2_and2_1 _6509_ (.A(_2152_),
    .B(_2590_),
    .X(_2598_));
 sg13g2_a221oi_1 _6510_ (.B2(_1756_),
    .C1(net879),
    .B1(_2598_),
    .A1(_2596_),
    .Y(_2599_),
    .A2(_2597_));
 sg13g2_a21oi_1 _6511_ (.A1(_1274_),
    .A2(_1297_),
    .Y(_2600_),
    .B1(_2599_));
 sg13g2_inv_1 _6512_ (.Y(_2601_),
    .A(_2600_));
 sg13g2_a21oi_1 _6513_ (.A1(_2173_),
    .A2(_2593_),
    .Y(_2602_),
    .B1(_2601_));
 sg13g2_xnor2_1 _6514_ (.Y(_2603_),
    .A(_2172_),
    .B(_2593_));
 sg13g2_xnor2_1 _6515_ (.Y(_2604_),
    .A(_2601_),
    .B(_2603_));
 sg13g2_or2_1 _6516_ (.X(_2605_),
    .B(_2604_),
    .A(_2595_));
 sg13g2_nor2_1 _6517_ (.A(_2187_),
    .B(_2219_),
    .Y(_2606_));
 sg13g2_mux2_1 _6518_ (.A0(_2587_),
    .A1(_2606_),
    .S(net834),
    .X(_2607_));
 sg13g2_a21oi_1 _6519_ (.A1(net872),
    .A2(_2607_),
    .Y(_2608_),
    .B1(_2236_));
 sg13g2_a21o_1 _6520_ (.A2(_2607_),
    .A1(net871),
    .B1(_2236_),
    .X(_2609_));
 sg13g2_nor2_1 _6521_ (.A(_2153_),
    .B(_2179_),
    .Y(_2610_));
 sg13g2_nor4_1 _6522_ (.A(net836),
    .B(_2153_),
    .C(_2156_),
    .D(_2178_),
    .Y(_2611_));
 sg13g2_a21oi_1 _6523_ (.A1(_2155_),
    .A2(_2157_),
    .Y(_2612_),
    .B1(_2611_));
 sg13g2_a21o_1 _6524_ (.A2(_2157_),
    .A1(_2155_),
    .B1(_2611_),
    .X(_2613_));
 sg13g2_nor2_1 _6525_ (.A(_2608_),
    .B(_2613_),
    .Y(_2614_));
 sg13g2_nand2b_1 _6526_ (.Y(_2615_),
    .B(_2580_),
    .A_N(net832));
 sg13g2_nand2_1 _6527_ (.Y(_2616_),
    .A(_2211_),
    .B(_2218_));
 sg13g2_a21oi_1 _6528_ (.A1(net832),
    .A2(_2616_),
    .Y(_2617_),
    .B1(_1322_));
 sg13g2_a21oi_2 _6529_ (.B1(_2205_),
    .Y(_2618_),
    .A2(_2617_),
    .A1(_2615_));
 sg13g2_nor2_2 _6530_ (.A(net879),
    .B(_2618_),
    .Y(_2619_));
 sg13g2_nand2_1 _6531_ (.Y(_2620_),
    .A(_2243_),
    .B(_2599_));
 sg13g2_a22oi_1 _6532_ (.Y(_2621_),
    .B1(_2619_),
    .B2(_2620_),
    .A2(_2600_),
    .A1(_2244_));
 sg13g2_nand2b_1 _6533_ (.Y(_2622_),
    .B(_2621_),
    .A_N(_2614_));
 sg13g2_or2_1 _6534_ (.X(_2623_),
    .B(_2606_),
    .A(net832));
 sg13g2_nand2_1 _6535_ (.Y(_2624_),
    .A(_2210_),
    .B(_2221_));
 sg13g2_a21oi_1 _6536_ (.A1(net832),
    .A2(_2624_),
    .Y(_2625_),
    .B1(net866));
 sg13g2_a21oi_2 _6537_ (.B1(_2203_),
    .Y(_2626_),
    .A2(_2625_),
    .A1(_2623_));
 sg13g2_nor2_1 _6538_ (.A(net879),
    .B(_2626_),
    .Y(_2627_));
 sg13g2_o21ai_1 _6539_ (.B1(net951),
    .Y(_2628_),
    .A1(net878),
    .A2(_2626_));
 sg13g2_nor3_1 _6540_ (.A(net878),
    .B(net951),
    .C(_2626_),
    .Y(_2629_));
 sg13g2_xor2_1 _6541_ (.B(_2627_),
    .A(net951),
    .X(_2630_));
 sg13g2_xnor2_1 _6542_ (.Y(_2631_),
    .A(_2619_),
    .B(_2630_));
 sg13g2_o21ai_1 _6543_ (.B1(_2628_),
    .Y(_2632_),
    .A1(_2619_),
    .A2(_2629_));
 sg13g2_a21oi_1 _6544_ (.A1(_2609_),
    .A2(_2612_),
    .Y(_2633_),
    .B1(_2251_));
 sg13g2_nor3_1 _6545_ (.A(_2252_),
    .B(_2608_),
    .C(_2613_),
    .Y(_2634_));
 sg13g2_or3_1 _6546_ (.A(_2584_),
    .B(_2633_),
    .C(_2634_),
    .X(_2635_));
 sg13g2_o21ai_1 _6547_ (.B1(_2584_),
    .Y(_2636_),
    .A1(_2633_),
    .A2(_2634_));
 sg13g2_a21o_1 _6548_ (.A2(_2636_),
    .A1(_2635_),
    .B1(_2632_),
    .X(_2637_));
 sg13g2_nor2b_1 _6549_ (.A(_2621_),
    .B_N(_2614_),
    .Y(_2638_));
 sg13g2_o21ai_1 _6550_ (.B1(_2622_),
    .Y(_2639_),
    .A1(_2631_),
    .A2(_2638_));
 sg13g2_nand3_1 _6551_ (.B(_2635_),
    .C(_2636_),
    .A(_2632_),
    .Y(_2640_));
 sg13g2_nor2b_1 _6552_ (.A(_2633_),
    .B_N(_2635_),
    .Y(_2641_));
 sg13g2_xnor2_1 _6553_ (.Y(_2642_),
    .A(_2593_),
    .B(_2594_));
 sg13g2_o21ai_1 _6554_ (.B1(_2640_),
    .Y(_2643_),
    .A1(_2641_),
    .A2(_2642_));
 sg13g2_a21oi_1 _6555_ (.A1(_2637_),
    .A2(_2639_),
    .Y(_2644_),
    .B1(_2643_));
 sg13g2_a22oi_1 _6556_ (.Y(_2645_),
    .B1(_2641_),
    .B2(_2642_),
    .A2(_2604_),
    .A1(_2595_));
 sg13g2_inv_1 _6557_ (.Y(_2646_),
    .A(_2645_));
 sg13g2_o21ai_1 _6558_ (.B1(_2605_),
    .Y(_2647_),
    .A1(_2644_),
    .A2(_2646_));
 sg13g2_o21ai_1 _6559_ (.B1(_2601_),
    .Y(_2648_),
    .A1(_2173_),
    .A2(_2593_));
 sg13g2_nor2b_1 _6560_ (.A(_2602_),
    .B_N(_2648_),
    .Y(_2649_));
 sg13g2_nor2_1 _6561_ (.A(_2647_),
    .B(_2649_),
    .Y(_2650_));
 sg13g2_nand2_1 _6562_ (.Y(_2651_),
    .A(_2647_),
    .B(_2649_));
 sg13g2_a21oi_1 _6563_ (.A1(_2647_),
    .A2(_2649_),
    .Y(_2652_),
    .B1(_2274_));
 sg13g2_nor2b_1 _6564_ (.A(_2650_),
    .B_N(_2652_),
    .Y(_0317_));
 sg13g2_a21oi_1 _6565_ (.A1(_2648_),
    .A2(_2651_),
    .Y(_0318_),
    .B1(_2274_));
 sg13g2_nand2_1 _6566_ (.Y(_2653_),
    .A(\vgademo.b_sin[0] ),
    .B(_2458_));
 sg13g2_xnor2_1 _6567_ (.Y(_2654_),
    .A(net379),
    .B(_2458_));
 sg13g2_a22oi_1 _6568_ (.Y(_2655_),
    .B1(net905),
    .B2(\vgademo.a_sin[3] ),
    .A2(net926),
    .A1(net379));
 sg13g2_o21ai_1 _6569_ (.B1(net380),
    .Y(_0319_),
    .A1(_2422_),
    .A2(_2654_));
 sg13g2_nand2_1 _6570_ (.Y(_2656_),
    .A(\vgademo.b_sin[1] ),
    .B(_2467_));
 sg13g2_xnor2_1 _6571_ (.Y(_2657_),
    .A(\vgademo.b_sin[1] ),
    .B(_2467_));
 sg13g2_xnor2_1 _6572_ (.Y(_2658_),
    .A(_2653_),
    .B(_2657_));
 sg13g2_a22oi_1 _6573_ (.Y(_2659_),
    .B1(net905),
    .B2(net346),
    .A2(net926),
    .A1(net356));
 sg13g2_o21ai_1 _6574_ (.B1(_2659_),
    .Y(_0320_),
    .A1(_2422_),
    .A2(_2658_));
 sg13g2_o21ai_1 _6575_ (.B1(_2656_),
    .Y(_2660_),
    .A1(_2653_),
    .A2(_2657_));
 sg13g2_nand2_1 _6576_ (.Y(_2661_),
    .A(\vgademo.b_sin[2] ),
    .B(_2472_));
 sg13g2_xnor2_1 _6577_ (.Y(_2662_),
    .A(\vgademo.b_sin[2] ),
    .B(_2472_));
 sg13g2_nand2b_1 _6578_ (.Y(_2663_),
    .B(_2660_),
    .A_N(_2662_));
 sg13g2_xor2_1 _6579_ (.B(_2662_),
    .A(_2660_),
    .X(_2664_));
 sg13g2_a22oi_1 _6580_ (.Y(_2665_),
    .B1(net906),
    .B2(net341),
    .A2(net926),
    .A1(\vgademo.b_sin[2] ));
 sg13g2_o21ai_1 _6581_ (.B1(net342),
    .Y(_0321_),
    .A1(_2422_),
    .A2(_2664_));
 sg13g2_nand2_1 _6582_ (.Y(_2666_),
    .A(net414),
    .B(_2479_));
 sg13g2_xnor2_1 _6583_ (.Y(_2667_),
    .A(\vgademo.b_sin[3] ),
    .B(_2479_));
 sg13g2_nand3_1 _6584_ (.B(_2663_),
    .C(_2667_),
    .A(_2661_),
    .Y(_2668_));
 sg13g2_a21o_1 _6585_ (.A2(_2663_),
    .A1(_2661_),
    .B1(_2667_),
    .X(_2669_));
 sg13g2_nand3_1 _6586_ (.B(_2668_),
    .C(_2669_),
    .A(net903),
    .Y(_2670_));
 sg13g2_a22oi_1 _6587_ (.Y(_2671_),
    .B1(net906),
    .B2(\vgademo.a_sin[6] ),
    .A2(net928),
    .A1(net414));
 sg13g2_nand2_1 _6588_ (.Y(_0322_),
    .A(_2670_),
    .B(net415));
 sg13g2_xnor2_1 _6589_ (.Y(_2672_),
    .A(\vgademo.b_sin[4] ),
    .B(net851));
 sg13g2_nand3_1 _6590_ (.B(_2669_),
    .C(_2672_),
    .A(_2666_),
    .Y(_2673_));
 sg13g2_a21oi_2 _6591_ (.B1(_2672_),
    .Y(_2674_),
    .A2(_2669_),
    .A1(_2666_));
 sg13g2_inv_1 _6592_ (.Y(_2675_),
    .A(_2674_));
 sg13g2_nand2_1 _6593_ (.Y(_2676_),
    .A(net903),
    .B(_2673_));
 sg13g2_a22oi_1 _6594_ (.Y(_2677_),
    .B1(net907),
    .B2(\vgademo.a_sin[7] ),
    .A2(net928),
    .A1(net456));
 sg13g2_o21ai_1 _6595_ (.B1(net457),
    .Y(_0323_),
    .A1(_2674_),
    .A2(_2676_));
 sg13g2_nand2_1 _6596_ (.Y(_2678_),
    .A(net260),
    .B(net927));
 sg13g2_xnor2_1 _6597_ (.Y(_2679_),
    .A(\vgademo.b_sin[5] ),
    .B(net850));
 sg13g2_a21o_1 _6598_ (.A2(net850),
    .A1(\vgademo.b_sin[4] ),
    .B1(_2674_),
    .X(_2680_));
 sg13g2_o21ai_1 _6599_ (.B1(net932),
    .Y(_2681_),
    .A1(_2679_),
    .A2(_2680_));
 sg13g2_a21oi_1 _6600_ (.A1(_2679_),
    .A2(_2680_),
    .Y(_2682_),
    .B1(_2681_));
 sg13g2_o21ai_1 _6601_ (.B1(net929),
    .Y(_2683_),
    .A1(\vgademo.a_sin[8] ),
    .A2(net932));
 sg13g2_o21ai_1 _6602_ (.B1(_2678_),
    .Y(_0324_),
    .A1(_2682_),
    .A2(_2683_));
 sg13g2_xnor2_1 _6603_ (.Y(_2684_),
    .A(\vgademo.b_sin[6] ),
    .B(net849));
 sg13g2_o21ai_1 _6604_ (.B1(net849),
    .Y(_2685_),
    .A1(\vgademo.b_sin[4] ),
    .A2(\vgademo.b_sin[5] ));
 sg13g2_nor2_1 _6605_ (.A(_2675_),
    .B(_2679_),
    .Y(_2686_));
 sg13g2_nor2b_1 _6606_ (.A(_2686_),
    .B_N(_2685_),
    .Y(_2687_));
 sg13g2_nor2_1 _6607_ (.A(_2684_),
    .B(_2687_),
    .Y(_2688_));
 sg13g2_a21o_1 _6608_ (.A2(_2687_),
    .A1(_2684_),
    .B1(_2422_),
    .X(_2689_));
 sg13g2_a22oi_1 _6609_ (.Y(_2690_),
    .B1(net907),
    .B2(\vgademo.a_sin[9] ),
    .A2(net927),
    .A1(net440));
 sg13g2_o21ai_1 _6610_ (.B1(net441),
    .Y(_0325_),
    .A1(_2688_),
    .A2(_2689_));
 sg13g2_nand2_1 _6611_ (.Y(_2691_),
    .A(net267),
    .B(net927));
 sg13g2_xnor2_1 _6612_ (.Y(_2692_),
    .A(_3148_),
    .B(net849));
 sg13g2_a21oi_1 _6613_ (.A1(\vgademo.b_sin[6] ),
    .A2(net849),
    .Y(_2693_),
    .B1(_2688_));
 sg13g2_o21ai_1 _6614_ (.B1(net932),
    .Y(_2694_),
    .A1(_2692_),
    .A2(_2693_));
 sg13g2_a21oi_1 _6615_ (.A1(_2692_),
    .A2(_2693_),
    .Y(_2695_),
    .B1(_2694_));
 sg13g2_o21ai_1 _6616_ (.B1(net929),
    .Y(_2696_),
    .A1(\vgademo.a_sin[10] ),
    .A2(net932));
 sg13g2_o21ai_1 _6617_ (.B1(_2691_),
    .Y(_0326_),
    .A1(_2695_),
    .A2(_2696_));
 sg13g2_nand2_1 _6618_ (.Y(_2697_),
    .A(\vgademo.b_sin[8] ),
    .B(net849));
 sg13g2_xnor2_1 _6619_ (.Y(_2698_),
    .A(\vgademo.b_sin[8] ),
    .B(net849));
 sg13g2_nor2b_1 _6620_ (.A(_2684_),
    .B_N(_2692_),
    .Y(_2699_));
 sg13g2_o21ai_1 _6621_ (.B1(net849),
    .Y(_2700_),
    .A1(\vgademo.b_sin[7] ),
    .A2(\vgademo.b_sin[6] ));
 sg13g2_nand2_1 _6622_ (.Y(_2701_),
    .A(_2685_),
    .B(_2700_));
 sg13g2_a21oi_1 _6623_ (.A1(_2686_),
    .A2(_2699_),
    .Y(_2702_),
    .B1(_2701_));
 sg13g2_or2_1 _6624_ (.X(_2703_),
    .B(_2702_),
    .A(_2698_));
 sg13g2_a21oi_1 _6625_ (.A1(_2698_),
    .A2(_2702_),
    .Y(_2704_),
    .B1(_2422_));
 sg13g2_nand2_1 _6626_ (.Y(_2705_),
    .A(_2703_),
    .B(_2704_));
 sg13g2_a22oi_1 _6627_ (.Y(_2706_),
    .B1(net907),
    .B2(\vgademo.a_sin[11] ),
    .A2(net927),
    .A1(net481));
 sg13g2_nand2_1 _6628_ (.Y(_0327_),
    .A(_2705_),
    .B(net482));
 sg13g2_nand2_1 _6629_ (.Y(_2707_),
    .A(net382),
    .B(net927));
 sg13g2_o21ai_1 _6630_ (.B1(net929),
    .Y(_2708_),
    .A1(\vgademo.a_sin[12] ),
    .A2(net932));
 sg13g2_nand2_1 _6631_ (.Y(_2709_),
    .A(_2697_),
    .B(_2703_));
 sg13g2_xnor2_1 _6632_ (.Y(_2710_),
    .A(\vgademo.b_sin[9] ),
    .B(net849));
 sg13g2_o21ai_1 _6633_ (.B1(net932),
    .Y(_2711_),
    .A1(_2709_),
    .A2(_2710_));
 sg13g2_a21oi_1 _6634_ (.A1(_2709_),
    .A2(_2710_),
    .Y(_2712_),
    .B1(_2711_));
 sg13g2_o21ai_1 _6635_ (.B1(_2707_),
    .Y(_0328_),
    .A1(_2708_),
    .A2(_2712_));
 sg13g2_nand2_1 _6636_ (.Y(_2713_),
    .A(\vgademo.b_sin[10] ),
    .B(net851));
 sg13g2_xnor2_1 _6637_ (.Y(_2714_),
    .A(\vgademo.b_sin[10] ),
    .B(net850));
 sg13g2_a21o_1 _6638_ (.A2(net850),
    .A1(\vgademo.b_sin[9] ),
    .B1(_2709_),
    .X(_2715_));
 sg13g2_o21ai_1 _6639_ (.B1(_2715_),
    .Y(_2716_),
    .A1(\vgademo.b_sin[9] ),
    .A2(net850));
 sg13g2_or2_1 _6640_ (.X(_2717_),
    .B(_2716_),
    .A(_2714_));
 sg13g2_a21oi_1 _6641_ (.A1(_2714_),
    .A2(_2716_),
    .Y(_2718_),
    .B1(_2422_));
 sg13g2_nand2_1 _6642_ (.Y(_2719_),
    .A(_2717_),
    .B(_2718_));
 sg13g2_a22oi_1 _6643_ (.Y(_2720_),
    .B1(net907),
    .B2(net458),
    .A2(net927),
    .A1(net490));
 sg13g2_nand2_1 _6644_ (.Y(_0329_),
    .A(_2719_),
    .B(_2720_));
 sg13g2_nand2_1 _6645_ (.Y(_2721_),
    .A(net965),
    .B(net928));
 sg13g2_nand2_1 _6646_ (.Y(_2722_),
    .A(_2713_),
    .B(_2717_));
 sg13g2_xnor2_1 _6647_ (.Y(_2723_),
    .A(\vgademo.b_cos[11] ),
    .B(_2481_));
 sg13g2_o21ai_1 _6648_ (.B1(net934),
    .Y(_2724_),
    .A1(_2722_),
    .A2(_2723_));
 sg13g2_a21oi_1 _6649_ (.A1(_2722_),
    .A2(_2723_),
    .Y(_2725_),
    .B1(_2724_));
 sg13g2_o21ai_1 _6650_ (.B1(net929),
    .Y(_2726_),
    .A1(net972),
    .A2(net934));
 sg13g2_o21ai_1 _6651_ (.B1(_2721_),
    .Y(_0330_),
    .A1(_2725_),
    .A2(_2726_));
 sg13g2_o21ai_1 _6652_ (.B1(net1078),
    .Y(_2727_),
    .A1(net941),
    .A2(_2270_));
 sg13g2_inv_1 _6653_ (.Y(_2728_),
    .A(net900));
 sg13g2_nand2_1 _6654_ (.Y(_2729_),
    .A(net211),
    .B(\vgademo.plane_du[0] ));
 sg13g2_nand2_1 _6655_ (.Y(_2730_),
    .A(net283),
    .B(net310));
 sg13g2_xor2_1 _6656_ (.B(\vgademo.plane_du[1] ),
    .A(\vgademo.plane_u[1] ),
    .X(_2731_));
 sg13g2_nand2b_1 _6657_ (.Y(_2732_),
    .B(_2731_),
    .A_N(_2729_));
 sg13g2_xor2_1 _6658_ (.B(_2731_),
    .A(_2729_),
    .X(_2733_));
 sg13g2_nor2_1 _6659_ (.A(net938),
    .B(_2733_),
    .Y(_2734_));
 sg13g2_a21oi_1 _6660_ (.A1(\vgademo.plane_dx[0] ),
    .A2(net937),
    .Y(_2735_),
    .B1(_2734_));
 sg13g2_nand2_1 _6661_ (.Y(_2736_),
    .A(net283),
    .B(net900));
 sg13g2_o21ai_1 _6662_ (.B1(_2736_),
    .Y(_0331_),
    .A1(net900),
    .A2(_2735_));
 sg13g2_nand2_1 _6663_ (.Y(_2737_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_xnor2_1 _6664_ (.Y(_2738_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_nand3_1 _6665_ (.B(_2732_),
    .C(_2738_),
    .A(_2730_),
    .Y(_2739_));
 sg13g2_a21o_1 _6666_ (.A2(_2732_),
    .A1(_2730_),
    .B1(_2738_),
    .X(_2740_));
 sg13g2_nand3_1 _6667_ (.B(_2739_),
    .C(_2740_),
    .A(net935),
    .Y(_2741_));
 sg13g2_nand2_1 _6668_ (.Y(_2742_),
    .A(_3095_),
    .B(net968));
 sg13g2_xnor2_1 _6669_ (.Y(_2743_),
    .A(\vgademo.plane_dx[1] ),
    .B(net968));
 sg13g2_a21oi_1 _6670_ (.A1(net937),
    .A2(_2743_),
    .Y(_2744_),
    .B1(net899));
 sg13g2_a22oi_1 _6671_ (.Y(_0332_),
    .B1(_2741_),
    .B2(_2744_),
    .A2(net899),
    .A1(_3169_));
 sg13g2_nand2_1 _6672_ (.Y(_2745_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_xnor2_1 _6673_ (.Y(_2746_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_nand3_1 _6674_ (.B(_2740_),
    .C(_2746_),
    .A(_2737_),
    .Y(_2747_));
 sg13g2_a21o_1 _6675_ (.A2(_2740_),
    .A1(_2737_),
    .B1(_2746_),
    .X(_2748_));
 sg13g2_nor2_1 _6676_ (.A(\vgademo.plane_dx[2] ),
    .B(_2742_),
    .Y(_2749_));
 sg13g2_xnor2_1 _6677_ (.Y(_2750_),
    .A(\vgademo.plane_dx[2] ),
    .B(_2742_));
 sg13g2_a21oi_1 _6678_ (.A1(_2747_),
    .A2(_2748_),
    .Y(_2751_),
    .B1(net938));
 sg13g2_a21oi_1 _6679_ (.A1(net937),
    .A2(_2750_),
    .Y(_2752_),
    .B1(_2751_));
 sg13g2_mux2_1 _6680_ (.A0(net331),
    .A1(_2752_),
    .S(_2728_),
    .X(_0333_));
 sg13g2_xnor2_1 _6681_ (.Y(_2753_),
    .A(\vgademo.plane_u[4] ),
    .B(\vgademo.plane_du[4] ));
 sg13g2_nand3_1 _6682_ (.B(_2748_),
    .C(_2753_),
    .A(_2745_),
    .Y(_2754_));
 sg13g2_a21oi_1 _6683_ (.A1(_2745_),
    .A2(_2748_),
    .Y(_2755_),
    .B1(_2753_));
 sg13g2_nor2_1 _6684_ (.A(net937),
    .B(_2755_),
    .Y(_2756_));
 sg13g2_nor2_1 _6685_ (.A(\vgademo.plane_dx[3] ),
    .B(_2749_),
    .Y(_2757_));
 sg13g2_xnor2_1 _6686_ (.Y(_2758_),
    .A(\vgademo.plane_dx[3] ),
    .B(_2749_));
 sg13g2_a221oi_1 _6687_ (.B2(net937),
    .C1(net899),
    .B1(_2758_),
    .A1(_2754_),
    .Y(_2759_),
    .A2(_2756_));
 sg13g2_a21oi_1 _6688_ (.A1(_3170_),
    .A2(net899),
    .Y(_0334_),
    .B1(_2759_));
 sg13g2_a21o_1 _6689_ (.A2(\vgademo.plane_du[4] ),
    .A1(\vgademo.plane_u[4] ),
    .B1(_2755_),
    .X(_2760_));
 sg13g2_nand2_1 _6690_ (.Y(_2761_),
    .A(_3172_),
    .B(_3173_));
 sg13g2_nand2_1 _6691_ (.Y(_2762_),
    .A(\vgademo.plane_u[5] ),
    .B(\vgademo.plane_du[5] ));
 sg13g2_nand3_1 _6692_ (.B(_2761_),
    .C(_2762_),
    .A(_2760_),
    .Y(_2763_));
 sg13g2_a21oi_1 _6693_ (.A1(_2761_),
    .A2(_2762_),
    .Y(_2764_),
    .B1(_2760_));
 sg13g2_nor2_1 _6694_ (.A(net937),
    .B(_2764_),
    .Y(_2765_));
 sg13g2_nand2b_1 _6695_ (.Y(_2766_),
    .B(\vgademo.plane_dx[0] ),
    .A_N(_0023_));
 sg13g2_xnor2_1 _6696_ (.Y(_2767_),
    .A(\vgademo.plane_dx[0] ),
    .B(net1044));
 sg13g2_nand2_1 _6697_ (.Y(_2768_),
    .A(_0022_),
    .B(_2767_));
 sg13g2_xnor2_1 _6698_ (.Y(_2769_),
    .A(_0022_),
    .B(_2767_));
 sg13g2_a21oi_1 _6699_ (.A1(_2757_),
    .A2(_2769_),
    .Y(_2770_),
    .B1(net935));
 sg13g2_o21ai_1 _6700_ (.B1(_2770_),
    .Y(_2771_),
    .A1(_2757_),
    .A2(_2769_));
 sg13g2_a21oi_1 _6701_ (.A1(_2763_),
    .A2(_2765_),
    .Y(_2772_),
    .B1(net899));
 sg13g2_a22oi_1 _6702_ (.Y(_0335_),
    .B1(_2771_),
    .B2(_2772_),
    .A2(net899),
    .A1(_3172_));
 sg13g2_xnor2_1 _6703_ (.Y(_2773_),
    .A(\vgademo.plane_u[6] ),
    .B(\vgademo.plane_du[6] ));
 sg13g2_nand2_1 _6704_ (.Y(_2774_),
    .A(_2760_),
    .B(_2761_));
 sg13g2_nand3_1 _6705_ (.B(_2773_),
    .C(_2774_),
    .A(_2762_),
    .Y(_2775_));
 sg13g2_a21oi_1 _6706_ (.A1(_2762_),
    .A2(_2774_),
    .Y(_2776_),
    .B1(_2773_));
 sg13g2_nor2_1 _6707_ (.A(net937),
    .B(_2776_),
    .Y(_2777_));
 sg13g2_nand2_1 _6708_ (.Y(_2778_),
    .A(net1042),
    .B(\vgademo.plane_dx[1] ));
 sg13g2_xor2_1 _6709_ (.B(\vgademo.plane_dx[1] ),
    .A(net1043),
    .X(_2779_));
 sg13g2_nand2b_1 _6710_ (.Y(_2780_),
    .B(_2779_),
    .A_N(_2766_));
 sg13g2_xnor2_1 _6711_ (.Y(_2781_),
    .A(_2766_),
    .B(_2779_));
 sg13g2_xnor2_1 _6712_ (.Y(_2782_),
    .A(net968),
    .B(_2781_));
 sg13g2_nand2b_1 _6713_ (.Y(_2783_),
    .B(_2782_),
    .A_N(_2767_));
 sg13g2_xnor2_1 _6714_ (.Y(_2784_),
    .A(_2767_),
    .B(_2782_));
 sg13g2_o21ai_1 _6715_ (.B1(_2768_),
    .Y(_2785_),
    .A1(_2757_),
    .A2(_2769_));
 sg13g2_nand2_1 _6716_ (.Y(_2786_),
    .A(_2784_),
    .B(_2785_));
 sg13g2_nor2_1 _6717_ (.A(_2784_),
    .B(_2785_),
    .Y(_2787_));
 sg13g2_nor2_1 _6718_ (.A(net935),
    .B(_2787_),
    .Y(_2788_));
 sg13g2_a221oi_1 _6719_ (.B2(_2788_),
    .C1(net900),
    .B1(_2786_),
    .A1(_2775_),
    .Y(_2789_),
    .A2(_2777_));
 sg13g2_a21oi_1 _6720_ (.A1(_3174_),
    .A2(net899),
    .Y(_0336_),
    .B1(_2789_));
 sg13g2_xnor2_1 _6721_ (.Y(_2790_),
    .A(\vgademo.plane_u[7] ),
    .B(\vgademo.plane_du[7] ));
 sg13g2_a21oi_1 _6722_ (.A1(\vgademo.plane_u[6] ),
    .A2(\vgademo.plane_du[6] ),
    .Y(_2791_),
    .B1(_2776_));
 sg13g2_nand2_1 _6723_ (.Y(_2792_),
    .A(_2790_),
    .B(_2791_));
 sg13g2_nor2_1 _6724_ (.A(_2790_),
    .B(_2791_),
    .Y(_2793_));
 sg13g2_nor2_1 _6725_ (.A(net937),
    .B(_2793_),
    .Y(_2794_));
 sg13g2_nand2_1 _6726_ (.Y(_2795_),
    .A(\vgademo.plane_dx[0] ),
    .B(_2781_));
 sg13g2_xnor2_1 _6727_ (.Y(_2796_),
    .A(\vgademo.plane_dx_div.q[5] ),
    .B(\vgademo.plane_dx[2] ));
 sg13g2_a21oi_1 _6728_ (.A1(_2778_),
    .A2(_2780_),
    .Y(_2797_),
    .B1(_2796_));
 sg13g2_nand3_1 _6729_ (.B(_2780_),
    .C(_2796_),
    .A(_2778_),
    .Y(_2798_));
 sg13g2_nor2b_1 _6730_ (.A(_2797_),
    .B_N(_2798_),
    .Y(_2799_));
 sg13g2_xnor2_1 _6731_ (.Y(_2800_),
    .A(_0024_),
    .B(_2799_));
 sg13g2_nand2b_1 _6732_ (.Y(_2801_),
    .B(_2795_),
    .A_N(_2800_));
 sg13g2_xor2_1 _6733_ (.B(_2800_),
    .A(_2795_),
    .X(_2802_));
 sg13g2_nor2_1 _6734_ (.A(_2782_),
    .B(_2802_),
    .Y(_2803_));
 sg13g2_xnor2_1 _6735_ (.Y(_2804_),
    .A(_2782_),
    .B(_2802_));
 sg13g2_nand3_1 _6736_ (.B(_2786_),
    .C(_2804_),
    .A(_2783_),
    .Y(_2805_));
 sg13g2_a21o_1 _6737_ (.A2(_2786_),
    .A1(_2783_),
    .B1(_2804_),
    .X(_2806_));
 sg13g2_nand3_1 _6738_ (.B(_2805_),
    .C(_2806_),
    .A(net938),
    .Y(_2807_));
 sg13g2_a21oi_1 _6739_ (.A1(_2792_),
    .A2(_2794_),
    .Y(_2808_),
    .B1(net901));
 sg13g2_a22oi_1 _6740_ (.Y(_0337_),
    .B1(_2807_),
    .B2(_2808_),
    .A2(net898),
    .A1(_3175_));
 sg13g2_nand2_1 _6741_ (.Y(_2809_),
    .A(\vgademo.plane_u[8] ),
    .B(\vgademo.plane_du[8] ));
 sg13g2_nor2_1 _6742_ (.A(\vgademo.plane_u[8] ),
    .B(net963),
    .Y(_2810_));
 sg13g2_xor2_1 _6743_ (.B(net963),
    .A(\vgademo.plane_u[8] ),
    .X(_2811_));
 sg13g2_a21oi_1 _6744_ (.A1(\vgademo.plane_u[7] ),
    .A2(\vgademo.plane_du[7] ),
    .Y(_2812_),
    .B1(_2793_));
 sg13g2_xnor2_1 _6745_ (.Y(_2813_),
    .A(_2811_),
    .B(_2812_));
 sg13g2_nor2b_1 _6746_ (.A(_2803_),
    .B_N(_2806_),
    .Y(_2814_));
 sg13g2_nand2_1 _6747_ (.Y(_2815_),
    .A(\vgademo.plane_dx[1] ),
    .B(_2799_));
 sg13g2_a21oi_1 _6748_ (.A1(\vgademo.plane_dx_div.q[5] ),
    .A2(_3178_),
    .Y(_2816_),
    .B1(_2797_));
 sg13g2_xor2_1 _6749_ (.B(\vgademo.plane_dx[3] ),
    .A(net1040),
    .X(_2817_));
 sg13g2_nand2b_1 _6750_ (.Y(_2818_),
    .B(_2817_),
    .A_N(_2816_));
 sg13g2_xnor2_1 _6751_ (.Y(_2819_),
    .A(_2816_),
    .B(_2817_));
 sg13g2_xnor2_1 _6752_ (.Y(_2820_),
    .A(_0025_),
    .B(_2819_));
 sg13g2_nand2b_1 _6753_ (.Y(_2821_),
    .B(_2815_),
    .A_N(_2820_));
 sg13g2_xor2_1 _6754_ (.B(_2820_),
    .A(_2815_),
    .X(_2822_));
 sg13g2_xnor2_1 _6755_ (.Y(_2823_),
    .A(_2801_),
    .B(_2822_));
 sg13g2_or2_1 _6756_ (.X(_2824_),
    .B(_2823_),
    .A(_2814_));
 sg13g2_a21oi_1 _6757_ (.A1(_2814_),
    .A2(_2823_),
    .Y(_2825_),
    .B1(net935));
 sg13g2_a221oi_1 _6758_ (.B2(_2825_),
    .C1(net898),
    .B1(_2824_),
    .A1(net935),
    .Y(_2826_),
    .A2(_2813_));
 sg13g2_a21oi_1 _6759_ (.A1(_3177_),
    .A2(net901),
    .Y(_0338_),
    .B1(_2826_));
 sg13g2_nand2_1 _6760_ (.Y(_2827_),
    .A(net353),
    .B(\vgademo.plane_du[9] ));
 sg13g2_xnor2_1 _6761_ (.Y(_2828_),
    .A(\vgademo.plane_u[9] ),
    .B(net962));
 sg13g2_o21ai_1 _6762_ (.B1(_2809_),
    .Y(_2829_),
    .A1(_2810_),
    .A2(_2812_));
 sg13g2_xnor2_1 _6763_ (.Y(_2830_),
    .A(_2828_),
    .B(_2829_));
 sg13g2_o21ai_1 _6764_ (.B1(_2824_),
    .Y(_2831_),
    .A1(_2801_),
    .A2(_2822_));
 sg13g2_xor2_1 _6765_ (.B(net968),
    .A(\vgademo.plane_dx[3] ),
    .X(_2832_));
 sg13g2_nor2_1 _6766_ (.A(net1044),
    .B(_0026_),
    .Y(_2833_));
 sg13g2_nand2_1 _6767_ (.Y(_2834_),
    .A(net1044),
    .B(_0026_));
 sg13g2_nand2b_1 _6768_ (.Y(_2835_),
    .B(_2834_),
    .A_N(_2833_));
 sg13g2_o21ai_1 _6769_ (.B1(_2818_),
    .Y(_2836_),
    .A1(_3093_),
    .A2(_0022_));
 sg13g2_xnor2_1 _6770_ (.Y(_2837_),
    .A(_2835_),
    .B(_2836_));
 sg13g2_nor2_1 _6771_ (.A(_2832_),
    .B(_2837_),
    .Y(_2838_));
 sg13g2_xnor2_1 _6772_ (.Y(_2839_),
    .A(_2832_),
    .B(_2837_));
 sg13g2_nand2_1 _6773_ (.Y(_2840_),
    .A(\vgademo.plane_dx[2] ),
    .B(_2819_));
 sg13g2_nand2b_1 _6774_ (.Y(_2841_),
    .B(_2840_),
    .A_N(_2839_));
 sg13g2_xor2_1 _6775_ (.B(_2840_),
    .A(_2839_),
    .X(_2842_));
 sg13g2_xor2_1 _6776_ (.B(_2842_),
    .A(_2821_),
    .X(_2843_));
 sg13g2_nor2_1 _6777_ (.A(_2831_),
    .B(_2843_),
    .Y(_2844_));
 sg13g2_nand2_1 _6778_ (.Y(_2845_),
    .A(_2831_),
    .B(_2843_));
 sg13g2_nor2_1 _6779_ (.A(net933),
    .B(_2844_),
    .Y(_2846_));
 sg13g2_a221oi_1 _6780_ (.B2(_2846_),
    .C1(net898),
    .B1(_2845_),
    .A1(net933),
    .Y(_2847_),
    .A2(_2830_));
 sg13g2_a21oi_1 _6781_ (.A1(_3179_),
    .A2(net898),
    .Y(_0339_),
    .B1(_2847_));
 sg13g2_nand2_1 _6782_ (.Y(_2848_),
    .A(\vgademo.plane_u[10] ),
    .B(\vgademo.plane_du[10] ));
 sg13g2_xnor2_1 _6783_ (.Y(_2849_),
    .A(\vgademo.plane_u[10] ),
    .B(\vgademo.plane_du[10] ));
 sg13g2_o21ai_1 _6784_ (.B1(_2829_),
    .Y(_2850_),
    .A1(\vgademo.plane_u[9] ),
    .A2(net962));
 sg13g2_nand3_1 _6785_ (.B(_2849_),
    .C(_2850_),
    .A(_2827_),
    .Y(_2851_));
 sg13g2_a21o_1 _6786_ (.A2(_2850_),
    .A1(_2827_),
    .B1(_2849_),
    .X(_2852_));
 sg13g2_nand3_1 _6787_ (.B(_2851_),
    .C(_2852_),
    .A(net933),
    .Y(_2853_));
 sg13g2_o21ai_1 _6788_ (.B1(_2845_),
    .Y(_2854_),
    .A1(_2821_),
    .A2(_2842_));
 sg13g2_xor2_1 _6789_ (.B(net1044),
    .A(\vgademo.plane_dx[1] ),
    .X(_2855_));
 sg13g2_a21oi_1 _6790_ (.A1(_2834_),
    .A2(_2836_),
    .Y(_2856_),
    .B1(_2833_));
 sg13g2_nand2_1 _6791_ (.Y(_2857_),
    .A(net1037),
    .B(net1043));
 sg13g2_nor2_1 _6792_ (.A(net1037),
    .B(net1043),
    .Y(_2858_));
 sg13g2_xor2_1 _6793_ (.B(net1043),
    .A(net1037),
    .X(_2859_));
 sg13g2_xnor2_1 _6794_ (.Y(_2860_),
    .A(_2856_),
    .B(_2859_));
 sg13g2_nor2_1 _6795_ (.A(_2855_),
    .B(_2860_),
    .Y(_2861_));
 sg13g2_xor2_1 _6796_ (.B(_2860_),
    .A(_2855_),
    .X(_2862_));
 sg13g2_a21oi_1 _6797_ (.A1(_3094_),
    .A2(net968),
    .Y(_2863_),
    .B1(_2838_));
 sg13g2_nand2b_1 _6798_ (.Y(_2864_),
    .B(_2862_),
    .A_N(_2863_));
 sg13g2_xor2_1 _6799_ (.B(_2863_),
    .A(_2862_),
    .X(_2865_));
 sg13g2_nor2_1 _6800_ (.A(_2841_),
    .B(_2865_),
    .Y(_2866_));
 sg13g2_xor2_1 _6801_ (.B(_2865_),
    .A(_2841_),
    .X(_2867_));
 sg13g2_nor2_1 _6802_ (.A(_2854_),
    .B(_2867_),
    .Y(_2868_));
 sg13g2_nand2_1 _6803_ (.Y(_2869_),
    .A(_2854_),
    .B(_2867_));
 sg13g2_nor2_1 _6804_ (.A(net933),
    .B(_2868_),
    .Y(_2870_));
 sg13g2_a21oi_1 _6805_ (.A1(_2869_),
    .A2(_2870_),
    .Y(_2871_),
    .B1(net898));
 sg13g2_a22oi_1 _6806_ (.Y(_0340_),
    .B1(_2853_),
    .B2(_2871_),
    .A2(net898),
    .A1(_3180_));
 sg13g2_a21oi_2 _6807_ (.B1(_0027_),
    .Y(_2872_),
    .A2(_2852_),
    .A1(_2848_));
 sg13g2_nand3_1 _6808_ (.B(_2848_),
    .C(_2852_),
    .A(_0027_),
    .Y(_2873_));
 sg13g2_nor2_1 _6809_ (.A(net938),
    .B(_2872_),
    .Y(_2874_));
 sg13g2_a21oi_1 _6810_ (.A1(_2854_),
    .A2(_2867_),
    .Y(_2875_),
    .B1(_2866_));
 sg13g2_xnor2_1 _6811_ (.Y(_2876_),
    .A(\vgademo.plane_dx_div.q[9] ),
    .B(\vgademo.plane_dx_div.q[5] ));
 sg13g2_o21ai_1 _6812_ (.B1(_2857_),
    .Y(_2877_),
    .A1(_2856_),
    .A2(_2858_));
 sg13g2_nor2b_1 _6813_ (.A(_2876_),
    .B_N(_2877_),
    .Y(_2878_));
 sg13g2_xor2_1 _6814_ (.B(_2877_),
    .A(_2876_),
    .X(_2879_));
 sg13g2_xor2_1 _6815_ (.B(\vgademo.plane_dx[2] ),
    .A(net1042),
    .X(_2880_));
 sg13g2_nand2_1 _6816_ (.Y(_2881_),
    .A(_2879_),
    .B(_2880_));
 sg13g2_xnor2_1 _6817_ (.Y(_2882_),
    .A(_2879_),
    .B(_2880_));
 sg13g2_a21oi_1 _6818_ (.A1(net1044),
    .A2(_0024_),
    .Y(_2883_),
    .B1(_2861_));
 sg13g2_nor2_1 _6819_ (.A(_2882_),
    .B(_2883_),
    .Y(_2884_));
 sg13g2_xnor2_1 _6820_ (.Y(_2885_),
    .A(_2882_),
    .B(_2883_));
 sg13g2_xnor2_1 _6821_ (.Y(_2886_),
    .A(_2864_),
    .B(_2885_));
 sg13g2_nor2_1 _6822_ (.A(_2875_),
    .B(_2886_),
    .Y(_2887_));
 sg13g2_inv_1 _6823_ (.Y(_2888_),
    .A(_2887_));
 sg13g2_a21oi_1 _6824_ (.A1(_2875_),
    .A2(_2886_),
    .Y(_2889_),
    .B1(net933));
 sg13g2_a221oi_1 _6825_ (.B2(_2889_),
    .C1(net898),
    .B1(_2888_),
    .A1(_2873_),
    .Y(_2890_),
    .A2(_2874_));
 sg13g2_a21oi_1 _6826_ (.A1(_3181_),
    .A2(net898),
    .Y(_0341_),
    .B1(_2890_));
 sg13g2_a21oi_1 _6827_ (.A1(_0028_),
    .A2(_2872_),
    .Y(_2891_),
    .B1(net939));
 sg13g2_o21ai_1 _6828_ (.B1(_2891_),
    .Y(_2892_),
    .A1(_0028_),
    .A2(_2872_));
 sg13g2_o21ai_1 _6829_ (.B1(_2888_),
    .Y(_2893_),
    .A1(_2864_),
    .A2(_2885_));
 sg13g2_a21oi_1 _6830_ (.A1(net1036),
    .A2(net1041),
    .Y(_2894_),
    .B1(_2878_));
 sg13g2_nand2b_2 _6831_ (.Y(_2895_),
    .B(net1040),
    .A_N(_2894_));
 sg13g2_xnor2_1 _6832_ (.Y(_2896_),
    .A(net1040),
    .B(_2894_));
 sg13g2_xor2_1 _6833_ (.B(\vgademo.plane_dx[3] ),
    .A(net1041),
    .X(_2897_));
 sg13g2_nand2b_1 _6834_ (.Y(_2898_),
    .B(_2897_),
    .A_N(_2896_));
 sg13g2_xnor2_1 _6835_ (.Y(_2899_),
    .A(_2896_),
    .B(_2897_));
 sg13g2_o21ai_1 _6836_ (.B1(_2881_),
    .Y(_2900_),
    .A1(net1042),
    .A2(_3178_));
 sg13g2_nand2_1 _6837_ (.Y(_2901_),
    .A(_2899_),
    .B(_2900_));
 sg13g2_xor2_1 _6838_ (.B(_2900_),
    .A(_2899_),
    .X(_2902_));
 sg13g2_xnor2_1 _6839_ (.Y(_2903_),
    .A(_2884_),
    .B(_2902_));
 sg13g2_nor2b_1 _6840_ (.A(_2903_),
    .B_N(_2893_),
    .Y(_2904_));
 sg13g2_xor2_1 _6841_ (.B(_2903_),
    .A(_2893_),
    .X(_2905_));
 sg13g2_a21oi_1 _6842_ (.A1(net939),
    .A2(_2905_),
    .Y(_2906_),
    .B1(net902));
 sg13g2_a22oi_1 _6843_ (.Y(_2907_),
    .B1(_2892_),
    .B2(_2906_),
    .A2(net902),
    .A1(net424));
 sg13g2_inv_1 _6844_ (.Y(_0342_),
    .A(net425));
 sg13g2_a21oi_1 _6845_ (.A1(_2884_),
    .A2(_2902_),
    .Y(_2908_),
    .B1(_2904_));
 sg13g2_nand2_1 _6846_ (.Y(_2909_),
    .A(_3093_),
    .B(net1044));
 sg13g2_xor2_1 _6847_ (.B(net1044),
    .A(net1040),
    .X(_2910_));
 sg13g2_nor2_1 _6848_ (.A(net1039),
    .B(_2895_),
    .Y(_2911_));
 sg13g2_xor2_1 _6849_ (.B(_2895_),
    .A(net1039),
    .X(_2912_));
 sg13g2_xnor2_1 _6850_ (.Y(_2913_),
    .A(_2910_),
    .B(_2912_));
 sg13g2_nand2b_1 _6851_ (.Y(_2914_),
    .B(_0022_),
    .A_N(net1041));
 sg13g2_and2_1 _6852_ (.A(_2898_),
    .B(_2914_),
    .X(_2915_));
 sg13g2_or2_1 _6853_ (.X(_2916_),
    .B(_2915_),
    .A(_2913_));
 sg13g2_xor2_1 _6854_ (.B(_2915_),
    .A(_2913_),
    .X(_2917_));
 sg13g2_nand2b_1 _6855_ (.Y(_2918_),
    .B(_2917_),
    .A_N(_2901_));
 sg13g2_xnor2_1 _6856_ (.Y(_2919_),
    .A(_2901_),
    .B(_2917_));
 sg13g2_nand2b_1 _6857_ (.Y(_2920_),
    .B(_2908_),
    .A_N(_2919_));
 sg13g2_nand2b_1 _6858_ (.Y(_2921_),
    .B(_2919_),
    .A_N(_2908_));
 sg13g2_nand3_1 _6859_ (.B(_2920_),
    .C(_2921_),
    .A(net939),
    .Y(_2922_));
 sg13g2_nand3_1 _6860_ (.B(\vgademo.plane_u[13] ),
    .C(_2872_),
    .A(\vgademo.plane_u[12] ),
    .Y(_2923_));
 sg13g2_a21oi_1 _6861_ (.A1(net424),
    .A2(_2872_),
    .Y(_2924_),
    .B1(net434));
 sg13g2_nor2_1 _6862_ (.A(net939),
    .B(_2924_),
    .Y(_2925_));
 sg13g2_a21oi_1 _6863_ (.A1(_2923_),
    .A2(_2925_),
    .Y(_2926_),
    .B1(net902));
 sg13g2_a22oi_1 _6864_ (.Y(_0343_),
    .B1(_2922_),
    .B2(_2926_),
    .A2(net902),
    .A1(_3182_));
 sg13g2_and2_1 _6865_ (.A(_2918_),
    .B(_2921_),
    .X(_2927_));
 sg13g2_nor2b_1 _6866_ (.A(net1042),
    .B_N(net1039),
    .Y(_2928_));
 sg13g2_xnor2_1 _6867_ (.Y(_2929_),
    .A(net1042),
    .B(net1039));
 sg13g2_nor3_1 _6868_ (.A(_3092_),
    .B(net1039),
    .C(_2895_),
    .Y(_2930_));
 sg13g2_xnor2_1 _6869_ (.Y(_2931_),
    .A(net1037),
    .B(_2911_));
 sg13g2_xor2_1 _6870_ (.B(_2931_),
    .A(_2929_),
    .X(_2932_));
 sg13g2_o21ai_1 _6871_ (.B1(_2909_),
    .Y(_2933_),
    .A1(_2910_),
    .A2(_2912_));
 sg13g2_nand2_1 _6872_ (.Y(_2934_),
    .A(_2932_),
    .B(_2933_));
 sg13g2_xnor2_1 _6873_ (.Y(_2935_),
    .A(_2932_),
    .B(_2933_));
 sg13g2_nor2_1 _6874_ (.A(_2916_),
    .B(_2935_),
    .Y(_2936_));
 sg13g2_xor2_1 _6875_ (.B(_2935_),
    .A(_2916_),
    .X(_2937_));
 sg13g2_nor2b_1 _6876_ (.A(_2927_),
    .B_N(_2937_),
    .Y(_2938_));
 sg13g2_xor2_1 _6877_ (.B(_2937_),
    .A(_2927_),
    .X(_2939_));
 sg13g2_xnor2_1 _6878_ (.Y(_2940_),
    .A(_3183_),
    .B(_2923_));
 sg13g2_nand2_1 _6879_ (.Y(_2941_),
    .A(net936),
    .B(_2940_));
 sg13g2_a21oi_1 _6880_ (.A1(net940),
    .A2(_2939_),
    .Y(_2942_),
    .B1(net897));
 sg13g2_a22oi_1 _6881_ (.Y(_2943_),
    .B1(_2941_),
    .B2(_2942_),
    .A2(net897),
    .A1(net392));
 sg13g2_inv_1 _6882_ (.Y(_0344_),
    .A(_2943_));
 sg13g2_nor2_1 _6883_ (.A(net1038),
    .B(net1041),
    .Y(_2944_));
 sg13g2_xor2_1 _6884_ (.B(net1041),
    .A(net1038),
    .X(_2945_));
 sg13g2_xnor2_1 _6885_ (.Y(_2946_),
    .A(\vgademo.plane_dx_div.q[9] ),
    .B(_2930_));
 sg13g2_xnor2_1 _6886_ (.Y(_2947_),
    .A(_2945_),
    .B(_2946_));
 sg13g2_a21oi_1 _6887_ (.A1(_2929_),
    .A2(_2931_),
    .Y(_2948_),
    .B1(_2928_));
 sg13g2_nor2_1 _6888_ (.A(_2947_),
    .B(_2948_),
    .Y(_2949_));
 sg13g2_xor2_1 _6889_ (.B(_2948_),
    .A(_2947_),
    .X(_2950_));
 sg13g2_nand2b_1 _6890_ (.Y(_2951_),
    .B(_2950_),
    .A_N(_2934_));
 sg13g2_xnor2_1 _6891_ (.Y(_2952_),
    .A(_2934_),
    .B(_2950_));
 sg13g2_o21ai_1 _6892_ (.B1(_2952_),
    .Y(_2953_),
    .A1(_2936_),
    .A2(_2938_));
 sg13g2_nor3_1 _6893_ (.A(_2936_),
    .B(_2938_),
    .C(_2952_),
    .Y(_2954_));
 sg13g2_nor2_1 _6894_ (.A(net936),
    .B(_2954_),
    .Y(_2955_));
 sg13g2_nor2_1 _6895_ (.A(_0029_),
    .B(_2923_),
    .Y(_2956_));
 sg13g2_xnor2_1 _6896_ (.Y(_2957_),
    .A(_3184_),
    .B(_2956_));
 sg13g2_a221oi_1 _6897_ (.B2(net936),
    .C1(net897),
    .B1(_2957_),
    .A1(_2953_),
    .Y(_2958_),
    .A2(_2955_));
 sg13g2_a21oi_1 _6898_ (.A1(_3184_),
    .A2(net897),
    .Y(_0345_),
    .B1(_2958_));
 sg13g2_nand2_1 _6899_ (.Y(_2959_),
    .A(net1036),
    .B(net1040));
 sg13g2_or2_1 _6900_ (.X(_2960_),
    .B(net1040),
    .A(net1036));
 sg13g2_a21oi_1 _6901_ (.A1(_2959_),
    .A2(_2960_),
    .Y(_2961_),
    .B1(_2930_));
 sg13g2_a21oi_1 _6902_ (.A1(_2945_),
    .A2(_2946_),
    .Y(_2962_),
    .B1(_2944_));
 sg13g2_nor2b_1 _6903_ (.A(_2962_),
    .B_N(_2961_),
    .Y(_2963_));
 sg13g2_xnor2_1 _6904_ (.Y(_2964_),
    .A(_2961_),
    .B(_2962_));
 sg13g2_xnor2_1 _6905_ (.Y(_2965_),
    .A(_2949_),
    .B(_2964_));
 sg13g2_a21oi_1 _6906_ (.A1(_2951_),
    .A2(_2953_),
    .Y(_2966_),
    .B1(_2965_));
 sg13g2_and3_1 _6907_ (.X(_2967_),
    .A(_2951_),
    .B(_2953_),
    .C(_2965_));
 sg13g2_nor3_2 _6908_ (.A(_3183_),
    .B(_3184_),
    .C(_2923_),
    .Y(_2968_));
 sg13g2_o21ai_1 _6909_ (.B1(net940),
    .Y(_2969_),
    .A1(_2966_),
    .A2(_2967_));
 sg13g2_xor2_1 _6910_ (.B(_2968_),
    .A(_0030_),
    .X(_2970_));
 sg13g2_a21oi_1 _6911_ (.A1(net936),
    .A2(_2970_),
    .Y(_2971_),
    .B1(net896));
 sg13g2_a22oi_1 _6912_ (.Y(_2972_),
    .B1(_2969_),
    .B2(_2971_),
    .A2(net896),
    .A1(net364));
 sg13g2_inv_1 _6913_ (.Y(_0346_),
    .A(net365));
 sg13g2_a21oi_1 _6914_ (.A1(_2949_),
    .A2(_2964_),
    .Y(_2973_),
    .B1(_2966_));
 sg13g2_nand2_1 _6915_ (.Y(_2974_),
    .A(net1039),
    .B(_2959_));
 sg13g2_xor2_1 _6916_ (.B(_2959_),
    .A(net1039),
    .X(_2975_));
 sg13g2_xnor2_1 _6917_ (.Y(_2976_),
    .A(_2963_),
    .B(_2975_));
 sg13g2_nor2_1 _6918_ (.A(_2973_),
    .B(_2976_),
    .Y(_2977_));
 sg13g2_a21oi_1 _6919_ (.A1(_2973_),
    .A2(_2976_),
    .Y(_2978_),
    .B1(net936));
 sg13g2_nand2b_1 _6920_ (.Y(_2979_),
    .B(_2978_),
    .A_N(_2977_));
 sg13g2_and3_1 _6921_ (.X(_2980_),
    .A(\vgademo.plane_u[16] ),
    .B(\vgademo.plane_u[17] ),
    .C(_2968_));
 sg13g2_a21oi_1 _6922_ (.A1(net364),
    .A2(_2968_),
    .Y(_2981_),
    .B1(net426));
 sg13g2_nor3_1 _6923_ (.A(net940),
    .B(_2980_),
    .C(_2981_),
    .Y(_2982_));
 sg13g2_nor2_1 _6924_ (.A(net896),
    .B(_2982_),
    .Y(_2983_));
 sg13g2_a22oi_1 _6925_ (.Y(_0347_),
    .B1(_2979_),
    .B2(_2983_),
    .A2(net896),
    .A1(_3185_));
 sg13g2_a21oi_1 _6926_ (.A1(_2963_),
    .A2(_2975_),
    .Y(_2984_),
    .B1(_2977_));
 sg13g2_xnor2_1 _6927_ (.Y(_2985_),
    .A(_3092_),
    .B(_2974_));
 sg13g2_or2_1 _6928_ (.X(_2986_),
    .B(_2985_),
    .A(_2984_));
 sg13g2_a21oi_1 _6929_ (.A1(_2984_),
    .A2(_2985_),
    .Y(_2987_),
    .B1(net931));
 sg13g2_xnor2_1 _6930_ (.Y(_2988_),
    .A(_3186_),
    .B(_2980_));
 sg13g2_a221oi_1 _6931_ (.B2(net931),
    .C1(net895),
    .B1(_2988_),
    .A1(_2986_),
    .Y(_2989_),
    .A2(_2987_));
 sg13g2_a21oi_1 _6932_ (.A1(_3186_),
    .A2(net895),
    .Y(_0348_),
    .B1(_2989_));
 sg13g2_o21ai_1 _6933_ (.B1(_2986_),
    .Y(_2990_),
    .A1(_3092_),
    .A2(_2974_));
 sg13g2_xnor2_1 _6934_ (.Y(_2991_),
    .A(net1036),
    .B(net1037));
 sg13g2_xnor2_1 _6935_ (.Y(_2992_),
    .A(_2990_),
    .B(_2991_));
 sg13g2_nand2_1 _6936_ (.Y(_2993_),
    .A(net941),
    .B(_2992_));
 sg13g2_nor2b_1 _6937_ (.A(_0031_),
    .B_N(_2980_),
    .Y(_2994_));
 sg13g2_xnor2_1 _6938_ (.Y(_2995_),
    .A(net419),
    .B(_2994_));
 sg13g2_a21oi_1 _6939_ (.A1(net931),
    .A2(_2995_),
    .Y(_2996_),
    .B1(net895));
 sg13g2_a22oi_1 _6940_ (.Y(_2997_),
    .B1(_2993_),
    .B2(_2996_),
    .A2(net895),
    .A1(net419));
 sg13g2_inv_1 _6941_ (.Y(_0349_),
    .A(net420));
 sg13g2_nand4_1 _6942_ (.B(net1037),
    .C(_2974_),
    .A(net1036),
    .Y(_2998_),
    .D(_2984_));
 sg13g2_nor3_1 _6943_ (.A(net1036),
    .B(net1037),
    .C(_2986_),
    .Y(_2999_));
 sg13g2_nor2_1 _6944_ (.A(net931),
    .B(_2999_),
    .Y(_3000_));
 sg13g2_nand2b_1 _6945_ (.Y(_3001_),
    .B(net941),
    .A_N(_2999_));
 sg13g2_nand3_1 _6946_ (.B(\vgademo.plane_u[19] ),
    .C(_2980_),
    .A(\vgademo.plane_u[18] ),
    .Y(_3002_));
 sg13g2_xnor2_1 _6947_ (.Y(_3003_),
    .A(net255),
    .B(_3002_));
 sg13g2_a221oi_1 _6948_ (.B2(net931),
    .C1(net895),
    .B1(_3003_),
    .A1(_2998_),
    .Y(_3004_),
    .A2(_3000_));
 sg13g2_a21oi_1 _6949_ (.A1(_3187_),
    .A2(net895),
    .Y(_0350_),
    .B1(_3004_));
 sg13g2_nor2_1 _6950_ (.A(_0032_),
    .B(_3002_),
    .Y(_3005_));
 sg13g2_xnor2_1 _6951_ (.Y(_3006_),
    .A(_3188_),
    .B(_3005_));
 sg13g2_a21oi_1 _6952_ (.A1(net931),
    .A2(_3006_),
    .Y(_3007_),
    .B1(net895));
 sg13g2_a22oi_1 _6953_ (.Y(_0351_),
    .B1(_3001_),
    .B2(_3007_),
    .A2(net895),
    .A1(_3188_));
 sg13g2_o21ai_1 _6954_ (.B1(_1861_),
    .Y(_3008_),
    .A1(_1810_),
    .A2(_1828_));
 sg13g2_and3_1 _6955_ (.X(_3009_),
    .A(net873),
    .B(net832),
    .C(_3008_));
 sg13g2_o21ai_1 _6956_ (.B1(net836),
    .Y(_3010_),
    .A1(_2142_),
    .A2(_3009_));
 sg13g2_a21oi_2 _6957_ (.B1(_1298_),
    .Y(_3011_),
    .A2(_3010_),
    .A1(_2180_));
 sg13g2_nor2_1 _6958_ (.A(_2162_),
    .B(_2183_),
    .Y(_3012_));
 sg13g2_o21ai_1 _6959_ (.B1(net833),
    .Y(_3013_),
    .A1(_2162_),
    .A2(_2183_));
 sg13g2_a21oi_1 _6960_ (.A1(net872),
    .A2(_3013_),
    .Y(_3014_),
    .B1(_2589_));
 sg13g2_nand2b_1 _6961_ (.Y(_3015_),
    .B(_2156_),
    .A_N(_2178_));
 sg13g2_a21oi_1 _6962_ (.A1(_2591_),
    .A2(_3015_),
    .Y(_3016_),
    .B1(_3014_));
 sg13g2_a21oi_2 _6963_ (.B1(_1298_),
    .Y(_3017_),
    .A2(_3016_),
    .A1(_1275_));
 sg13g2_o21ai_1 _6964_ (.B1(_3011_),
    .Y(_3018_),
    .A1(_2173_),
    .A2(_3017_));
 sg13g2_and2_1 _6965_ (.A(_2173_),
    .B(_3017_),
    .X(_3019_));
 sg13g2_o21ai_1 _6966_ (.B1(_3018_),
    .Y(_3020_),
    .A1(_3011_),
    .A2(_3019_));
 sg13g2_xor2_1 _6967_ (.B(_1804_),
    .A(_1791_),
    .X(_3021_));
 sg13g2_a21o_2 _6968_ (.A2(_3021_),
    .A1(_2184_),
    .B1(_2188_),
    .X(_3022_));
 sg13g2_mux2_1 _6969_ (.A0(_3008_),
    .A1(_3022_),
    .S(net833),
    .X(_3023_));
 sg13g2_or2_1 _6970_ (.X(_3024_),
    .B(_2192_),
    .A(_1756_));
 sg13g2_a21oi_1 _6971_ (.A1(net873),
    .A2(_3023_),
    .Y(_3025_),
    .B1(_3024_));
 sg13g2_o21ai_1 _6972_ (.B1(_1275_),
    .Y(_3026_),
    .A1(_2610_),
    .A2(_3025_));
 sg13g2_and2_1 _6973_ (.A(net953),
    .B(_3026_),
    .X(_3027_));
 sg13g2_or2_1 _6974_ (.X(_3028_),
    .B(_3026_),
    .A(net953));
 sg13g2_xnor2_1 _6975_ (.Y(_3029_),
    .A(_2171_),
    .B(_3026_));
 sg13g2_a21oi_1 _6976_ (.A1(_3017_),
    .A2(_3028_),
    .Y(_3030_),
    .B1(_3027_));
 sg13g2_xnor2_1 _6977_ (.Y(_3031_),
    .A(_2172_),
    .B(_3017_));
 sg13g2_xnor2_1 _6978_ (.Y(_3032_),
    .A(_3011_),
    .B(_3031_));
 sg13g2_nand2_1 _6979_ (.Y(_3033_),
    .A(_3030_),
    .B(_3032_));
 sg13g2_xnor2_1 _6980_ (.Y(_3034_),
    .A(_1796_),
    .B(_1800_));
 sg13g2_a21oi_1 _6981_ (.A1(_2184_),
    .A2(_3034_),
    .Y(_3035_),
    .B1(_2222_));
 sg13g2_nand3_1 _6982_ (.B(_1793_),
    .C(_1802_),
    .A(_1792_),
    .Y(_3036_));
 sg13g2_nor2b_1 _6983_ (.A(_1803_),
    .B_N(_3036_),
    .Y(_3037_));
 sg13g2_a21oi_2 _6984_ (.B1(_2219_),
    .Y(_3038_),
    .A2(_3037_),
    .A1(_2184_));
 sg13g2_mux2_1 _6985_ (.A0(_3038_),
    .A1(_3035_),
    .S(net833),
    .X(_3039_));
 sg13g2_a21oi_1 _6986_ (.A1(net873),
    .A2(_3039_),
    .Y(_3040_),
    .B1(_2203_));
 sg13g2_nor2_1 _6987_ (.A(net879),
    .B(_3040_),
    .Y(_3041_));
 sg13g2_nor2b_1 _6988_ (.A(_3041_),
    .B_N(net951),
    .Y(_3042_));
 sg13g2_nand3_1 _6989_ (.B(_1795_),
    .C(_1801_),
    .A(_1794_),
    .Y(_3043_));
 sg13g2_nand2_2 _6990_ (.Y(_3044_),
    .A(_1802_),
    .B(_3043_));
 sg13g2_o21ai_1 _6991_ (.B1(_2211_),
    .Y(_3045_),
    .A1(_2185_),
    .A2(_3044_));
 sg13g2_mux2_1 _6992_ (.A0(_3022_),
    .A1(_3045_),
    .S(net833),
    .X(_3046_));
 sg13g2_nor2_1 _6993_ (.A(net866),
    .B(_3046_),
    .Y(_3047_));
 sg13g2_o21ai_1 _6994_ (.B1(_1275_),
    .Y(_3048_),
    .A1(_2205_),
    .A2(_3047_));
 sg13g2_nand2b_1 _6995_ (.Y(_3049_),
    .B(_3041_),
    .A_N(net952));
 sg13g2_xor2_1 _6996_ (.B(_3041_),
    .A(net952),
    .X(_3050_));
 sg13g2_a21o_1 _6997_ (.A2(_3049_),
    .A1(_3048_),
    .B1(_3042_),
    .X(_3051_));
 sg13g2_mux2_1 _6998_ (.A0(_3012_),
    .A1(_3038_),
    .S(net833),
    .X(_3052_));
 sg13g2_a21o_1 _6999_ (.A2(_3052_),
    .A1(net871),
    .B1(_2236_),
    .X(_3053_));
 sg13g2_a21o_1 _7000_ (.A2(_3053_),
    .A1(_2158_),
    .B1(_1298_),
    .X(_3054_));
 sg13g2_nor2_1 _7001_ (.A(_2251_),
    .B(_3054_),
    .Y(_3055_));
 sg13g2_xnor2_1 _7002_ (.Y(_3056_),
    .A(_2252_),
    .B(_3054_));
 sg13g2_xor2_1 _7003_ (.B(_3056_),
    .A(_3026_),
    .X(_3057_));
 sg13g2_nor2_1 _7004_ (.A(_2243_),
    .B(_3011_),
    .Y(_3058_));
 sg13g2_a21oi_1 _7005_ (.A1(_2243_),
    .A2(_3011_),
    .Y(_3059_),
    .B1(_3048_));
 sg13g2_nor3_1 _7006_ (.A(_3054_),
    .B(_3058_),
    .C(_3059_),
    .Y(_3060_));
 sg13g2_o21ai_1 _7007_ (.B1(_3054_),
    .Y(_3061_),
    .A1(_3058_),
    .A2(_3059_));
 sg13g2_xnor2_1 _7008_ (.Y(_3062_),
    .A(_3048_),
    .B(_3050_));
 sg13g2_a221oi_1 _7009_ (.B2(_3062_),
    .C1(_3060_),
    .B1(_3061_),
    .A1(_3051_),
    .Y(_3063_),
    .A2(_3057_));
 sg13g2_xnor2_1 _7010_ (.Y(_3064_),
    .A(_3017_),
    .B(_3029_));
 sg13g2_a21o_1 _7011_ (.A2(_3056_),
    .A1(_3026_),
    .B1(_3055_),
    .X(_3065_));
 sg13g2_nor2_1 _7012_ (.A(_3064_),
    .B(_3065_),
    .Y(_3066_));
 sg13g2_nor2_1 _7013_ (.A(_3051_),
    .B(_3057_),
    .Y(_3067_));
 sg13g2_nor3_1 _7014_ (.A(_3063_),
    .B(_3066_),
    .C(_3067_),
    .Y(_3068_));
 sg13g2_nand2_1 _7015_ (.Y(_3069_),
    .A(_3064_),
    .B(_3065_));
 sg13g2_o21ai_1 _7016_ (.B1(_3069_),
    .Y(_3070_),
    .A1(_3030_),
    .A2(_3032_));
 sg13g2_o21ai_1 _7017_ (.B1(_3033_),
    .Y(_3071_),
    .A1(_3068_),
    .A2(_3070_));
 sg13g2_or2_1 _7018_ (.X(_3072_),
    .B(_3071_),
    .A(_3020_));
 sg13g2_a21oi_1 _7019_ (.A1(_3020_),
    .A2(_3071_),
    .Y(_3073_),
    .B1(_2274_));
 sg13g2_and2_1 _7020_ (.A(_3072_),
    .B(_3073_),
    .X(_0352_));
 sg13g2_a21oi_1 _7021_ (.A1(_3018_),
    .A2(_3072_),
    .Y(_0353_),
    .B1(_2274_));
 sg13g2_nor2_1 _7022_ (.A(net290),
    .B(net911),
    .Y(_3074_));
 sg13g2_a21oi_1 _7023_ (.A1(_3096_),
    .A2(net910),
    .Y(_0354_),
    .B1(_3074_));
 sg13g2_nor2_1 _7024_ (.A(net310),
    .B(net910),
    .Y(_3075_));
 sg13g2_a21oi_1 _7025_ (.A1(_3095_),
    .A2(net910),
    .Y(_0355_),
    .B1(_3075_));
 sg13g2_mux2_1 _7026_ (.A0(net483),
    .A1(\vgademo.plane_dx[2] ),
    .S(net910),
    .X(_0356_));
 sg13g2_nor2_1 _7027_ (.A(net541),
    .B(net910),
    .Y(_3076_));
 sg13g2_a21oi_1 _7028_ (.A1(_3094_),
    .A2(net910),
    .Y(_0357_),
    .B1(_3076_));
 sg13g2_nor2_1 _7029_ (.A(\vgademo.plane_du[4] ),
    .B(net911),
    .Y(_3077_));
 sg13g2_a21oi_1 _7030_ (.A1(net1044),
    .A2(net910),
    .Y(_0358_),
    .B1(_3077_));
 sg13g2_nand2_1 _7031_ (.Y(_3078_),
    .A(net1042),
    .B(net909));
 sg13g2_o21ai_1 _7032_ (.B1(_3078_),
    .Y(_0359_),
    .A1(_3173_),
    .A2(net909));
 sg13g2_mux2_1 _7033_ (.A0(net583),
    .A1(net1041),
    .S(net909),
    .X(_0360_));
 sg13g2_nor2_1 _7034_ (.A(\vgademo.plane_du[7] ),
    .B(net909),
    .Y(_3079_));
 sg13g2_a21oi_1 _7035_ (.A1(_3093_),
    .A2(net911),
    .Y(_0361_),
    .B1(_3079_));
 sg13g2_nor2_1 _7036_ (.A(net963),
    .B(net909),
    .Y(_3080_));
 sg13g2_a21oi_1 _7037_ (.A1(net1039),
    .A2(net909),
    .Y(_0362_),
    .B1(_3080_));
 sg13g2_nor2_1 _7038_ (.A(net962),
    .B(net909),
    .Y(_3081_));
 sg13g2_a21oi_1 _7039_ (.A1(_3092_),
    .A2(net909),
    .Y(_0363_),
    .B1(_3081_));
 sg13g2_mux2_1 _7040_ (.A0(net534),
    .A1(net1036),
    .S(net910),
    .X(_0364_));
 sg13g2_a21oi_1 _7041_ (.A1(\vgademo.plane_du[0] ),
    .A2(_2728_),
    .Y(_3082_),
    .B1(net211));
 sg13g2_a21oi_1 _7042_ (.A1(net935),
    .A2(_2729_),
    .Y(_3083_),
    .B1(net899));
 sg13g2_nor2_1 _7043_ (.A(net212),
    .B(_3083_),
    .Y(_0365_));
 sg13g2_dfrbp_1 _7044_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net46),
    .D(_0112_),
    .Q_N(_3551_),
    .Q(\vgademo.linelfsr[0] ));
 sg13g2_dfrbp_1 _7045_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net159),
    .D(net553),
    .Q_N(_3550_),
    .Q(\vgademo.linelfsr[1] ));
 sg13g2_dfrbp_1 _7046_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net157),
    .D(net389),
    .Q_N(_3549_),
    .Q(\vgademo.linelfsr[2] ));
 sg13g2_dfrbp_1 _7047_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net155),
    .D(_0115_),
    .Q_N(_3548_),
    .Q(\vgademo.linelfsr[3] ));
 sg13g2_dfrbp_1 _7048_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net153),
    .D(net362),
    .Q_N(_3547_),
    .Q(\vgademo.linelfsr[4] ));
 sg13g2_dfrbp_1 _7049_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net151),
    .D(_0117_),
    .Q_N(_3546_),
    .Q(\vgademo.linelfsr[5] ));
 sg13g2_dfrbp_1 _7050_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net149),
    .D(net391),
    .Q_N(_3545_),
    .Q(\vgademo.linelfsr[6] ));
 sg13g2_dfrbp_1 _7051_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net147),
    .D(_0119_),
    .Q_N(_3544_),
    .Q(\vgademo.linelfsr[7] ));
 sg13g2_dfrbp_1 _7052_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net145),
    .D(net367),
    .Q_N(_3543_),
    .Q(\vgademo.linelfsr[8] ));
 sg13g2_dfrbp_1 _7053_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net143),
    .D(net377),
    .Q_N(_3542_),
    .Q(\vgademo.linelfsr[9] ));
 sg13g2_dfrbp_1 _7054_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net141),
    .D(_0122_),
    .Q_N(_3541_),
    .Q(\vgademo.linelfsr[10] ));
 sg13g2_dfrbp_1 _7055_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net139),
    .D(_0123_),
    .Q_N(_3540_),
    .Q(\vgademo.linelfsr[11] ));
 sg13g2_dfrbp_1 _7056_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(net300),
    .Q_N(_3539_),
    .Q(\vgademo.linelfsr[12] ));
 sg13g2_dfrbp_1 _7057_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1068),
    .D(net275),
    .Q_N(\vgademo.audio_songpos[0] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _7058_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1073),
    .D(_0126_),
    .Q_N(\vgademo.audio_songpos[1] ),
    .Q(_0087_));
 sg13g2_dfrbp_1 _7059_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1068),
    .D(_0127_),
    .Q_N(\vgademo.audio_songpos[2] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 _7060_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1073),
    .D(_0128_),
    .Q_N(\vgademo.audio_songpos[3] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _7061_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1068),
    .D(_0129_),
    .Q_N(\vgademo.audio_songpos[4] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _7062_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1068),
    .D(_0130_),
    .Q_N(\vgademo.audio_songpos[5] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _7063_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1073),
    .D(_0131_),
    .Q_N(\vgademo.audio_songpos[6] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 _7064_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1073),
    .D(_0132_),
    .Q_N(\vgademo.audio_songpos[7] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 _7065_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net119),
    .D(_0133_),
    .Q_N(_0024_),
    .Q(\vgademo.plane_dx[1] ));
 sg13g2_dfrbp_1 _7066_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net117),
    .D(_0134_),
    .Q_N(_0025_),
    .Q(\vgademo.plane_dx[2] ));
 sg13g2_dfrbp_1 _7067_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net115),
    .D(_0135_),
    .Q_N(_0022_),
    .Q(\vgademo.plane_dx[3] ));
 sg13g2_dfrbp_1 _7068_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net113),
    .D(_0136_),
    .Q_N(_0023_),
    .Q(\vgademo.plane_dx_div.q[3] ));
 sg13g2_dfrbp_1 _7069_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net111),
    .D(_0137_),
    .Q_N(_3538_),
    .Q(\vgademo.plane_dx_div.q[4] ));
 sg13g2_dfrbp_1 _7070_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net109),
    .D(_0138_),
    .Q_N(_3537_),
    .Q(\vgademo.plane_dx_div.q[5] ));
 sg13g2_dfrbp_1 _7071_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net107),
    .D(_0139_),
    .Q_N(_3536_),
    .Q(\vgademo.plane_dx_div.q[6] ));
 sg13g2_dfrbp_1 _7072_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net105),
    .D(_0140_),
    .Q_N(_0026_),
    .Q(\vgademo.plane_dx_div.q[7] ));
 sg13g2_dfrbp_1 _7073_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net103),
    .D(_0141_),
    .Q_N(_3535_),
    .Q(\vgademo.plane_dx_div.q[8] ));
 sg13g2_dfrbp_1 _7074_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net101),
    .D(_0142_),
    .Q_N(_3534_),
    .Q(\vgademo.plane_dx_div.q[9] ));
 sg13g2_dfrbp_1 _7075_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net99),
    .D(net169),
    .Q_N(_0085_),
    .Q(\vgademo.plane_dx_div.i[0] ));
 sg13g2_dfrbp_1 _7076_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net97),
    .D(_0144_),
    .Q_N(_3533_),
    .Q(\vgademo.plane_dx_div.i[1] ));
 sg13g2_dfrbp_1 _7077_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net95),
    .D(net544),
    .Q_N(_3532_),
    .Q(\vgademo.plane_dx_div.i[2] ));
 sg13g2_dfrbp_1 _7078_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net47),
    .D(_0146_),
    .Q_N(_3552_),
    .Q(\vgademo.plane_dx_div.i[3] ));
 sg13g2_dfrbp_1 _7079_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1070),
    .D(\vgademo.soundtrack.sigma_delta_accum_[0] ),
    .Q_N(_3553_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[0] ));
 sg13g2_dfrbp_1 _7080_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1070),
    .D(\vgademo.soundtrack.sigma_delta_accum_[1] ),
    .Q_N(_3554_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[1] ));
 sg13g2_dfrbp_1 _7081_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1070),
    .D(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .Q_N(_3555_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[2] ));
 sg13g2_dfrbp_1 _7082_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1069),
    .D(net537),
    .Q_N(_3556_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[3] ));
 sg13g2_dfrbp_1 _7083_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1069),
    .D(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .Q_N(_3557_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[4] ));
 sg13g2_dfrbp_1 _7084_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1069),
    .D(net533),
    .Q_N(_3558_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[5] ));
 sg13g2_dfrbp_1 _7085_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1069),
    .D(\vgademo.soundtrack.sigma_delta_accum_[6] ),
    .Q_N(_3559_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[6] ));
 sg13g2_dfrbp_1 _7086_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1069),
    .D(net528),
    .Q_N(_3560_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[7] ));
 sg13g2_dfrbp_1 _7087_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1069),
    .D(net517),
    .Q_N(_3561_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[8] ));
 sg13g2_dfrbp_1 _7088_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1067),
    .D(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .Q_N(_3562_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[9] ));
 sg13g2_dfrbp_1 _7089_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1067),
    .D(net505),
    .Q_N(_3563_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[10] ));
 sg13g2_dfrbp_1 _7090_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1067),
    .D(net495),
    .Q_N(_3564_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[11] ));
 sg13g2_dfrbp_1 _7091_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1067),
    .D(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .Q_N(_3565_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[12] ));
 sg13g2_dfrbp_1 _7092_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1067),
    .D(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .Q_N(_3566_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[13] ));
 sg13g2_dfrbp_1 _7093_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1067),
    .D(\vgademo.soundtrack.sigma_delta_accum_[14] ),
    .Q_N(_3567_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[14] ));
 sg13g2_dfrbp_1 _7094_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1067),
    .D(\vgademo.soundtrack.sigma_delta_accum_[15] ),
    .Q_N(_3531_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[15] ));
 sg13g2_dfrbp_1 _7095_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1072),
    .D(_0147_),
    .Q_N(_0058_),
    .Q(\vgademo.audio_beat_out[0] ));
 sg13g2_dfrbp_1 _7096_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1072),
    .D(net375),
    .Q_N(_0059_),
    .Q(\vgademo.audio_beat_out[1] ));
 sg13g2_dfrbp_1 _7097_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1072),
    .D(_0149_),
    .Q_N(_0062_),
    .Q(\vgademo.audio_beat_out[2] ));
 sg13g2_dfrbp_1 _7098_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1072),
    .D(_0150_),
    .Q_N(_0057_),
    .Q(\vgademo.audio_beat_out[3] ));
 sg13g2_dfrbp_1 _7099_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1072),
    .D(_0151_),
    .Q_N(_0055_),
    .Q(\vgademo.audio_beat_out[4] ));
 sg13g2_dfrbp_1 _7100_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1084),
    .D(_0152_),
    .Q_N(_3530_),
    .Q(\vgademo.soundtrack.tri_osc_i[0] ));
 sg13g2_dfrbp_1 _7101_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1081),
    .D(_0153_),
    .Q_N(_3529_),
    .Q(\vgademo.soundtrack.tri_osc_i[1] ));
 sg13g2_dfrbp_1 _7102_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1071),
    .D(net452),
    .Q_N(_3528_),
    .Q(\vgademo.soundtrack.tri_osc_i[2] ));
 sg13g2_dfrbp_1 _7103_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1072),
    .D(_0155_),
    .Q_N(_3527_),
    .Q(\vgademo.soundtrack.tri_osc_i[3] ));
 sg13g2_dfrbp_1 _7104_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1071),
    .D(_0156_),
    .Q_N(_3526_),
    .Q(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_dfrbp_1 _7105_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1070),
    .D(_0157_),
    .Q_N(_3525_),
    .Q(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_dfrbp_1 _7106_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1070),
    .D(_0158_),
    .Q_N(_3524_),
    .Q(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_dfrbp_1 _7107_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1070),
    .D(_0159_),
    .Q_N(_3523_),
    .Q(\vgademo.soundtrack.tri_osc_i[7] ));
 sg13g2_dfrbp_1 _7108_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1070),
    .D(_0160_),
    .Q_N(_3522_),
    .Q(\vgademo.soundtrack.tri_osc_i[8] ));
 sg13g2_dfrbp_1 _7109_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net89),
    .D(net198),
    .Q_N(_3521_),
    .Q(audio));
 sg13g2_dfrbp_1 _7110_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1082),
    .D(net179),
    .Q_N(\vgademo.soundtrack.tick_div_[0] ),
    .Q(\vgademo.soundtrack.tick_div[0] ));
 sg13g2_dfrbp_1 _7111_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1082),
    .D(net498),
    .Q_N(_3520_),
    .Q(\vgademo.soundtrack.tick_div[1] ));
 sg13g2_dfrbp_1 _7112_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1082),
    .D(net265),
    .Q_N(_3519_),
    .Q(\vgademo.soundtrack.tick_div[2] ));
 sg13g2_dfrbp_1 _7113_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1082),
    .D(net244),
    .Q_N(_3518_),
    .Q(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_dfrbp_1 _7114_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1080),
    .D(net210),
    .Q_N(_3517_),
    .Q(\vgademo.soundtrack.tick_div[4] ));
 sg13g2_dfrbp_1 _7115_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1085),
    .D(net263),
    .Q_N(_3516_),
    .Q(\vgademo.soundtrack.tick_div[5] ));
 sg13g2_dfrbp_1 _7116_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1084),
    .D(net205),
    .Q_N(_3515_),
    .Q(\vgademo.soundtrack.tick_div[6] ));
 sg13g2_dfrbp_1 _7117_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(net231),
    .Q_N(_3514_),
    .Q(\vgademo.soundtrack.tick_div[7] ));
 sg13g2_dfrbp_1 _7118_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1080),
    .D(net171),
    .Q_N(\vgademo.soundtrack.noise_lfsr[0] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 _7119_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1080),
    .D(net167),
    .Q_N(\vgademo.soundtrack.noise_lfsr[1] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 _7120_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1080),
    .D(net183),
    .Q_N(\vgademo.soundtrack.noise_lfsr[2] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 _7121_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1081),
    .D(net229),
    .Q_N(\vgademo.soundtrack.noise_lfsr[3] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 _7122_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1081),
    .D(net234),
    .Q_N(_0040_),
    .Q(\vgademo.soundtrack.noise_lfsr[4] ));
 sg13g2_dfrbp_1 _7123_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1081),
    .D(net175),
    .Q_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 _7124_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1081),
    .D(net277),
    .Q_N(_0084_),
    .Q(\vgademo.soundtrack.noise_lfsr[6] ));
 sg13g2_dfrbp_1 _7125_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1081),
    .D(net177),
    .Q_N(\vgademo.soundtrack.noise_lfsr[7] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 _7126_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1081),
    .D(net324),
    .Q_N(_0083_),
    .Q(\vgademo.soundtrack.noise_lfsr[8] ));
 sg13g2_dfrbp_1 _7127_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1080),
    .D(net186),
    .Q_N(_3513_),
    .Q(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_dfrbp_1 _7128_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1070),
    .D(net181),
    .Q_N(\vgademo.soundtrack.noise_lfsr[10] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _7129_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1080),
    .D(net173),
    .Q_N(\vgademo.soundtrack.noise_lfsr[11] ),
    .Q(_0101_));
 sg13g2_dfrbp_1 _7130_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1080),
    .D(net202),
    .Q_N(\vgademo.soundtrack.noise_lfsr[12] ),
    .Q(_0102_));
 sg13g2_dfrbp_1 _7131_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1080),
    .D(net242),
    .Q_N(_0082_),
    .Q(\vgademo.soundtrack.noise_lfsr[13] ));
 sg13g2_dfrbp_1 _7132_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1083),
    .D(net333),
    .Q_N(_3512_),
    .Q(\vgademo.soundtrack.noise_lfsr[14] ));
 sg13g2_dfrbp_1 _7133_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1084),
    .D(net200),
    .Q_N(\vgademo.audio_snare_frames[0] ),
    .Q(_0103_));
 sg13g2_dfrbp_1 _7134_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1084),
    .D(net259),
    .Q_N(\vgademo.audio_snare_frames[1] ),
    .Q(_0104_));
 sg13g2_dfrbp_1 _7135_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1072),
    .D(net246),
    .Q_N(\vgademo.audio_snare_frames[2] ),
    .Q(_0105_));
 sg13g2_dfrbp_1 _7136_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1072),
    .D(net193),
    .Q_N(\vgademo.audio_snare_frames[3] ),
    .Q(_0106_));
 sg13g2_dfrbp_1 _7137_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net62),
    .D(_0189_),
    .Q_N(_3511_),
    .Q(\vgademo.soundtrack.pulse_osc_p[0] ));
 sg13g2_dfrbp_1 _7138_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net61),
    .D(net191),
    .Q_N(_0042_),
    .Q(\vgademo.soundtrack.pulse_osc_p[1] ));
 sg13g2_dfrbp_1 _7139_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net60),
    .D(_0191_),
    .Q_N(_3510_),
    .Q(\vgademo.soundtrack.pulse_osc_p[2] ));
 sg13g2_dfrbp_1 _7140_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net59),
    .D(net340),
    .Q_N(_3509_),
    .Q(\vgademo.soundtrack.pulse_osc_p[3] ));
 sg13g2_dfrbp_1 _7141_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net58),
    .D(_0193_),
    .Q_N(_3508_),
    .Q(\vgademo.soundtrack.pulse_osc_p[4] ));
 sg13g2_dfrbp_1 _7142_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net57),
    .D(_0194_),
    .Q_N(_3507_),
    .Q(\vgademo.soundtrack.pulse_osc_p[5] ));
 sg13g2_dfrbp_1 _7143_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net56),
    .D(_0195_),
    .Q_N(_3506_),
    .Q(\vgademo.soundtrack.pulse_osc_p[6] ));
 sg13g2_dfrbp_1 _7144_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net55),
    .D(_0196_),
    .Q_N(_3505_),
    .Q(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_dfrbp_1 _7145_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net54),
    .D(net225),
    .Q_N(_3504_),
    .Q(\vgademo.soundtrack.pulse_osc_p[8] ));
 sg13g2_dfrbp_1 _7146_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net53),
    .D(_0198_),
    .Q_N(_3503_),
    .Q(\vgademo.soundtrack.pulse_osc_p[9] ));
 sg13g2_dfrbp_1 _7147_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net52),
    .D(net196),
    .Q_N(_3502_),
    .Q(\vgademo.soundtrack.pulse_osc_p[10] ));
 sg13g2_dfrbp_1 _7148_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net51),
    .D(_0200_),
    .Q_N(_3501_),
    .Q(\vgademo.soundtrack.pulse_osc_p[11] ));
 sg13g2_dfrbp_1 _7149_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net50),
    .D(_0201_),
    .Q_N(_3500_),
    .Q(\vgademo.soundtrack.pulse_osc_p[12] ));
 sg13g2_dfrbp_1 _7150_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net49),
    .D(net252),
    .Q_N(_3499_),
    .Q(\vgademo.soundtrack.pulse_osc_p[13] ));
 sg13g2_dfrbp_1 _7151_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1084),
    .D(_0203_),
    .Q_N(_3498_),
    .Q(\vgademo.audio_kick_frames[0] ));
 sg13g2_dfrbp_1 _7152_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1085),
    .D(net455),
    .Q_N(_0068_),
    .Q(\vgademo.audio_kick_frames[1] ));
 sg13g2_dfrbp_1 _7153_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1085),
    .D(net387),
    .Q_N(_0060_),
    .Q(\vgademo.audio_kick_frames[2] ));
 sg13g2_dfrbp_1 _7154_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1068),
    .D(_0206_),
    .Q_N(\vgademo.soundtrack.pulse_vol[0] ),
    .Q(_0107_));
 sg13g2_dfrbp_1 _7155_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1069),
    .D(_0207_),
    .Q_N(\vgademo.soundtrack.pulse_vol[1] ),
    .Q(_0108_));
 sg13g2_dfrbp_1 _7156_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1068),
    .D(_0208_),
    .Q_N(\vgademo.soundtrack.pulse_vol[2] ),
    .Q(_0109_));
 sg13g2_dfrbp_1 _7157_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1068),
    .D(net221),
    .Q_N(\vgademo.soundtrack.pulse_vol[3] ),
    .Q(_0110_));
 sg13g2_dfrbp_1 _7158_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1082),
    .D(net165),
    .Q_N(\vgademo.soundtrack.sample_div_[0] ),
    .Q(\vgademo.soundtrack.sample_div[0] ));
 sg13g2_dfrbp_1 _7159_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1086),
    .D(net254),
    .Q_N(_3568_),
    .Q(\vgademo.soundtrack.sample_div[1] ));
 sg13g2_dfrbp_1 _7160_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1082),
    .D(net477),
    .Q_N(_3569_),
    .Q(\vgademo.soundtrack.sample_div[2] ));
 sg13g2_dfrbp_1 _7161_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1082),
    .D(net240),
    .Q_N(_3570_),
    .Q(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_dfrbp_1 _7162_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1082),
    .D(net227),
    .Q_N(_3571_),
    .Q(\vgademo.soundtrack.sample_div[4] ));
 sg13g2_dfrbp_1 _7163_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1091),
    .D(\vgademo.soundtrack.sample_div_[5] ),
    .Q_N(_3572_),
    .Q(\vgademo.soundtrack.sample_div[5] ));
 sg13g2_dfrbp_1 _7164_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1083),
    .D(\vgademo.soundtrack.sample_div_[6] ),
    .Q_N(_3573_),
    .Q(\vgademo.soundtrack.sample_div[6] ));
 sg13g2_dfrbp_1 _7165_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1083),
    .D(net248),
    .Q_N(_3574_),
    .Q(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_dfrbp_1 _7166_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1083),
    .D(net219),
    .Q_N(_3575_),
    .Q(\vgademo.soundtrack.sample_div[8] ));
 sg13g2_dfrbp_1 _7167_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1083),
    .D(\vgademo.soundtrack.sample_div_[9] ),
    .Q_N(_3497_),
    .Q(\vgademo.soundtrack.sample_div[9] ));
 sg13g2_dfrbp_1 _7168_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net38),
    .D(net207),
    .Q_N(_3496_),
    .Q(\vgademo.soundtrack.tri_osc_p[0] ));
 sg13g2_dfrbp_1 _7169_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net37),
    .D(net349),
    .Q_N(_3495_),
    .Q(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_dfrbp_1 _7170_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net36),
    .D(_0212_),
    .Q_N(_3494_),
    .Q(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_dfrbp_1 _7171_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net35),
    .D(net398),
    .Q_N(_3493_),
    .Q(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_dfrbp_1 _7172_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net34),
    .D(_0214_),
    .Q_N(_3492_),
    .Q(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_dfrbp_1 _7173_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net33),
    .D(_0215_),
    .Q_N(_3491_),
    .Q(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_dfrbp_1 _7174_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net32),
    .D(net418),
    .Q_N(_3490_),
    .Q(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_dfrbp_1 _7175_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net31),
    .D(_0217_),
    .Q_N(_3489_),
    .Q(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_dfrbp_1 _7176_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net30),
    .D(_0218_),
    .Q_N(_3488_),
    .Q(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_dfrbp_1 _7177_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net29),
    .D(net373),
    .Q_N(_0041_),
    .Q(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_dfrbp_1 _7178_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net28),
    .D(net282),
    .Q_N(_3487_),
    .Q(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_dfrbp_1 _7179_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net27),
    .D(net359),
    .Q_N(_3486_),
    .Q(\vgademo.soundtrack.tri_osc_p[11] ));
 sg13g2_dfrbp_1 _7180_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net26),
    .D(_0222_),
    .Q_N(_3485_),
    .Q(\vgademo.soundtrack.tri_osc_p[12] ));
 sg13g2_dfrbp_1 _7181_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net25),
    .D(net306),
    .Q_N(_3484_),
    .Q(\vgademo.soundtrack.tri_osc_p[13] ));
 sg13g2_dfrbp_1 _7182_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net24),
    .D(net355),
    .Q_N(_3483_),
    .Q(\vgademo.soundtrack.tri_osc_p[14] ));
 sg13g2_dfrbp_1 _7183_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net23),
    .D(net432),
    .Q_N(_3482_),
    .Q(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_dfrbp_1 _7184_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net22),
    .D(_0226_),
    .Q_N(_3481_),
    .Q(\vgademo.plane_dx_div.d[16] ));
 sg13g2_dfrbp_1 _7185_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net21),
    .D(_0227_),
    .Q_N(_0070_),
    .Q(\vgademo.plane_dx_div.d[17] ));
 sg13g2_dfrbp_1 _7186_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net20),
    .D(_0228_),
    .Q_N(_0073_),
    .Q(\vgademo.plane_dx_div.d[18] ));
 sg13g2_dfrbp_1 _7187_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net19),
    .D(_0229_),
    .Q_N(_0076_),
    .Q(\vgademo.plane_dx_div.d[19] ));
 sg13g2_dfrbp_1 _7188_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net18),
    .D(_0230_),
    .Q_N(_0079_),
    .Q(\vgademo.plane_dx_div.d[20] ));
 sg13g2_dfrbp_1 _7189_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net17),
    .D(_0231_),
    .Q_N(_0081_),
    .Q(\vgademo.plane_dx_div.d[21] ));
 sg13g2_dfrbp_1 _7190_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net16),
    .D(_0232_),
    .Q_N(_0013_),
    .Q(\vgademo.plane_dx_div.d[22] ));
 sg13g2_dfrbp_1 _7191_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net15),
    .D(_0233_),
    .Q_N(_0017_),
    .Q(\vgademo.plane_dx_div.d[23] ));
 sg13g2_dfrbp_1 _7192_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net91),
    .D(_0234_),
    .Q_N(_0020_),
    .Q(\vgademo.plane_dx_div.d[24] ));
 sg13g2_dfrbp_1 _7193_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net92),
    .D(_0012_),
    .Q_N(_3576_),
    .Q(\vgademo.vsync ));
 sg13g2_dfrbp_1 _7194_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net93),
    .D(_0011_),
    .Q_N(_3577_),
    .Q(hsync));
 sg13g2_dfrbp_1 _7195_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1078),
    .D(_0000_),
    .Q_N(_3578_),
    .Q(\vgademo.h_count[0] ));
 sg13g2_dfrbp_1 _7196_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1067),
    .D(_0002_),
    .Q_N(_3579_),
    .Q(\vgademo.h_count[1] ));
 sg13g2_dfrbp_1 _7197_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1068),
    .D(_0003_),
    .Q_N(_0033_),
    .Q(\vgademo.h_count[2] ));
 sg13g2_dfrbp_1 _7198_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1075),
    .D(_0004_),
    .Q_N(_0034_),
    .Q(\vgademo.h_count[3] ));
 sg13g2_dfrbp_1 _7199_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1075),
    .D(_0005_),
    .Q_N(_0044_),
    .Q(\vgademo.h_count[4] ));
 sg13g2_dfrbp_1 _7200_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1075),
    .D(_0006_),
    .Q_N(_0035_),
    .Q(\vgademo.h_count[5] ));
 sg13g2_dfrbp_1 _7201_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1075),
    .D(_0007_),
    .Q_N(_0036_),
    .Q(\vgademo.h_count[6] ));
 sg13g2_dfrbp_1 _7202_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1075),
    .D(_0008_),
    .Q_N(_0037_),
    .Q(\vgademo.h_count[7] ));
 sg13g2_dfrbp_1 _7203_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1075),
    .D(net582),
    .Q_N(_0038_),
    .Q(\vgademo.h_count[8] ));
 sg13g2_dfrbp_1 _7204_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1075),
    .D(net236),
    .Q_N(_0039_),
    .Q(\vgademo.h_count[9] ));
 sg13g2_dfrbp_1 _7205_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(_0001_),
    .Q_N(_0061_),
    .Q(\vgademo.h_count[10] ));
 sg13g2_dfrbp_1 _7206_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1078),
    .D(_0235_),
    .Q_N(_0064_),
    .Q(\vgademo.a_scrolly[3] ));
 sg13g2_dfrbp_1 _7207_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net1077),
    .D(_0236_),
    .Q_N(_0069_),
    .Q(\vgademo.a_scrolly[4] ));
 sg13g2_dfrbp_1 _7208_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1078),
    .D(net501),
    .Q_N(_0056_),
    .Q(\vgademo.a_scrolly[5] ));
 sg13g2_dfrbp_1 _7209_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1076),
    .D(_0238_),
    .Q_N(_0075_),
    .Q(\vgademo.a_scrolly[6] ));
 sg13g2_dfrbp_1 _7210_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(net530),
    .Q_N(_0078_),
    .Q(\vgademo.a_scrolly[7] ));
 sg13g2_dfrbp_1 _7211_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1076),
    .D(net319),
    .Q_N(_0080_),
    .Q(\vgademo.a_scrolly[8] ));
 sg13g2_dfrbp_1 _7212_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1077),
    .D(_0241_),
    .Q_N(_0065_),
    .Q(\vgademo.a_scrolly[9] ));
 sg13g2_dfrbp_1 _7213_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1077),
    .D(net444),
    .Q_N(_0015_),
    .Q(\vgademo.a_scrolly[10] ));
 sg13g2_dfrbp_1 _7214_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net1077),
    .D(_0243_),
    .Q_N(_0019_),
    .Q(\vgademo.a_scrolly[11] ));
 sg13g2_dfrbp_1 _7215_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1077),
    .D(_0244_),
    .Q_N(_0067_),
    .Q(\vgademo.a_scrolly[12] ));
 sg13g2_dfrbp_1 _7216_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net1077),
    .D(net569),
    .Q_N(_0066_),
    .Q(\vgademo.a_scrolly[13] ));
 sg13g2_dfrbp_1 _7217_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1078),
    .D(_0246_),
    .Q_N(_3480_),
    .Q(\vgademo.bayer_j[0] ));
 sg13g2_dfrbp_1 _7218_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1079),
    .D(_0247_),
    .Q_N(_0072_),
    .Q(\vgademo.bayer_j[1] ));
 sg13g2_dfrbp_1 _7219_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1092),
    .D(net471),
    .Q_N(_0071_),
    .Q(\vgademo.v_count[2] ));
 sg13g2_dfrbp_1 _7220_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1092),
    .D(net474),
    .Q_N(_0074_),
    .Q(\vgademo.v_count[3] ));
 sg13g2_dfrbp_1 _7221_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1092),
    .D(net303),
    .Q_N(_0077_),
    .Q(\vgademo.v_count[4] ));
 sg13g2_dfrbp_1 _7222_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1091),
    .D(_0251_),
    .Q_N(_0063_),
    .Q(\vgademo.v_count[5] ));
 sg13g2_dfrbp_1 _7223_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1091),
    .D(net562),
    .Q_N(_0016_),
    .Q(\vgademo.v_count[6] ));
 sg13g2_dfrbp_1 _7224_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1078),
    .D(net288),
    .Q_N(_0014_),
    .Q(\vgademo.v_count[7] ));
 sg13g2_dfrbp_1 _7225_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1078),
    .D(net524),
    .Q_N(_0018_),
    .Q(\vgademo.v_count[8] ));
 sg13g2_dfrbp_1 _7226_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1078),
    .D(net439),
    .Q_N(_0021_),
    .Q(\vgademo.v_count[9] ));
 sg13g2_dfrbp_1 _7227_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net163),
    .D(_0256_),
    .Q_N(_3479_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7228_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net162),
    .D(_0257_),
    .Q_N(_3478_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7229_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1088),
    .D(net238),
    .Q_N(_3477_),
    .Q(\vgademo.a_cos[0] ));
 sg13g2_dfrbp_1 _7230_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1088),
    .D(_0259_),
    .Q_N(_3476_),
    .Q(\vgademo.a_cos[1] ));
 sg13g2_dfrbp_1 _7231_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1089),
    .D(_0260_),
    .Q_N(_3475_),
    .Q(\vgademo.a_cos[2] ));
 sg13g2_dfrbp_1 _7232_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1089),
    .D(_0261_),
    .Q_N(_3474_),
    .Q(\vgademo.a_cos[3] ));
 sg13g2_dfrbp_1 _7233_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1089),
    .D(_0262_),
    .Q_N(_3473_),
    .Q(\vgademo.a_cos[4] ));
 sg13g2_dfrbp_1 _7234_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1090),
    .D(_0263_),
    .Q_N(_3472_),
    .Q(\vgademo.a_cos[5] ));
 sg13g2_dfrbp_1 _7235_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1089),
    .D(_0264_),
    .Q_N(_3471_),
    .Q(\vgademo.a_cos[6] ));
 sg13g2_dfrbp_1 _7236_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1090),
    .D(_0265_),
    .Q_N(_3470_),
    .Q(\vgademo.a_cos[7] ));
 sg13g2_dfrbp_1 _7237_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1086),
    .D(_0266_),
    .Q_N(_3469_),
    .Q(\vgademo.a_cos[8] ));
 sg13g2_dfrbp_1 _7238_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(_0267_),
    .Q_N(_3468_),
    .Q(\vgademo.a_cos[9] ));
 sg13g2_dfrbp_1 _7239_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1085),
    .D(_0268_),
    .Q_N(_3467_),
    .Q(\vgademo.a_cos[10] ));
 sg13g2_dfrbp_1 _7240_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1085),
    .D(_0269_),
    .Q_N(_3466_),
    .Q(\vgademo.a_cos[11] ));
 sg13g2_dfrbp_1 _7241_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1086),
    .D(_0270_),
    .Q_N(_3465_),
    .Q(\vgademo.a_cos[12] ));
 sg13g2_dfrbp_1 _7242_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1088),
    .D(_0271_),
    .Q_N(\vgademo.a_cos[13] ),
    .Q(_0111_));
 sg13g2_dfrbp_1 _7243_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1088),
    .D(_0272_),
    .Q_N(_3464_),
    .Q(\vgademo.a_cos[14] ));
 sg13g2_dfrbp_1 _7244_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1088),
    .D(_0273_),
    .Q_N(_3463_),
    .Q(\vgademo.a_sin[0] ));
 sg13g2_dfrbp_1 _7245_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1088),
    .D(net297),
    .Q_N(_3462_),
    .Q(\vgademo.a_sin[1] ));
 sg13g2_dfrbp_1 _7246_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1086),
    .D(_0275_),
    .Q_N(_3461_),
    .Q(\vgademo.a_sin[2] ));
 sg13g2_dfrbp_1 _7247_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1086),
    .D(_0276_),
    .Q_N(_3460_),
    .Q(\vgademo.a_sin[3] ));
 sg13g2_dfrbp_1 _7248_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(_0277_),
    .Q_N(_3459_),
    .Q(\vgademo.a_sin[4] ));
 sg13g2_dfrbp_1 _7249_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1086),
    .D(_0278_),
    .Q_N(_3458_),
    .Q(\vgademo.a_sin[5] ));
 sg13g2_dfrbp_1 _7250_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1086),
    .D(_0279_),
    .Q_N(_3457_),
    .Q(\vgademo.a_sin[6] ));
 sg13g2_dfrbp_1 _7251_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1088),
    .D(_0280_),
    .Q_N(_3456_),
    .Q(\vgademo.a_sin[7] ));
 sg13g2_dfrbp_1 _7252_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1089),
    .D(net575),
    .Q_N(_3455_),
    .Q(\vgademo.a_sin[8] ));
 sg13g2_dfrbp_1 _7253_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1089),
    .D(_0282_),
    .Q_N(_3454_),
    .Q(\vgademo.a_sin[9] ));
 sg13g2_dfrbp_1 _7254_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1089),
    .D(_0283_),
    .Q_N(_3453_),
    .Q(\vgademo.a_sin[10] ));
 sg13g2_dfrbp_1 _7255_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1090),
    .D(_0284_),
    .Q_N(_3452_),
    .Q(\vgademo.a_sin[11] ));
 sg13g2_dfrbp_1 _7256_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1089),
    .D(_0285_),
    .Q_N(_3451_),
    .Q(\vgademo.a_sin[12] ));
 sg13g2_dfrbp_1 _7257_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1090),
    .D(_0286_),
    .Q_N(_3450_),
    .Q(\vgademo.a_sin[13] ));
 sg13g2_dfrbp_1 _7258_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1088),
    .D(net503),
    .Q_N(_3449_),
    .Q(\vgademo.a_sin[14] ));
 sg13g2_dfrbp_1 _7259_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net160),
    .D(_0288_),
    .Q_N(_3448_),
    .Q(\vgademo.scanline_audio_sample[0] ));
 sg13g2_dfrbp_1 _7260_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net158),
    .D(_0289_),
    .Q_N(_3447_),
    .Q(\vgademo.scanline_audio_sample[1] ));
 sg13g2_dfrbp_1 _7261_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net156),
    .D(_0290_),
    .Q_N(_3446_),
    .Q(\vgademo.scanline_audio_sample[2] ));
 sg13g2_dfrbp_1 _7262_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net154),
    .D(_0291_),
    .Q_N(_3445_),
    .Q(\vgademo.scanline_audio_sample[3] ));
 sg13g2_dfrbp_1 _7263_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net152),
    .D(_0292_),
    .Q_N(_3444_),
    .Q(\vgademo.scanline_audio_sample[4] ));
 sg13g2_dfrbp_1 _7264_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net150),
    .D(_0293_),
    .Q_N(_0043_),
    .Q(\vgademo.scanline_audio_sample[5] ));
 sg13g2_dfrbp_1 _7265_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net148),
    .D(_0294_),
    .Q_N(_3443_),
    .Q(\vgademo.scanline_audio_sample[6] ));
 sg13g2_dfrbp_1 _7266_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net146),
    .D(net294),
    .Q_N(_3442_),
    .Q(\vgademo.b_cos[0] ));
 sg13g2_dfrbp_1 _7267_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net144),
    .D(_0296_),
    .Q_N(_3441_),
    .Q(\vgademo.b_cos[1] ));
 sg13g2_dfrbp_1 _7268_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net142),
    .D(_0297_),
    .Q_N(_3440_),
    .Q(\vgademo.b_cos[2] ));
 sg13g2_dfrbp_1 _7269_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net140),
    .D(net326),
    .Q_N(_3439_),
    .Q(\vgademo.b_cos[3] ));
 sg13g2_dfrbp_1 _7270_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net138),
    .D(net403),
    .Q_N(_3438_),
    .Q(\vgademo.b_cos[4] ));
 sg13g2_dfrbp_1 _7271_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net136),
    .D(_0300_),
    .Q_N(_3437_),
    .Q(\vgademo.b_cos[5] ));
 sg13g2_dfrbp_1 _7272_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net135),
    .D(_0301_),
    .Q_N(_3436_),
    .Q(\vgademo.b_cos[6] ));
 sg13g2_dfrbp_1 _7273_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net134),
    .D(net488),
    .Q_N(_3435_),
    .Q(\vgademo.b_cos[7] ));
 sg13g2_dfrbp_1 _7274_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net133),
    .D(net467),
    .Q_N(_3434_),
    .Q(\vgademo.b_cos[8] ));
 sg13g2_dfrbp_1 _7275_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net132),
    .D(_0304_),
    .Q_N(_3433_),
    .Q(\vgademo.b_cos[9] ));
 sg13g2_dfrbp_1 _7276_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net131),
    .D(_0305_),
    .Q_N(_3432_),
    .Q(\vgademo.b_cos[10] ));
 sg13g2_dfrbp_1 _7277_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net130),
    .D(_0306_),
    .Q_N(_3431_),
    .Q(\vgademo.b_cos[11] ));
 sg13g2_dfrbp_1 _7278_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net129),
    .D(net337),
    .Q_N(_3430_),
    .Q(\vgademo.plane_dx_div.r[16] ));
 sg13g2_dfrbp_1 _7279_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net128),
    .D(_0308_),
    .Q_N(_3429_),
    .Q(\vgademo.plane_dx_div.r[17] ));
 sg13g2_dfrbp_1 _7280_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net127),
    .D(net328),
    .Q_N(_3428_),
    .Q(\vgademo.plane_dx_div.r[18] ));
 sg13g2_dfrbp_1 _7281_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net126),
    .D(_0310_),
    .Q_N(_3427_),
    .Q(\vgademo.plane_dx_div.r[19] ));
 sg13g2_dfrbp_1 _7282_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net125),
    .D(_0311_),
    .Q_N(_3426_),
    .Q(\vgademo.plane_dx_div.r[20] ));
 sg13g2_dfrbp_1 _7283_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net124),
    .D(_0312_),
    .Q_N(_3425_),
    .Q(\vgademo.plane_dx_div.r[21] ));
 sg13g2_dfrbp_1 _7284_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net123),
    .D(net322),
    .Q_N(_3424_),
    .Q(\vgademo.plane_dx_div.r[22] ));
 sg13g2_dfrbp_1 _7285_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net122),
    .D(_0314_),
    .Q_N(_3423_),
    .Q(\vgademo.plane_dx_div.r[23] ));
 sg13g2_dfrbp_1 _7286_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net121),
    .D(net316),
    .Q_N(_3422_),
    .Q(\vgademo.plane_dx_div.r[24] ));
 sg13g2_dfrbp_1 _7287_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net120),
    .D(_0316_),
    .Q_N(\vgademo.plane_dx[0] ),
    .Q(\vgademo.plane_dx_div.r[25] ));
 sg13g2_dfrbp_1 _7288_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net118),
    .D(_0317_),
    .Q_N(_3421_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7289_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net116),
    .D(_0318_),
    .Q_N(_3420_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7290_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net114),
    .D(_0319_),
    .Q_N(_3419_),
    .Q(\vgademo.b_sin[0] ));
 sg13g2_dfrbp_1 _7291_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net112),
    .D(net357),
    .Q_N(_3418_),
    .Q(\vgademo.b_sin[1] ));
 sg13g2_dfrbp_1 _7292_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net110),
    .D(net343),
    .Q_N(_3417_),
    .Q(\vgademo.b_sin[2] ));
 sg13g2_dfrbp_1 _7293_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net108),
    .D(net416),
    .Q_N(_3416_),
    .Q(\vgademo.b_sin[3] ));
 sg13g2_dfrbp_1 _7294_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net106),
    .D(_0323_),
    .Q_N(_3415_),
    .Q(\vgademo.b_sin[4] ));
 sg13g2_dfrbp_1 _7295_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net104),
    .D(net261),
    .Q_N(_3414_),
    .Q(\vgademo.b_sin[5] ));
 sg13g2_dfrbp_1 _7296_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net102),
    .D(_0325_),
    .Q_N(_3413_),
    .Q(\vgademo.b_sin[6] ));
 sg13g2_dfrbp_1 _7297_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net100),
    .D(_0326_),
    .Q_N(_3412_),
    .Q(\vgademo.b_sin[7] ));
 sg13g2_dfrbp_1 _7298_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net98),
    .D(_0327_),
    .Q_N(_3411_),
    .Q(\vgademo.b_sin[8] ));
 sg13g2_dfrbp_1 _7299_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net96),
    .D(net383),
    .Q_N(_3410_),
    .Q(\vgademo.b_sin[9] ));
 sg13g2_dfrbp_1 _7300_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net94),
    .D(_0329_),
    .Q_N(_3409_),
    .Q(\vgademo.b_sin[10] ));
 sg13g2_dfrbp_1 _7301_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net90),
    .D(_0330_),
    .Q_N(_3408_),
    .Q(\vgademo.b_sin[11] ));
 sg13g2_dfrbp_1 _7302_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net88),
    .D(net284),
    .Q_N(_3407_),
    .Q(\vgademo.plane_u[1] ));
 sg13g2_dfrbp_1 _7303_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net87),
    .D(_0332_),
    .Q_N(_3406_),
    .Q(\vgademo.plane_u[2] ));
 sg13g2_dfrbp_1 _7304_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net86),
    .D(_0333_),
    .Q_N(_3405_),
    .Q(\vgademo.plane_u[3] ));
 sg13g2_dfrbp_1 _7305_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net85),
    .D(_0334_),
    .Q_N(_3404_),
    .Q(\vgademo.plane_u[4] ));
 sg13g2_dfrbp_1 _7306_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net84),
    .D(_0335_),
    .Q_N(_3403_),
    .Q(\vgademo.plane_u[5] ));
 sg13g2_dfrbp_1 _7307_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net83),
    .D(_0336_),
    .Q_N(_3402_),
    .Q(\vgademo.plane_u[6] ));
 sg13g2_dfrbp_1 _7308_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net82),
    .D(_0337_),
    .Q_N(_3401_),
    .Q(\vgademo.plane_u[7] ));
 sg13g2_dfrbp_1 _7309_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net81),
    .D(_0338_),
    .Q_N(_3400_),
    .Q(\vgademo.plane_u[8] ));
 sg13g2_dfrbp_1 _7310_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net80),
    .D(_0339_),
    .Q_N(_3399_),
    .Q(\vgademo.plane_u[9] ));
 sg13g2_dfrbp_1 _7311_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net79),
    .D(net410),
    .Q_N(_3398_),
    .Q(\vgademo.plane_u[10] ));
 sg13g2_dfrbp_1 _7312_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net78),
    .D(net279),
    .Q_N(_0027_),
    .Q(\vgademo.plane_u[11] ));
 sg13g2_dfrbp_1 _7313_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net77),
    .D(_0342_),
    .Q_N(_0028_),
    .Q(\vgademo.plane_u[12] ));
 sg13g2_dfrbp_1 _7314_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net76),
    .D(net435),
    .Q_N(_0048_),
    .Q(\vgademo.plane_u[13] ));
 sg13g2_dfrbp_1 _7315_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net75),
    .D(_0344_),
    .Q_N(_0029_),
    .Q(\vgademo.plane_u[14] ));
 sg13g2_dfrbp_1 _7316_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net74),
    .D(net493),
    .Q_N(_0047_),
    .Q(\vgademo.plane_u[15] ));
 sg13g2_dfrbp_1 _7317_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net73),
    .D(_0346_),
    .Q_N(_0030_),
    .Q(\vgademo.plane_u[16] ));
 sg13g2_dfrbp_1 _7318_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net72),
    .D(_0347_),
    .Q_N(_0046_),
    .Q(\vgademo.plane_u[17] ));
 sg13g2_dfrbp_1 _7319_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net71),
    .D(_0348_),
    .Q_N(_0031_),
    .Q(\vgademo.plane_u[18] ));
 sg13g2_dfrbp_1 _7320_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net70),
    .D(_0349_),
    .Q_N(_0045_),
    .Q(\vgademo.plane_u[19] ));
 sg13g2_dfrbp_1 _7321_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net69),
    .D(_0350_),
    .Q_N(_0032_),
    .Q(\vgademo.plane_u[20] ));
 sg13g2_dfrbp_1 _7322_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net68),
    .D(net400),
    .Q_N(_3397_),
    .Q(\vgademo.plane_u[21] ));
 sg13g2_dfrbp_1 _7323_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net67),
    .D(_0352_),
    .Q_N(_3396_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7324_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net66),
    .D(_0353_),
    .Q_N(_3395_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7325_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net65),
    .D(net291),
    .Q_N(_3394_),
    .Q(\vgademo.plane_du[0] ));
 sg13g2_dfrbp_1 _7326_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net64),
    .D(net311),
    .Q_N(_3393_),
    .Q(\vgademo.plane_du[1] ));
 sg13g2_dfrbp_1 _7327_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net63),
    .D(net484),
    .Q_N(_3392_),
    .Q(\vgademo.plane_du[2] ));
 sg13g2_dfrbp_1 _7328_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net48),
    .D(_0357_),
    .Q_N(_0050_),
    .Q(\vgademo.plane_du[3] ));
 sg13g2_dfrbp_1 _7329_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net45),
    .D(net521),
    .Q_N(_0049_),
    .Q(\vgademo.plane_du[4] ));
 sg13g2_dfrbp_1 _7330_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net44),
    .D(_0359_),
    .Q_N(_0051_),
    .Q(\vgademo.plane_du[5] ));
 sg13g2_dfrbp_1 _7331_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net43),
    .D(_0360_),
    .Q_N(_0052_),
    .Q(\vgademo.plane_du[6] ));
 sg13g2_dfrbp_1 _7332_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net42),
    .D(net412),
    .Q_N(_0053_),
    .Q(\vgademo.plane_du[7] ));
 sg13g2_dfrbp_1 _7333_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net41),
    .D(net564),
    .Q_N(_0054_),
    .Q(\vgademo.plane_du[8] ));
 sg13g2_dfrbp_1 _7334_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net40),
    .D(_0363_),
    .Q_N(_3391_),
    .Q(\vgademo.plane_du[9] ));
 sg13g2_dfrbp_1 _7335_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net39),
    .D(_0364_),
    .Q_N(_3390_),
    .Q(\vgademo.plane_du[10] ));
 sg13g2_dfrbp_1 _7336_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net161),
    .D(net213),
    .Q_N(_3389_),
    .Q(\vgademo.plane_u[0] ));
 sg13g2_tiehi _7190__16 (.L_HI(net16));
 sg13g2_tiehi _7189__17 (.L_HI(net17));
 sg13g2_tiehi _7188__18 (.L_HI(net18));
 sg13g2_tiehi _7187__19 (.L_HI(net19));
 sg13g2_tiehi _7186__20 (.L_HI(net20));
 sg13g2_tiehi _7185__21 (.L_HI(net21));
 sg13g2_tiehi _7184__22 (.L_HI(net22));
 sg13g2_tiehi _7183__23 (.L_HI(net23));
 sg13g2_tiehi _7182__24 (.L_HI(net24));
 sg13g2_tiehi _7181__25 (.L_HI(net25));
 sg13g2_tiehi _7180__26 (.L_HI(net26));
 sg13g2_tiehi _7179__27 (.L_HI(net27));
 sg13g2_tiehi _7178__28 (.L_HI(net28));
 sg13g2_tiehi _7177__29 (.L_HI(net29));
 sg13g2_tiehi _7176__30 (.L_HI(net30));
 sg13g2_tiehi _7175__31 (.L_HI(net31));
 sg13g2_tiehi _7174__32 (.L_HI(net32));
 sg13g2_tiehi _7173__33 (.L_HI(net33));
 sg13g2_tiehi _7172__34 (.L_HI(net34));
 sg13g2_tiehi _7171__35 (.L_HI(net35));
 sg13g2_tiehi _7170__36 (.L_HI(net36));
 sg13g2_tiehi _7169__37 (.L_HI(net37));
 sg13g2_tiehi _7168__38 (.L_HI(net38));
 sg13g2_tiehi _7335__39 (.L_HI(net39));
 sg13g2_tiehi _7334__40 (.L_HI(net40));
 sg13g2_tiehi _7333__41 (.L_HI(net41));
 sg13g2_tiehi _7332__42 (.L_HI(net42));
 sg13g2_tiehi _7331__43 (.L_HI(net43));
 sg13g2_tiehi _7330__44 (.L_HI(net44));
 sg13g2_tiehi _7329__45 (.L_HI(net45));
 sg13g2_tiehi _7044__46 (.L_HI(net46));
 sg13g2_tiehi _7078__47 (.L_HI(net47));
 sg13g2_tiehi _7328__48 (.L_HI(net48));
 sg13g2_tiehi _7150__49 (.L_HI(net49));
 sg13g2_tiehi _7149__50 (.L_HI(net50));
 sg13g2_tiehi _7148__51 (.L_HI(net51));
 sg13g2_tiehi _7147__52 (.L_HI(net52));
 sg13g2_tiehi _7146__53 (.L_HI(net53));
 sg13g2_tiehi _7145__54 (.L_HI(net54));
 sg13g2_tiehi _7144__55 (.L_HI(net55));
 sg13g2_tiehi _7143__56 (.L_HI(net56));
 sg13g2_tiehi _7142__57 (.L_HI(net57));
 sg13g2_tiehi _7141__58 (.L_HI(net58));
 sg13g2_tiehi _7140__59 (.L_HI(net59));
 sg13g2_tiehi _7139__60 (.L_HI(net60));
 sg13g2_tiehi _7138__61 (.L_HI(net61));
 sg13g2_tiehi _7137__62 (.L_HI(net62));
 sg13g2_tiehi _7327__63 (.L_HI(net63));
 sg13g2_tiehi _7326__64 (.L_HI(net64));
 sg13g2_tiehi _7325__65 (.L_HI(net65));
 sg13g2_tiehi _7324__66 (.L_HI(net66));
 sg13g2_tiehi _7323__67 (.L_HI(net67));
 sg13g2_tiehi _7322__68 (.L_HI(net68));
 sg13g2_tiehi _7321__69 (.L_HI(net69));
 sg13g2_tiehi _7320__70 (.L_HI(net70));
 sg13g2_tiehi _7319__71 (.L_HI(net71));
 sg13g2_tiehi _7318__72 (.L_HI(net72));
 sg13g2_tiehi _7317__73 (.L_HI(net73));
 sg13g2_tiehi _7316__74 (.L_HI(net74));
 sg13g2_tiehi _7315__75 (.L_HI(net75));
 sg13g2_tiehi _7314__76 (.L_HI(net76));
 sg13g2_tiehi _7313__77 (.L_HI(net77));
 sg13g2_tiehi _7312__78 (.L_HI(net78));
 sg13g2_tiehi _7311__79 (.L_HI(net79));
 sg13g2_tiehi _7310__80 (.L_HI(net80));
 sg13g2_tiehi _7309__81 (.L_HI(net81));
 sg13g2_tiehi _7308__82 (.L_HI(net82));
 sg13g2_tiehi _7307__83 (.L_HI(net83));
 sg13g2_tiehi _7306__84 (.L_HI(net84));
 sg13g2_tiehi _7305__85 (.L_HI(net85));
 sg13g2_tiehi _7304__86 (.L_HI(net86));
 sg13g2_tiehi _7303__87 (.L_HI(net87));
 sg13g2_tiehi _7302__88 (.L_HI(net88));
 sg13g2_tiehi _7109__89 (.L_HI(net89));
 sg13g2_tiehi _7301__90 (.L_HI(net90));
 sg13g2_tiehi _7192__91 (.L_HI(net91));
 sg13g2_tiehi _7193__92 (.L_HI(net92));
 sg13g2_tiehi _7194__93 (.L_HI(net93));
 sg13g2_tiehi _7300__94 (.L_HI(net94));
 sg13g2_tiehi _7077__95 (.L_HI(net95));
 sg13g2_tiehi _7299__96 (.L_HI(net96));
 sg13g2_tiehi _7076__97 (.L_HI(net97));
 sg13g2_tiehi _7298__98 (.L_HI(net98));
 sg13g2_tiehi _7075__99 (.L_HI(net99));
 sg13g2_tiehi _7297__100 (.L_HI(net100));
 sg13g2_tiehi _7074__101 (.L_HI(net101));
 sg13g2_tiehi _7296__102 (.L_HI(net102));
 sg13g2_tiehi _7073__103 (.L_HI(net103));
 sg13g2_tiehi _7295__104 (.L_HI(net104));
 sg13g2_tiehi _7072__105 (.L_HI(net105));
 sg13g2_tiehi _7294__106 (.L_HI(net106));
 sg13g2_tiehi _7071__107 (.L_HI(net107));
 sg13g2_tiehi _7293__108 (.L_HI(net108));
 sg13g2_tiehi _7070__109 (.L_HI(net109));
 sg13g2_tiehi _7292__110 (.L_HI(net110));
 sg13g2_tiehi _7069__111 (.L_HI(net111));
 sg13g2_tiehi _7291__112 (.L_HI(net112));
 sg13g2_tiehi _7068__113 (.L_HI(net113));
 sg13g2_tiehi _7290__114 (.L_HI(net114));
 sg13g2_tiehi _7067__115 (.L_HI(net115));
 sg13g2_tiehi _7289__116 (.L_HI(net116));
 sg13g2_tiehi _7066__117 (.L_HI(net117));
 sg13g2_tiehi _7288__118 (.L_HI(net118));
 sg13g2_tiehi _7065__119 (.L_HI(net119));
 sg13g2_tiehi _7287__120 (.L_HI(net120));
 sg13g2_tiehi _7286__121 (.L_HI(net121));
 sg13g2_tiehi _7285__122 (.L_HI(net122));
 sg13g2_tiehi _7284__123 (.L_HI(net123));
 sg13g2_tiehi _7283__124 (.L_HI(net124));
 sg13g2_tiehi _7282__125 (.L_HI(net125));
 sg13g2_tiehi _7281__126 (.L_HI(net126));
 sg13g2_tiehi _7280__127 (.L_HI(net127));
 sg13g2_tiehi _7279__128 (.L_HI(net128));
 sg13g2_tiehi _7278__129 (.L_HI(net129));
 sg13g2_tiehi _7277__130 (.L_HI(net130));
 sg13g2_tiehi _7276__131 (.L_HI(net131));
 sg13g2_tiehi _7275__132 (.L_HI(net132));
 sg13g2_tiehi _7274__133 (.L_HI(net133));
 sg13g2_tiehi _7273__134 (.L_HI(net134));
 sg13g2_tiehi _7272__135 (.L_HI(net135));
 sg13g2_tiehi _7271__136 (.L_HI(net136));
 sg13g2_tiehi _7056__137 (.L_HI(net137));
 sg13g2_tiehi _7270__138 (.L_HI(net138));
 sg13g2_tiehi _7055__139 (.L_HI(net139));
 sg13g2_tiehi _7269__140 (.L_HI(net140));
 sg13g2_tiehi _7054__141 (.L_HI(net141));
 sg13g2_tiehi _7268__142 (.L_HI(net142));
 sg13g2_tiehi _7053__143 (.L_HI(net143));
 sg13g2_tiehi _7267__144 (.L_HI(net144));
 sg13g2_tiehi _7052__145 (.L_HI(net145));
 sg13g2_tiehi _7266__146 (.L_HI(net146));
 sg13g2_tiehi _7051__147 (.L_HI(net147));
 sg13g2_tiehi _7265__148 (.L_HI(net148));
 sg13g2_tiehi _7050__149 (.L_HI(net149));
 sg13g2_tiehi _7264__150 (.L_HI(net150));
 sg13g2_tiehi _7049__151 (.L_HI(net151));
 sg13g2_tiehi _7263__152 (.L_HI(net152));
 sg13g2_tiehi _7048__153 (.L_HI(net153));
 sg13g2_tiehi _7262__154 (.L_HI(net154));
 sg13g2_tiehi _7047__155 (.L_HI(net155));
 sg13g2_tiehi _7261__156 (.L_HI(net156));
 sg13g2_tiehi _7046__157 (.L_HI(net157));
 sg13g2_tiehi _7260__158 (.L_HI(net158));
 sg13g2_tiehi _7045__159 (.L_HI(net159));
 sg13g2_tiehi _7259__160 (.L_HI(net160));
 sg13g2_tiehi _7336__161 (.L_HI(net161));
 sg13g2_tiehi _7228__162 (.L_HI(net162));
 sg13g2_tiehi _7227__163 (.L_HI(net163));
 sg13g2_tiehi tt_um_a1k0n_demo_164 (.L_HI(net164));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_a1k0n_demo_2 (.L_LO(net2));
 sg13g2_tielo tt_um_a1k0n_demo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_a1k0n_demo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_a1k0n_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_a1k0n_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_a1k0n_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_a1k0n_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_a1k0n_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_a1k0n_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_a1k0n_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_a1k0n_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_a1k0n_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_a1k0n_demo_14 (.L_LO(net14));
 sg13g2_tiehi _7191__15 (.L_HI(net15));
 sg13g2_buf_2 _7501_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_1 _7502_ (.A(\vgademo.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7503_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout832 (.A(_1779_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_1779_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_1779_),
    .X(net834));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(_1757_));
 sg13g2_buf_1 fanout836 (.A(_1757_),
    .X(net836));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(net838));
 sg13g2_buf_2 fanout838 (.A(_2348_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_1465_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_1464_),
    .X(net841));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(net843));
 sg13g2_buf_2 fanout843 (.A(_1428_),
    .X(net843));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(_1427_));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_1426_),
    .X(net846));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(_1425_));
 sg13g2_buf_2 fanout848 (.A(_1425_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_2483_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_1461_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_1411_),
    .X(net854));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(_1342_));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(_1449_));
 sg13g2_buf_2 fanout857 (.A(_1448_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_1437_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_1408_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_1407_),
    .X(net860));
 sg13g2_buf_4 fanout861 (.X(net861),
    .A(_1341_));
 sg13g2_buf_2 fanout862 (.A(_1445_),
    .X(net862));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(_1434_));
 sg13g2_buf_2 fanout864 (.A(_1434_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_1433_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_1322_),
    .X(net866));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(_0682_));
 sg13g2_buf_1 fanout868 (.A(_0682_),
    .X(net868));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(_0626_));
 sg13g2_buf_1 fanout870 (.A(_0626_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(net873),
    .X(net871));
 sg13g2_buf_1 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_1 fanout873 (.A(net876),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net876),
    .X(net874));
 sg13g2_buf_4 fanout875 (.X(net875),
    .A(net876));
 sg13g2_buf_4 fanout876 (.X(net876),
    .A(_1321_));
 sg13g2_buf_2 fanout877 (.A(_0622_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(net879),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_1274_),
    .X(net879));
 sg13g2_buf_4 fanout880 (.X(net880),
    .A(_0810_));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_1 fanout882 (.A(net885),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(net885),
    .X(net883));
 sg13g2_buf_1 fanout884 (.A(net885),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_0809_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_0577_),
    .X(net886));
 sg13g2_buf_1 fanout887 (.A(_0577_),
    .X(net887));
 sg13g2_buf_4 fanout888 (.X(net888),
    .A(net889));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(_0576_));
 sg13g2_buf_4 fanout890 (.X(net890),
    .A(_1191_));
 sg13g2_buf_2 fanout891 (.A(_0594_),
    .X(net891));
 sg13g2_buf_1 fanout892 (.A(_0594_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_0594_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(net897),
    .X(net895));
 sg13g2_buf_1 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_2727_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(net901),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net901),
    .X(net899));
 sg13g2_buf_1 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_2727_),
    .X(net902));
 sg13g2_buf_4 fanout903 (.X(net903),
    .A(net904));
 sg13g2_buf_2 fanout904 (.A(_2421_),
    .X(net904));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(net908));
 sg13g2_buf_2 fanout906 (.A(net908),
    .X(net906));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(net908));
 sg13g2_buf_2 fanout908 (.A(_0585_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(net911),
    .X(net909));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(net911));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_4 fanout912 (.X(net912),
    .A(_2418_));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(net914));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(_0648_));
 sg13g2_buf_2 fanout915 (.A(net916),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_0647_),
    .X(net916));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(net921));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(net921),
    .X(net919));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(net921));
 sg13g2_buf_4 fanout921 (.X(net921),
    .A(_0591_));
 sg13g2_buf_2 fanout922 (.A(net925),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(_0590_));
 sg13g2_buf_2 fanout926 (.A(net928),
    .X(net926));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(net928));
 sg13g2_buf_2 fanout928 (.A(_0584_),
    .X(net928));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(_0583_));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_4 fanout931 (.X(net931),
    .A(_0582_));
 sg13g2_buf_2 fanout932 (.A(net934),
    .X(net932));
 sg13g2_buf_1 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(net936),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_0582_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(net938),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(_0581_));
 sg13g2_buf_2 fanout942 (.A(_1042_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_1042_),
    .X(net943));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(_0646_));
 sg13g2_buf_2 fanout945 (.A(net947),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(net947),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_0645_),
    .X(net947));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(_3212_));
 sg13g2_buf_1 fanout949 (.A(_3212_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_0694_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_2229_),
    .X(net951));
 sg13g2_buf_1 fanout952 (.A(_2229_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_2171_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_3290_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_3126_),
    .X(net956));
 sg13g2_buf_4 fanout957 (.X(net957),
    .A(_3118_));
 sg13g2_buf_4 fanout958 (.X(net958),
    .A(_3106_));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(_3105_));
 sg13g2_buf_2 fanout960 (.A(_3103_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_3103_),
    .X(net961));
 sg13g2_buf_4 fanout962 (.X(net962),
    .A(net584));
 sg13g2_buf_4 fanout963 (.X(net963),
    .A(\vgademo.plane_du[8] ));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(net965));
 sg13g2_buf_2 fanout965 (.A(net535),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(net969),
    .X(net967));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(net969));
 sg13g2_buf_2 fanout969 (.A(net590),
    .X(net969));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(\vgademo.b_cos[10] ));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(net572));
 sg13g2_buf_4 fanout972 (.X(net972),
    .A(\vgademo.a_sin[14] ));
 sg13g2_buf_4 fanout973 (.X(net973),
    .A(\vgademo.v_count[9] ));
 sg13g2_buf_4 fanout974 (.X(net974),
    .A(\vgademo.v_count[7] ));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(net561));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(\vgademo.v_count[5] ));
 sg13g2_buf_2 fanout977 (.A(net468),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(\vgademo.v_count[4] ),
    .X(net978));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(net573));
 sg13g2_buf_2 fanout980 (.A(\vgademo.a_scrolly[13] ),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(net982),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(\vgademo.a_scrolly[12] ),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(net551),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(net986),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(net986),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(\vgademo.a_scrolly[10] ),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(net989),
    .X(net987));
 sg13g2_buf_1 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(\vgademo.a_scrolly[9] ));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(net991));
 sg13g2_buf_4 fanout991 (.X(net991),
    .A(\vgademo.a_scrolly[8] ));
 sg13g2_buf_4 fanout992 (.X(net992),
    .A(net993));
 sg13g2_buf_4 fanout993 (.X(net993),
    .A(\vgademo.a_scrolly[7] ));
 sg13g2_buf_2 fanout994 (.A(net529),
    .X(net994));
 sg13g2_buf_4 fanout995 (.X(net995),
    .A(net996));
 sg13g2_buf_4 fanout996 (.X(net996),
    .A(\vgademo.a_scrolly[6] ));
 sg13g2_buf_4 fanout997 (.X(net997),
    .A(net1000));
 sg13g2_buf_1 fanout998 (.A(net1000),
    .X(net998));
 sg13g2_buf_4 fanout999 (.X(net999),
    .A(net1000));
 sg13g2_buf_2 fanout1000 (.A(net500),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_4 fanout1002 (.X(net1002),
    .A(net531));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(net1004));
 sg13g2_buf_4 fanout1004 (.X(net1004),
    .A(net1005));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(net554));
 sg13g2_buf_2 fanout1006 (.A(_0061_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(\vgademo.h_count[8] ),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(\vgademo.h_count[6] ),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(net507),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(\vgademo.h_count[3] ),
    .X(net1010));
 sg13g2_buf_1 fanout1011 (.A(\vgademo.h_count[3] ),
    .X(net1011));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(net1013));
 sg13g2_buf_2 fanout1013 (.A(\vgademo.h_count[2] ),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(\vgademo.h_count[1] ),
    .X(net1015));
 sg13g2_buf_4 fanout1016 (.X(net1016),
    .A(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_buf_4 fanout1017 (.X(net1017),
    .A(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_buf_2 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_1 fanout1019 (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_1 fanout1022 (.A(net1023),
    .X(net1022));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(\vgademo.audio_snare_frames[3] ));
 sg13g2_buf_2 fanout1024 (.A(net1026),
    .X(net1024));
 sg13g2_buf_1 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(net1027),
    .X(net1026));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(\vgademo.audio_snare_frames[2] ));
 sg13g2_buf_2 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(\vgademo.audio_snare_frames[1] ),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1034),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net1035),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(\vgademo.audio_snare_frames[0] ),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(net545),
    .X(net1036));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(\vgademo.plane_dx_div.q[8] ));
 sg13g2_buf_2 fanout1038 (.A(net250),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(net563),
    .X(net1039));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(net411));
 sg13g2_buf_2 fanout1041 (.A(net514),
    .X(net1041));
 sg13g2_buf_4 fanout1042 (.X(net1042),
    .A(net249));
 sg13g2_buf_2 fanout1043 (.A(\vgademo.plane_dx_div.q[4] ),
    .X(net1043));
 sg13g2_buf_4 fanout1044 (.X(net1044),
    .A(net520));
 sg13g2_buf_2 fanout1045 (.A(\vgademo.audio_songpos[7] ),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(net1047),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(net1048),
    .X(net1047));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(\vgademo.audio_songpos[5] ));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(net1051));
 sg13g2_buf_2 fanout1051 (.A(\vgademo.audio_songpos[4] ),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(net1054));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(\vgademo.audio_songpos[3] ));
 sg13g2_buf_2 fanout1055 (.A(net1057),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(\vgademo.audio_songpos[2] ),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(\vgademo.audio_songpos[1] ),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(\vgademo.audio_songpos[0] ),
    .X(net1061));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(\vgademo.audio_songpos[0] ));
 sg13g2_buf_2 fanout1063 (.A(\vgademo.linelfsr[1] ),
    .X(net1063));
 sg13g2_buf_1 fanout1064 (.A(\vgademo.linelfsr[1] ),
    .X(net1064));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(\vgademo.linelfsr[0] ));
 sg13g2_buf_2 fanout1066 (.A(net464),
    .X(net1066));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(net1074));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(net1069));
 sg13g2_buf_4 fanout1069 (.X(net1069),
    .A(net1074));
 sg13g2_buf_8 fanout1070 (.A(net1074),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(net1074),
    .X(net1071));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1073));
 sg13g2_buf_2 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(net1092));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(net1076));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_4 fanout1077 (.X(net1077),
    .A(net1079));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(net1079));
 sg13g2_buf_2 fanout1079 (.A(net1092),
    .X(net1079));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1087));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(net1087));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net1083));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(net1087));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(net1085));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(net1086));
 sg13g2_buf_4 fanout1086 (.X(net1086),
    .A(net1087));
 sg13g2_buf_2 fanout1087 (.A(net1091),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(net1090));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(net1090));
 sg13g2_buf_4 fanout1090 (.X(net1090),
    .A(net1091));
 sg13g2_buf_4 fanout1091 (.X(net1091),
    .A(net1092));
 sg13g2_buf_4 fanout1092 (.X(net1092),
    .A(rst_n));
 sg13g2_tielo tt_um_a1k0n_demo_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_1_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_55_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_2_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_4_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_51_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_52_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_54_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_49_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_50_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_14_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_17_clk));
 sg13g2_inv_8 clkload31 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_44_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_34_clk));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_40_clk));
 sg13g2_inv_1 clkload37 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload39 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload41 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload42 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload43 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload44 (.A(clknet_leaf_36_clk));
 sg13g2_inv_2 clkload45 (.A(clknet_leaf_37_clk));
 sg13g2_inv_1 clkload46 (.A(clknet_leaf_27_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vgademo.soundtrack.sample_div_[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold2 (.A(\vgademo.soundtrack.noise_lfsr[2] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0171_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0085_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0143_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold6 (.A(\vgademo.soundtrack.noise_lfsr[1] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0170_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold8 (.A(\vgademo.soundtrack.noise_lfsr[12] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0181_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0084_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0175_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0083_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0177_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold14 (.A(\vgademo.soundtrack.tick_div_[0] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0162_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold16 (.A(\vgademo.soundtrack.noise_lfsr[11] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0180_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold18 (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0172_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0090_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold21 (.A(\vgademo.soundtrack.noise_lfsr[10] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0179_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold23 (.A(\vgademo.plane_dx_div.q[3] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0652_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0089_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold26 (.A(\vgademo.soundtrack.pulse_osc_p[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0190_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0106_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0188_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold30 (.A(\vgademo.soundtrack.pulse_osc_p[10] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0933_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0199_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold33 (.A(audio),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0161_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0103_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0185_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0082_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0182_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold39 (.A(\vgademo.soundtrack.tick_div[6] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0781_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0168_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vgademo.soundtrack.tri_osc_p[0] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0210_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0108_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold45 (.A(\vgademo.soundtrack.tick_div[4] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0166_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold47 (.A(\vgademo.plane_u[0] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold48 (.A(_3082_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0365_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vgademo.soundtrack.sigma_delta_accum[0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold51 (.A(\vgademo.a_sin[0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold52 (.A(\vgademo.plane_dx_div.q[7] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0656_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vgademo.soundtrack.sample_div[8] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold55 (.A(\vgademo.soundtrack.sample_div_[8] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0110_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0209_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0107_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0109_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold60 (.A(\vgademo.soundtrack.pulse_osc_p[8] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0197_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold62 (.A(\vgademo.soundtrack.sample_div[4] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold63 (.A(\vgademo.soundtrack.sample_div_[4] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0097_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0173_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold66 (.A(\vgademo.soundtrack.tick_div[7] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0169_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0111_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold69 (.A(\vgademo.soundtrack.noise_lfsr[4] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0174_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0039_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0010_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold73 (.A(\vgademo.a_cos[0] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0258_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold75 (.A(\vgademo.soundtrack.sample_div[3] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold76 (.A(\vgademo.soundtrack.sample_div_[3] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold77 (.A(\vgademo.soundtrack.noise_lfsr[13] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0183_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold79 (.A(\vgademo.soundtrack.tick_div[3] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0165_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0105_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0187_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold83 (.A(\vgademo.soundtrack.sample_div[7] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold84 (.A(\vgademo.soundtrack.sample_div_[7] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold85 (.A(\vgademo.plane_dx_div.q[4] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold86 (.A(\vgademo.plane_dx_div.q[8] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold87 (.A(\vgademo.soundtrack.pulse_osc_p[13] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0202_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold89 (.A(\vgademo.soundtrack.sample_div[0] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold90 (.A(\vgademo.soundtrack.sample_div_[1] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold91 (.A(\vgademo.plane_u[20] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold92 (.A(\vgademo.soundtrack.pulse_osc_p[9] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold93 (.A(\vgademo.soundtrack.pulse_osc_p[11] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0104_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0186_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold96 (.A(\vgademo.b_sin[5] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0324_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold98 (.A(\vgademo.soundtrack.tick_div[5] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0167_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold100 (.A(\vgademo.soundtrack.tick_div[2] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0164_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold102 (.A(\vgademo.soundtrack.sample_div[9] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vgademo.b_sin[7] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold104 (.A(\vgademo.soundtrack.sample_div[5] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0087_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold106 (.A(\vgademo.plane_dx_div.r[21] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0093_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0088_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0091_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0086_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0125_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold112 (.A(\vgademo.soundtrack.noise_lfsr[7] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0176_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold114 (.A(\vgademo.plane_u[11] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0341_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0092_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold117 (.A(\vgademo.soundtrack.tri_osc_p[10] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0220_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold119 (.A(\vgademo.plane_u[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0331_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold121 (.A(\vgademo.plane_dx_div.d[23] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold122 (.A(\vgademo.soundtrack.pulse_osc_p[0] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold123 (.A(\vgademo.v_count[7] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0253_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold125 (.A(\vgademo.plane_dx_div.d[18] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold126 (.A(\vgademo.plane_du[0] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0354_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold128 (.A(\vgademo.plane_u[4] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold129 (.A(\vgademo.b_cos[0] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0295_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold131 (.A(\vgademo.a_sin[2] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold132 (.A(\vgademo.a_sin[1] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0274_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold134 (.A(\vgademo.plane_dx_div.d[20] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold135 (.A(\vgademo.linelfsr[12] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0124_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold137 (.A(\vgademo.plane_dx_div.d[22] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold138 (.A(\vgademo.v_count[4] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0250_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold140 (.A(\vgademo.plane_u[6] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold141 (.A(\vgademo.soundtrack.tri_osc_p[13] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0223_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold143 (.A(\vgademo.plane_dx_div.d[24] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold144 (.A(\vgademo.a_cos[1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold145 (.A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold146 (.A(\vgademo.plane_du[1] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0355_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold148 (.A(\vgademo.plane_dx_div.r[20] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold149 (.A(\vgademo.soundtrack.pulse_osc_p[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold150 (.A(\vgademo.plane_u[5] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold151 (.A(\vgademo.plane_dx_div.r[24] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0315_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold153 (.A(\vgademo.scanline_audio_sample[0] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold154 (.A(\vgademo.a_scrolly[8] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0240_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold156 (.A(\vgademo.a_cos[2] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold157 (.A(\vgademo.plane_dx_div.r[22] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0313_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold159 (.A(\vgademo.soundtrack.noise_lfsr[8] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0178_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold161 (.A(\vgademo.b_cos[3] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0298_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold163 (.A(\vgademo.plane_dx_div.r[18] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0309_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0034_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold166 (.A(_3218_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold167 (.A(\vgademo.plane_u[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold168 (.A(\vgademo.soundtrack.noise_lfsr[14] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0184_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold170 (.A(\vgademo.plane_dx_div.r[19] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold171 (.A(\vgademo.linelfsr[11] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold172 (.A(\vgademo.plane_dx_div.r[16] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0307_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold174 (.A(\vgademo.plane_u[8] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold175 (.A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0192_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold177 (.A(\vgademo.a_sin[5] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold178 (.A(_2665_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0321_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold180 (.A(\vgademo.plane_u[7] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold181 (.A(\vgademo.plane_u[2] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold182 (.A(\vgademo.a_sin[4] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold183 (.A(\vgademo.scanline_audio_sample[2] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold184 (.A(\vgademo.soundtrack.tri_osc_p[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0211_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold186 (.A(\vgademo.soundtrack.pulse_osc_p[7] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold187 (.A(\vgademo.audio_beat_out[0] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold188 (.A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold189 (.A(\vgademo.plane_u[9] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold190 (.A(\vgademo.soundtrack.tri_osc_p[14] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0224_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold192 (.A(\vgademo.b_sin[1] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0320_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold194 (.A(\vgademo.soundtrack.tri_osc_p[11] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0221_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold196 (.A(\vgademo.scanline_audio_sample[5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold197 (.A(\vgademo.linelfsr[4] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0116_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold199 (.A(\vgademo.plane_dx_div.d[19] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold200 (.A(\vgademo.plane_u[16] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold201 (.A(_2972_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold202 (.A(\vgademo.linelfsr[8] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0120_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold204 (.A(\vgademo.a_cos[12] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold205 (.A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold206 (.A(\vgademo.plane_dx_div.d[21] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0041_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold208 (.A(_1010_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0219_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold210 (.A(\vgademo.audio_beat_out[1] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0148_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold212 (.A(\vgademo.linelfsr[9] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0121_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold214 (.A(\vgademo.scanline_audio_sample[1] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold215 (.A(\vgademo.b_sin[0] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold216 (.A(_2655_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold217 (.A(\vgademo.soundtrack.sigma_delta_accum[1] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold218 (.A(\vgademo.b_sin[9] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0328_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold220 (.A(\vgademo.plane_dx_div.d[17] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold221 (.A(\vgademo.audio_kick_frames[2] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0940_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0205_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold224 (.A(\vgademo.linelfsr[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0114_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold226 (.A(\vgademo.linelfsr[6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0118_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold228 (.A(\vgademo.plane_u[14] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold229 (.A(\vgademo.linelfsr[10] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold230 (.A(\vgademo.plane_dx_div.i[0] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0659_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold232 (.A(\vgademo.linelfsr[5] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold233 (.A(\vgademo.soundtrack.tri_osc_p[3] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0213_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold235 (.A(\vgademo.plane_u[21] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0351_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold237 (.A(\vgademo.soundtrack.tri_osc_p[2] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold238 (.A(\vgademo.b_cos[4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0299_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold240 (.A(\vgademo.plane_dx_div.r[23] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold241 (.A(\vgademo.linelfsr[7] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold242 (.A(\vgademo.a_sin[3] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold243 (.A(\vgademo.plane_dx_div.i[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0662_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold245 (.A(\vgademo.plane_u[10] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0340_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold247 (.A(\vgademo.plane_dx_div.q[6] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0361_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold249 (.A(\vgademo.soundtrack.tri_osc_p[5] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold250 (.A(\vgademo.b_sin[3] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold251 (.A(_2671_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0322_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold253 (.A(\vgademo.soundtrack.tri_osc_p[6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0216_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold255 (.A(\vgademo.plane_u[19] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold256 (.A(_2997_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold257 (.A(\vgademo.soundtrack.tri_osc_p[4] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold258 (.A(\vgademo.b_cos[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold259 (.A(_2434_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold260 (.A(\vgademo.plane_u[12] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold261 (.A(_2907_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold262 (.A(\vgademo.plane_u[17] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold263 (.A(\vgademo.plane_dx_div.d[16] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold264 (.A(\vgademo.plane_dx_div.r[17] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold265 (.A(\vgademo.a_sin[6] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold266 (.A(\vgademo.scanline_audio_sample[4] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold267 (.A(\vgademo.soundtrack.tri_osc_p[12] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0225_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold269 (.A(\vgademo.b_cos[1] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold270 (.A(\vgademo.plane_u[13] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0343_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold272 (.A(\vgademo.a_cos[5] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0021_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold274 (.A(_1247_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0255_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold276 (.A(\vgademo.b_sin[6] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold277 (.A(_2690_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0015_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold279 (.A(_1211_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0242_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0037_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold282 (.A(_3226_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold283 (.A(\vgademo.soundtrack.tri_osc_p[7] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0019_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold285 (.A(_1217_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold286 (.A(\vgademo.a_sin[9] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold287 (.A(\vgademo.soundtrack.tri_osc_i[2] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0154_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold289 (.A(\vgademo.soundtrack.tri_osc_p[8] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold290 (.A(\vgademo.audio_kick_frames[1] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0204_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold292 (.A(\vgademo.b_sin[4] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold293 (.A(_2677_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold294 (.A(\vgademo.a_sin[13] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold295 (.A(\vgademo.a_cos[3] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0035_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold297 (.A(_3222_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold298 (.A(\vgademo.soundtrack.sample_div[6] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold299 (.A(\vgademo.scanline_audio_sample[6] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold300 (.A(\vgademo.linelfsr[0] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0062_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold302 (.A(\vgademo.a_cos[11] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0303_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold304 (.A(\vgademo.v_count[5] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold305 (.A(\vgademo.a_cos[4] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0071_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0248_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold308 (.A(\vgademo.a_cos[14] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold309 (.A(\vgademo.v_count[3] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0249_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold311 (.A(\vgademo.soundtrack.sample_div[2] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0569_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold313 (.A(\vgademo.soundtrack.sample_div_[2] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold314 (.A(\vgademo.a_sin[12] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold315 (.A(\vgademo.audio_beat_out[4] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0674_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold317 (.A(\vgademo.b_sin[8] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold318 (.A(_2706_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold319 (.A(\vgademo.plane_du[2] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0356_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold321 (.A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold322 (.A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold323 (.A(\vgademo.a_cos[10] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0302_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0063_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold326 (.A(\vgademo.b_sin[10] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold327 (.A(\vgademo.a_sin[11] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold328 (.A(\vgademo.plane_u[15] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0345_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold330 (.A(\vgademo.soundtrack.sigma_delta_accum[11] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold331 (.A(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold332 (.A(\vgademo.soundtrack.tick_div[1] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0780_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0163_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold335 (.A(\vgademo.a_cos[6] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold336 (.A(\vgademo.a_scrolly[5] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0237_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold338 (.A(\vgademo.a_sin[14] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0287_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold340 (.A(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold341 (.A(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0033_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold343 (.A(\vgademo.h_count[4] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold344 (.A(\vgademo.soundtrack.pulse_osc_p[12] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold345 (.A(\vgademo.scanline_audio_sample[3] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold346 (.A(\vgademo.soundtrack.tri_osc_i[3] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold347 (.A(\vgademo.a_cos[9] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold348 (.A(\vgademo.soundtrack.sigma_delta_accum[12] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold349 (.A(\vgademo.plane_u[18] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold350 (.A(\vgademo.plane_dx_div.q[5] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold351 (.A(\vgademo.soundtrack.sigma_delta_accum[13] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold352 (.A(\vgademo.soundtrack.sigma_delta_accum[8] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold353 (.A(\vgademo.soundtrack.sigma_delta_accum_[8] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold354 (.A(\vgademo.audio_beat_out[3] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold355 (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0023_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0358_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0018_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold359 (.A(_1243_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0254_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0065_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold362 (.A(\vgademo.soundtrack.sigma_delta_accum[9] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold363 (.A(\vgademo.soundtrack.sigma_delta_accum[7] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold364 (.A(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold365 (.A(\vgademo.a_scrolly[7] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0239_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold367 (.A(\vgademo.a_scrolly[4] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold368 (.A(\vgademo.soundtrack.sigma_delta_accum[5] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold369 (.A(\vgademo.soundtrack.sigma_delta_accum_[5] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold370 (.A(\vgademo.plane_du[10] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold371 (.A(\vgademo.b_sin[11] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold372 (.A(\vgademo.soundtrack.sigma_delta_accum[3] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold373 (.A(\vgademo.soundtrack.sigma_delta_accum_[3] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold374 (.A(\vgademo.plane_dx[3] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0651_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold376 (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold377 (.A(\vgademo.plane_du[3] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold378 (.A(\vgademo.plane_dx_div.i[2] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0660_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0145_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold381 (.A(\vgademo.plane_dx_div.q[9] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold382 (.A(\vgademo.h_count[0] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold383 (.A(\vgademo.plane_du[5] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold384 (.A(\vgademo.soundtrack.sigma_delta_accum[14] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold385 (.A(\vgademo.a_sin[10] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold386 (.A(\vgademo.a_sin[7] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold387 (.A(\vgademo.a_scrolly[11] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold388 (.A(\vgademo.linelfsr[2] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0113_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold390 (.A(\vgademo.a_scrolly[3] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold391 (.A(\vgademo.a_cos[8] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold392 (.A(_2448_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold393 (.A(\vgademo.soundtrack.tri_osc_i[8] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold394 (.A(\vgademo.b_cos[11] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold395 (.A(\vgademo.plane_dx[1] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0650_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold397 (.A(\vgademo.v_count[6] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0252_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0026_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0362_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold401 (.A(\vgademo.soundtrack.sigma_delta_accum[6] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold402 (.A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold403 (.A(\vgademo.plane_dx[0] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0066_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0245_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold406 (.A(\vgademo.soundtrack.sigma_delta_accum[2] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold407 (.A(\vgademo.a_cos[7] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold408 (.A(\vgademo.b_cos[6] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold409 (.A(\vgademo.bayer_j[0] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold410 (.A(\vgademo.a_sin[8] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0281_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0036_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold413 (.A(_3224_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold414 (.A(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold415 (.A(\vgademo.soundtrack.sigma_delta_accum[4] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0038_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold417 (.A(_3228_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0009_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold419 (.A(\vgademo.plane_du[6] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold420 (.A(\vgademo.plane_du[9] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold421 (.A(\vgademo.a_cos[13] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold422 (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold423 (.A(\vgademo.audio_kick_frames[0] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0075_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold425 (.A(\vgademo.bayer_j[1] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold426 (.A(\vgademo.plane_dx_div.r[25] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold427 (.A(\vgademo.h_count[9] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold428 (.A(_3233_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold429 (.A(\vgademo.h_count[8] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold430 (.A(\vgademo.b_cos[1] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold431 (.A(\vgademo.audio_beat_out[3] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold432 (.A(\vgademo.a_sin[8] ),
    .X(net596));
 sg13g2_antennanp ANTENNA_1 (.A(_0594_));
 sg13g2_antennanp ANTENNA_2 (.A(_0594_));
 sg13g2_antennanp ANTENNA_3 (.A(_0594_));
 sg13g2_antennanp ANTENNA_4 (.A(_0594_));
 sg13g2_antennanp ANTENNA_5 (.A(_0594_));
 sg13g2_antennanp ANTENNA_6 (.A(_0594_));
 sg13g2_antennanp ANTENNA_7 (.A(_0594_));
 sg13g2_antennanp ANTENNA_8 (.A(_0594_));
 sg13g2_antennanp ANTENNA_9 (.A(_0594_));
 sg13g2_antennanp ANTENNA_10 (.A(_0594_));
 sg13g2_antennanp ANTENNA_11 (.A(_0594_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_decap_8 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_104 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_decap_8 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_132 ();
 sg13g2_decap_4 FILLER_9_139 ();
 sg13g2_decap_8 FILLER_9_146 ();
 sg13g2_decap_8 FILLER_9_153 ();
 sg13g2_decap_8 FILLER_9_160 ();
 sg13g2_decap_8 FILLER_9_167 ();
 sg13g2_decap_8 FILLER_9_174 ();
 sg13g2_decap_8 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_188 ();
 sg13g2_decap_8 FILLER_9_195 ();
 sg13g2_decap_8 FILLER_9_202 ();
 sg13g2_decap_8 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_230 ();
 sg13g2_decap_8 FILLER_9_237 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_265 ();
 sg13g2_decap_8 FILLER_9_272 ();
 sg13g2_decap_8 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_8 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_8 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_9_433 ();
 sg13g2_decap_8 FILLER_9_440 ();
 sg13g2_decap_8 FILLER_9_447 ();
 sg13g2_decap_8 FILLER_9_454 ();
 sg13g2_decap_8 FILLER_9_461 ();
 sg13g2_decap_8 FILLER_9_468 ();
 sg13g2_decap_8 FILLER_9_475 ();
 sg13g2_decap_8 FILLER_9_482 ();
 sg13g2_decap_8 FILLER_9_489 ();
 sg13g2_decap_8 FILLER_9_496 ();
 sg13g2_decap_8 FILLER_9_503 ();
 sg13g2_decap_8 FILLER_9_510 ();
 sg13g2_decap_8 FILLER_9_517 ();
 sg13g2_decap_8 FILLER_9_524 ();
 sg13g2_decap_8 FILLER_9_531 ();
 sg13g2_decap_8 FILLER_9_538 ();
 sg13g2_decap_8 FILLER_9_545 ();
 sg13g2_decap_8 FILLER_9_552 ();
 sg13g2_decap_8 FILLER_9_559 ();
 sg13g2_decap_8 FILLER_9_566 ();
 sg13g2_decap_8 FILLER_9_573 ();
 sg13g2_decap_8 FILLER_9_580 ();
 sg13g2_decap_8 FILLER_9_587 ();
 sg13g2_decap_8 FILLER_9_594 ();
 sg13g2_decap_8 FILLER_9_601 ();
 sg13g2_decap_8 FILLER_9_608 ();
 sg13g2_decap_8 FILLER_9_615 ();
 sg13g2_decap_8 FILLER_9_622 ();
 sg13g2_decap_8 FILLER_9_629 ();
 sg13g2_decap_8 FILLER_9_636 ();
 sg13g2_decap_8 FILLER_9_643 ();
 sg13g2_decap_8 FILLER_9_650 ();
 sg13g2_decap_8 FILLER_9_657 ();
 sg13g2_decap_8 FILLER_9_664 ();
 sg13g2_decap_8 FILLER_9_671 ();
 sg13g2_decap_8 FILLER_9_678 ();
 sg13g2_decap_8 FILLER_9_685 ();
 sg13g2_decap_8 FILLER_9_692 ();
 sg13g2_decap_8 FILLER_9_699 ();
 sg13g2_decap_8 FILLER_9_706 ();
 sg13g2_decap_8 FILLER_9_713 ();
 sg13g2_decap_8 FILLER_9_720 ();
 sg13g2_decap_8 FILLER_9_727 ();
 sg13g2_decap_8 FILLER_9_734 ();
 sg13g2_decap_8 FILLER_9_741 ();
 sg13g2_decap_8 FILLER_9_748 ();
 sg13g2_decap_8 FILLER_9_755 ();
 sg13g2_decap_8 FILLER_9_762 ();
 sg13g2_decap_8 FILLER_9_769 ();
 sg13g2_decap_8 FILLER_9_776 ();
 sg13g2_decap_8 FILLER_9_783 ();
 sg13g2_decap_8 FILLER_9_790 ();
 sg13g2_decap_8 FILLER_9_797 ();
 sg13g2_decap_8 FILLER_9_804 ();
 sg13g2_decap_8 FILLER_9_811 ();
 sg13g2_decap_8 FILLER_9_818 ();
 sg13g2_decap_8 FILLER_9_825 ();
 sg13g2_decap_8 FILLER_9_832 ();
 sg13g2_decap_8 FILLER_9_839 ();
 sg13g2_decap_8 FILLER_9_846 ();
 sg13g2_decap_8 FILLER_9_853 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_4 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_4 FILLER_10_112 ();
 sg13g2_fill_1 FILLER_10_116 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_decap_8 FILLER_10_153 ();
 sg13g2_decap_8 FILLER_10_160 ();
 sg13g2_decap_8 FILLER_10_167 ();
 sg13g2_decap_8 FILLER_10_174 ();
 sg13g2_decap_8 FILLER_10_181 ();
 sg13g2_decap_8 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_195 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_fill_2 FILLER_10_216 ();
 sg13g2_decap_4 FILLER_10_223 ();
 sg13g2_decap_4 FILLER_10_237 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_fill_1 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_fill_2 FILLER_10_300 ();
 sg13g2_fill_1 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_fill_2 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_111 ();
 sg13g2_fill_1 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_132 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_fill_2 FILLER_11_186 ();
 sg13g2_fill_1 FILLER_11_188 ();
 sg13g2_fill_2 FILLER_11_215 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_253 ();
 sg13g2_fill_2 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_decap_8 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_11_415 ();
 sg13g2_decap_8 FILLER_11_422 ();
 sg13g2_decap_8 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_11_436 ();
 sg13g2_decap_8 FILLER_11_443 ();
 sg13g2_decap_8 FILLER_11_450 ();
 sg13g2_decap_8 FILLER_11_457 ();
 sg13g2_decap_8 FILLER_11_464 ();
 sg13g2_decap_8 FILLER_11_471 ();
 sg13g2_decap_8 FILLER_11_478 ();
 sg13g2_decap_8 FILLER_11_485 ();
 sg13g2_decap_8 FILLER_11_492 ();
 sg13g2_decap_8 FILLER_11_499 ();
 sg13g2_decap_8 FILLER_11_506 ();
 sg13g2_decap_8 FILLER_11_513 ();
 sg13g2_decap_8 FILLER_11_520 ();
 sg13g2_decap_8 FILLER_11_527 ();
 sg13g2_decap_8 FILLER_11_534 ();
 sg13g2_decap_8 FILLER_11_541 ();
 sg13g2_decap_8 FILLER_11_548 ();
 sg13g2_decap_8 FILLER_11_555 ();
 sg13g2_decap_8 FILLER_11_562 ();
 sg13g2_decap_8 FILLER_11_569 ();
 sg13g2_decap_8 FILLER_11_576 ();
 sg13g2_decap_8 FILLER_11_583 ();
 sg13g2_decap_8 FILLER_11_590 ();
 sg13g2_decap_8 FILLER_11_597 ();
 sg13g2_decap_8 FILLER_11_604 ();
 sg13g2_decap_8 FILLER_11_611 ();
 sg13g2_decap_8 FILLER_11_618 ();
 sg13g2_decap_8 FILLER_11_625 ();
 sg13g2_decap_8 FILLER_11_632 ();
 sg13g2_decap_8 FILLER_11_639 ();
 sg13g2_decap_8 FILLER_11_646 ();
 sg13g2_decap_8 FILLER_11_653 ();
 sg13g2_decap_8 FILLER_11_660 ();
 sg13g2_decap_8 FILLER_11_667 ();
 sg13g2_decap_8 FILLER_11_674 ();
 sg13g2_decap_8 FILLER_11_681 ();
 sg13g2_decap_8 FILLER_11_688 ();
 sg13g2_decap_8 FILLER_11_695 ();
 sg13g2_decap_8 FILLER_11_702 ();
 sg13g2_decap_8 FILLER_11_709 ();
 sg13g2_decap_8 FILLER_11_716 ();
 sg13g2_decap_8 FILLER_11_723 ();
 sg13g2_decap_8 FILLER_11_730 ();
 sg13g2_decap_8 FILLER_11_737 ();
 sg13g2_decap_8 FILLER_11_744 ();
 sg13g2_decap_8 FILLER_11_751 ();
 sg13g2_decap_8 FILLER_11_758 ();
 sg13g2_decap_8 FILLER_11_765 ();
 sg13g2_decap_8 FILLER_11_772 ();
 sg13g2_decap_8 FILLER_11_779 ();
 sg13g2_decap_8 FILLER_11_786 ();
 sg13g2_decap_8 FILLER_11_793 ();
 sg13g2_decap_8 FILLER_11_800 ();
 sg13g2_decap_8 FILLER_11_807 ();
 sg13g2_decap_8 FILLER_11_814 ();
 sg13g2_decap_8 FILLER_11_821 ();
 sg13g2_decap_8 FILLER_11_828 ();
 sg13g2_decap_8 FILLER_11_835 ();
 sg13g2_decap_8 FILLER_11_842 ();
 sg13g2_decap_8 FILLER_11_849 ();
 sg13g2_decap_4 FILLER_11_856 ();
 sg13g2_fill_2 FILLER_11_860 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_decap_4 FILLER_12_118 ();
 sg13g2_fill_2 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_144 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_173 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_decap_8 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_194 ();
 sg13g2_decap_8 FILLER_12_201 ();
 sg13g2_fill_2 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_decap_4 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_fill_2 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_8 FILLER_12_404 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_8 FILLER_12_425 ();
 sg13g2_decap_8 FILLER_12_432 ();
 sg13g2_decap_8 FILLER_12_439 ();
 sg13g2_decap_8 FILLER_12_446 ();
 sg13g2_decap_8 FILLER_12_453 ();
 sg13g2_decap_8 FILLER_12_460 ();
 sg13g2_decap_8 FILLER_12_467 ();
 sg13g2_decap_8 FILLER_12_474 ();
 sg13g2_decap_8 FILLER_12_481 ();
 sg13g2_decap_8 FILLER_12_488 ();
 sg13g2_decap_8 FILLER_12_495 ();
 sg13g2_decap_8 FILLER_12_502 ();
 sg13g2_decap_8 FILLER_12_509 ();
 sg13g2_decap_8 FILLER_12_516 ();
 sg13g2_decap_8 FILLER_12_523 ();
 sg13g2_decap_8 FILLER_12_530 ();
 sg13g2_decap_8 FILLER_12_537 ();
 sg13g2_decap_8 FILLER_12_544 ();
 sg13g2_decap_8 FILLER_12_551 ();
 sg13g2_decap_8 FILLER_12_558 ();
 sg13g2_decap_8 FILLER_12_565 ();
 sg13g2_decap_8 FILLER_12_572 ();
 sg13g2_decap_8 FILLER_12_579 ();
 sg13g2_decap_8 FILLER_12_586 ();
 sg13g2_decap_8 FILLER_12_593 ();
 sg13g2_decap_8 FILLER_12_600 ();
 sg13g2_decap_8 FILLER_12_607 ();
 sg13g2_decap_8 FILLER_12_614 ();
 sg13g2_decap_8 FILLER_12_621 ();
 sg13g2_decap_8 FILLER_12_628 ();
 sg13g2_decap_8 FILLER_12_635 ();
 sg13g2_decap_8 FILLER_12_642 ();
 sg13g2_decap_8 FILLER_12_649 ();
 sg13g2_decap_8 FILLER_12_656 ();
 sg13g2_decap_8 FILLER_12_663 ();
 sg13g2_decap_8 FILLER_12_670 ();
 sg13g2_decap_8 FILLER_12_677 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_decap_8 FILLER_12_691 ();
 sg13g2_decap_8 FILLER_12_698 ();
 sg13g2_decap_8 FILLER_12_705 ();
 sg13g2_decap_8 FILLER_12_712 ();
 sg13g2_decap_8 FILLER_12_719 ();
 sg13g2_decap_8 FILLER_12_726 ();
 sg13g2_decap_8 FILLER_12_733 ();
 sg13g2_decap_8 FILLER_12_740 ();
 sg13g2_decap_8 FILLER_12_747 ();
 sg13g2_decap_8 FILLER_12_754 ();
 sg13g2_decap_8 FILLER_12_761 ();
 sg13g2_decap_8 FILLER_12_768 ();
 sg13g2_decap_8 FILLER_12_775 ();
 sg13g2_decap_8 FILLER_12_782 ();
 sg13g2_decap_8 FILLER_12_789 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_decap_8 FILLER_12_803 ();
 sg13g2_decap_8 FILLER_12_810 ();
 sg13g2_decap_8 FILLER_12_817 ();
 sg13g2_decap_8 FILLER_12_824 ();
 sg13g2_decap_8 FILLER_12_831 ();
 sg13g2_decap_8 FILLER_12_838 ();
 sg13g2_decap_8 FILLER_12_845 ();
 sg13g2_decap_8 FILLER_12_852 ();
 sg13g2_fill_2 FILLER_12_859 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_73 ();
 sg13g2_decap_8 FILLER_13_80 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_156 ();
 sg13g2_decap_4 FILLER_13_206 ();
 sg13g2_fill_1 FILLER_13_210 ();
 sg13g2_decap_4 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_257 ();
 sg13g2_decap_4 FILLER_13_264 ();
 sg13g2_decap_4 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_fill_2 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_fill_1 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_8 FILLER_13_404 ();
 sg13g2_decap_8 FILLER_13_411 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_8 FILLER_13_425 ();
 sg13g2_decap_8 FILLER_13_432 ();
 sg13g2_decap_8 FILLER_13_439 ();
 sg13g2_decap_8 FILLER_13_446 ();
 sg13g2_decap_8 FILLER_13_453 ();
 sg13g2_decap_8 FILLER_13_460 ();
 sg13g2_decap_8 FILLER_13_467 ();
 sg13g2_decap_8 FILLER_13_474 ();
 sg13g2_decap_8 FILLER_13_481 ();
 sg13g2_decap_8 FILLER_13_488 ();
 sg13g2_decap_8 FILLER_13_495 ();
 sg13g2_decap_8 FILLER_13_502 ();
 sg13g2_decap_8 FILLER_13_509 ();
 sg13g2_decap_8 FILLER_13_516 ();
 sg13g2_decap_8 FILLER_13_523 ();
 sg13g2_decap_8 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_537 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_decap_8 FILLER_13_551 ();
 sg13g2_decap_8 FILLER_13_558 ();
 sg13g2_decap_8 FILLER_13_565 ();
 sg13g2_decap_8 FILLER_13_572 ();
 sg13g2_decap_8 FILLER_13_579 ();
 sg13g2_decap_8 FILLER_13_586 ();
 sg13g2_decap_8 FILLER_13_593 ();
 sg13g2_decap_8 FILLER_13_600 ();
 sg13g2_decap_8 FILLER_13_607 ();
 sg13g2_decap_8 FILLER_13_614 ();
 sg13g2_decap_8 FILLER_13_621 ();
 sg13g2_decap_8 FILLER_13_628 ();
 sg13g2_decap_8 FILLER_13_635 ();
 sg13g2_decap_8 FILLER_13_642 ();
 sg13g2_decap_8 FILLER_13_649 ();
 sg13g2_decap_8 FILLER_13_656 ();
 sg13g2_decap_8 FILLER_13_663 ();
 sg13g2_decap_8 FILLER_13_670 ();
 sg13g2_decap_8 FILLER_13_677 ();
 sg13g2_decap_8 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_691 ();
 sg13g2_decap_8 FILLER_13_698 ();
 sg13g2_decap_8 FILLER_13_705 ();
 sg13g2_decap_8 FILLER_13_712 ();
 sg13g2_decap_8 FILLER_13_719 ();
 sg13g2_decap_8 FILLER_13_726 ();
 sg13g2_decap_8 FILLER_13_733 ();
 sg13g2_decap_8 FILLER_13_740 ();
 sg13g2_decap_8 FILLER_13_747 ();
 sg13g2_decap_8 FILLER_13_754 ();
 sg13g2_decap_8 FILLER_13_761 ();
 sg13g2_decap_8 FILLER_13_768 ();
 sg13g2_decap_8 FILLER_13_775 ();
 sg13g2_decap_8 FILLER_13_782 ();
 sg13g2_decap_8 FILLER_13_789 ();
 sg13g2_decap_8 FILLER_13_796 ();
 sg13g2_decap_8 FILLER_13_803 ();
 sg13g2_decap_8 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_817 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_decap_8 FILLER_13_831 ();
 sg13g2_decap_8 FILLER_13_838 ();
 sg13g2_decap_8 FILLER_13_845 ();
 sg13g2_decap_8 FILLER_13_852 ();
 sg13g2_fill_2 FILLER_13_859 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_2 FILLER_14_53 ();
 sg13g2_fill_1 FILLER_14_55 ();
 sg13g2_fill_1 FILLER_14_59 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_143 ();
 sg13g2_decap_8 FILLER_14_150 ();
 sg13g2_decap_8 FILLER_14_157 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_fill_1 FILLER_14_168 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_198 ();
 sg13g2_decap_4 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_242 ();
 sg13g2_decap_4 FILLER_14_265 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_373 ();
 sg13g2_fill_2 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_424 ();
 sg13g2_decap_8 FILLER_14_431 ();
 sg13g2_decap_8 FILLER_14_438 ();
 sg13g2_decap_8 FILLER_14_445 ();
 sg13g2_decap_8 FILLER_14_452 ();
 sg13g2_decap_8 FILLER_14_459 ();
 sg13g2_decap_8 FILLER_14_466 ();
 sg13g2_decap_8 FILLER_14_473 ();
 sg13g2_decap_8 FILLER_14_480 ();
 sg13g2_decap_8 FILLER_14_487 ();
 sg13g2_decap_8 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_501 ();
 sg13g2_decap_8 FILLER_14_508 ();
 sg13g2_decap_8 FILLER_14_515 ();
 sg13g2_decap_8 FILLER_14_522 ();
 sg13g2_decap_8 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_536 ();
 sg13g2_decap_8 FILLER_14_543 ();
 sg13g2_decap_8 FILLER_14_550 ();
 sg13g2_decap_8 FILLER_14_557 ();
 sg13g2_decap_8 FILLER_14_564 ();
 sg13g2_decap_8 FILLER_14_571 ();
 sg13g2_decap_8 FILLER_14_578 ();
 sg13g2_decap_8 FILLER_14_585 ();
 sg13g2_decap_8 FILLER_14_592 ();
 sg13g2_decap_8 FILLER_14_599 ();
 sg13g2_decap_8 FILLER_14_606 ();
 sg13g2_decap_8 FILLER_14_613 ();
 sg13g2_decap_8 FILLER_14_620 ();
 sg13g2_decap_8 FILLER_14_627 ();
 sg13g2_decap_8 FILLER_14_634 ();
 sg13g2_decap_8 FILLER_14_641 ();
 sg13g2_decap_8 FILLER_14_648 ();
 sg13g2_decap_8 FILLER_14_655 ();
 sg13g2_decap_8 FILLER_14_662 ();
 sg13g2_decap_8 FILLER_14_669 ();
 sg13g2_decap_8 FILLER_14_676 ();
 sg13g2_decap_8 FILLER_14_683 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_decap_8 FILLER_14_697 ();
 sg13g2_decap_8 FILLER_14_704 ();
 sg13g2_decap_8 FILLER_14_711 ();
 sg13g2_decap_8 FILLER_14_718 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_14_739 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_753 ();
 sg13g2_decap_8 FILLER_14_760 ();
 sg13g2_decap_8 FILLER_14_767 ();
 sg13g2_decap_8 FILLER_14_774 ();
 sg13g2_decap_8 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_788 ();
 sg13g2_decap_8 FILLER_14_795 ();
 sg13g2_decap_8 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_809 ();
 sg13g2_decap_8 FILLER_14_816 ();
 sg13g2_decap_8 FILLER_14_823 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_837 ();
 sg13g2_decap_8 FILLER_14_844 ();
 sg13g2_decap_8 FILLER_14_851 ();
 sg13g2_decap_4 FILLER_14_858 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_48 ();
 sg13g2_decap_8 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_62 ();
 sg13g2_decap_8 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_83 ();
 sg13g2_decap_8 FILLER_15_90 ();
 sg13g2_fill_1 FILLER_15_97 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_144 ();
 sg13g2_fill_1 FILLER_15_146 ();
 sg13g2_decap_4 FILLER_15_190 ();
 sg13g2_decap_8 FILLER_15_199 ();
 sg13g2_decap_4 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_210 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_fill_2 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_decap_4 FILLER_15_305 ();
 sg13g2_fill_2 FILLER_15_309 ();
 sg13g2_decap_4 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_decap_4 FILLER_15_351 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_fill_2 FILLER_15_399 ();
 sg13g2_fill_1 FILLER_15_401 ();
 sg13g2_decap_8 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_15_436 ();
 sg13g2_decap_4 FILLER_15_443 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_4 FILLER_15_487 ();
 sg13g2_fill_2 FILLER_15_491 ();
 sg13g2_decap_8 FILLER_15_502 ();
 sg13g2_fill_2 FILLER_15_509 ();
 sg13g2_decap_8 FILLER_15_519 ();
 sg13g2_decap_8 FILLER_15_526 ();
 sg13g2_decap_8 FILLER_15_533 ();
 sg13g2_decap_8 FILLER_15_540 ();
 sg13g2_decap_8 FILLER_15_547 ();
 sg13g2_decap_8 FILLER_15_554 ();
 sg13g2_decap_8 FILLER_15_561 ();
 sg13g2_decap_8 FILLER_15_568 ();
 sg13g2_decap_8 FILLER_15_575 ();
 sg13g2_decap_8 FILLER_15_582 ();
 sg13g2_decap_8 FILLER_15_589 ();
 sg13g2_decap_8 FILLER_15_596 ();
 sg13g2_decap_8 FILLER_15_603 ();
 sg13g2_decap_8 FILLER_15_610 ();
 sg13g2_decap_8 FILLER_15_617 ();
 sg13g2_decap_8 FILLER_15_624 ();
 sg13g2_decap_8 FILLER_15_631 ();
 sg13g2_decap_8 FILLER_15_638 ();
 sg13g2_decap_8 FILLER_15_645 ();
 sg13g2_decap_8 FILLER_15_652 ();
 sg13g2_decap_8 FILLER_15_659 ();
 sg13g2_decap_8 FILLER_15_666 ();
 sg13g2_decap_8 FILLER_15_673 ();
 sg13g2_decap_8 FILLER_15_680 ();
 sg13g2_decap_8 FILLER_15_687 ();
 sg13g2_decap_8 FILLER_15_694 ();
 sg13g2_decap_8 FILLER_15_701 ();
 sg13g2_decap_8 FILLER_15_708 ();
 sg13g2_decap_8 FILLER_15_715 ();
 sg13g2_decap_8 FILLER_15_722 ();
 sg13g2_decap_8 FILLER_15_729 ();
 sg13g2_decap_8 FILLER_15_736 ();
 sg13g2_decap_8 FILLER_15_743 ();
 sg13g2_decap_8 FILLER_15_750 ();
 sg13g2_decap_8 FILLER_15_757 ();
 sg13g2_decap_8 FILLER_15_764 ();
 sg13g2_decap_8 FILLER_15_771 ();
 sg13g2_decap_8 FILLER_15_778 ();
 sg13g2_decap_8 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_792 ();
 sg13g2_decap_8 FILLER_15_799 ();
 sg13g2_decap_8 FILLER_15_806 ();
 sg13g2_decap_8 FILLER_15_813 ();
 sg13g2_decap_8 FILLER_15_820 ();
 sg13g2_decap_8 FILLER_15_827 ();
 sg13g2_decap_8 FILLER_15_834 ();
 sg13g2_decap_8 FILLER_15_841 ();
 sg13g2_decap_8 FILLER_15_848 ();
 sg13g2_decap_8 FILLER_15_855 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_23 ();
 sg13g2_fill_2 FILLER_16_50 ();
 sg13g2_decap_4 FILLER_16_55 ();
 sg13g2_decap_4 FILLER_16_87 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_2 FILLER_16_98 ();
 sg13g2_fill_1 FILLER_16_100 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_120 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_159 ();
 sg13g2_fill_2 FILLER_16_207 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_decap_8 FILLER_16_262 ();
 sg13g2_fill_2 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_283 ();
 sg13g2_decap_4 FILLER_16_290 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_299 ();
 sg13g2_fill_2 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_4 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_4 FILLER_16_352 ();
 sg13g2_fill_2 FILLER_16_394 ();
 sg13g2_fill_1 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_4 FILLER_16_434 ();
 sg13g2_fill_2 FILLER_16_438 ();
 sg13g2_decap_8 FILLER_16_471 ();
 sg13g2_decap_4 FILLER_16_478 ();
 sg13g2_fill_2 FILLER_16_482 ();
 sg13g2_decap_4 FILLER_16_503 ();
 sg13g2_fill_2 FILLER_16_507 ();
 sg13g2_fill_1 FILLER_16_518 ();
 sg13g2_fill_1 FILLER_16_529 ();
 sg13g2_decap_8 FILLER_16_534 ();
 sg13g2_decap_8 FILLER_16_541 ();
 sg13g2_decap_8 FILLER_16_548 ();
 sg13g2_decap_8 FILLER_16_555 ();
 sg13g2_decap_8 FILLER_16_562 ();
 sg13g2_decap_8 FILLER_16_569 ();
 sg13g2_decap_8 FILLER_16_576 ();
 sg13g2_decap_8 FILLER_16_583 ();
 sg13g2_decap_8 FILLER_16_590 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_decap_8 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_611 ();
 sg13g2_decap_8 FILLER_16_618 ();
 sg13g2_decap_8 FILLER_16_625 ();
 sg13g2_decap_8 FILLER_16_632 ();
 sg13g2_decap_8 FILLER_16_639 ();
 sg13g2_decap_8 FILLER_16_646 ();
 sg13g2_decap_8 FILLER_16_653 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_8 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_674 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_decap_8 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_709 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_80 ();
 sg13g2_fill_1 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_180 ();
 sg13g2_decap_4 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_decap_4 FILLER_17_249 ();
 sg13g2_decap_4 FILLER_17_284 ();
 sg13g2_fill_1 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_fill_1 FILLER_17_355 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_fill_2 FILLER_17_392 ();
 sg13g2_fill_1 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_405 ();
 sg13g2_fill_2 FILLER_17_412 ();
 sg13g2_fill_1 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_547 ();
 sg13g2_decap_8 FILLER_17_554 ();
 sg13g2_decap_8 FILLER_17_561 ();
 sg13g2_decap_8 FILLER_17_568 ();
 sg13g2_decap_8 FILLER_17_575 ();
 sg13g2_decap_8 FILLER_17_582 ();
 sg13g2_decap_8 FILLER_17_589 ();
 sg13g2_decap_8 FILLER_17_596 ();
 sg13g2_decap_8 FILLER_17_603 ();
 sg13g2_decap_8 FILLER_17_610 ();
 sg13g2_decap_8 FILLER_17_617 ();
 sg13g2_decap_8 FILLER_17_624 ();
 sg13g2_decap_8 FILLER_17_631 ();
 sg13g2_decap_8 FILLER_17_638 ();
 sg13g2_decap_8 FILLER_17_645 ();
 sg13g2_decap_8 FILLER_17_652 ();
 sg13g2_decap_8 FILLER_17_659 ();
 sg13g2_decap_8 FILLER_17_666 ();
 sg13g2_decap_8 FILLER_17_673 ();
 sg13g2_decap_8 FILLER_17_680 ();
 sg13g2_decap_8 FILLER_17_687 ();
 sg13g2_decap_8 FILLER_17_694 ();
 sg13g2_decap_8 FILLER_17_701 ();
 sg13g2_decap_8 FILLER_17_708 ();
 sg13g2_decap_8 FILLER_17_715 ();
 sg13g2_decap_8 FILLER_17_722 ();
 sg13g2_decap_8 FILLER_17_729 ();
 sg13g2_decap_8 FILLER_17_736 ();
 sg13g2_decap_8 FILLER_17_743 ();
 sg13g2_decap_8 FILLER_17_750 ();
 sg13g2_decap_8 FILLER_17_757 ();
 sg13g2_decap_8 FILLER_17_764 ();
 sg13g2_decap_8 FILLER_17_771 ();
 sg13g2_decap_8 FILLER_17_778 ();
 sg13g2_decap_8 FILLER_17_785 ();
 sg13g2_decap_8 FILLER_17_792 ();
 sg13g2_decap_8 FILLER_17_799 ();
 sg13g2_decap_8 FILLER_17_806 ();
 sg13g2_decap_8 FILLER_17_813 ();
 sg13g2_decap_8 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_decap_8 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_848 ();
 sg13g2_decap_8 FILLER_17_855 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_decap_4 FILLER_18_36 ();
 sg13g2_fill_2 FILLER_18_53 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_decap_4 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_72 ();
 sg13g2_decap_8 FILLER_18_82 ();
 sg13g2_decap_8 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_96 ();
 sg13g2_decap_4 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_decap_4 FILLER_18_163 ();
 sg13g2_fill_2 FILLER_18_167 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_decap_4 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_256 ();
 sg13g2_decap_4 FILLER_18_261 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_315 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_fill_2 FILLER_18_345 ();
 sg13g2_fill_1 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_fill_2 FILLER_18_385 ();
 sg13g2_fill_1 FILLER_18_387 ();
 sg13g2_decap_4 FILLER_18_440 ();
 sg13g2_fill_1 FILLER_18_444 ();
 sg13g2_fill_2 FILLER_18_454 ();
 sg13g2_fill_1 FILLER_18_456 ();
 sg13g2_fill_2 FILLER_18_491 ();
 sg13g2_fill_1 FILLER_18_493 ();
 sg13g2_fill_2 FILLER_18_508 ();
 sg13g2_fill_1 FILLER_18_510 ();
 sg13g2_decap_8 FILLER_18_552 ();
 sg13g2_fill_2 FILLER_18_559 ();
 sg13g2_fill_1 FILLER_18_561 ();
 sg13g2_decap_8 FILLER_18_570 ();
 sg13g2_decap_8 FILLER_18_577 ();
 sg13g2_decap_8 FILLER_18_584 ();
 sg13g2_decap_8 FILLER_18_591 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_decap_8 FILLER_18_605 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_8 FILLER_18_640 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_8 FILLER_18_654 ();
 sg13g2_decap_8 FILLER_18_661 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_4 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_43 ();
 sg13g2_fill_2 FILLER_19_58 ();
 sg13g2_fill_2 FILLER_19_94 ();
 sg13g2_fill_1 FILLER_19_96 ();
 sg13g2_decap_8 FILLER_19_114 ();
 sg13g2_decap_4 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_4 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_172 ();
 sg13g2_decap_4 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_185 ();
 sg13g2_fill_2 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_206 ();
 sg13g2_decap_8 FILLER_19_213 ();
 sg13g2_decap_4 FILLER_19_220 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_4 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_289 ();
 sg13g2_fill_2 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_335 ();
 sg13g2_fill_2 FILLER_19_343 ();
 sg13g2_fill_1 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_fill_2 FILLER_19_402 ();
 sg13g2_fill_1 FILLER_19_404 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_fill_2 FILLER_19_523 ();
 sg13g2_fill_1 FILLER_19_525 ();
 sg13g2_decap_4 FILLER_19_561 ();
 sg13g2_fill_2 FILLER_19_565 ();
 sg13g2_decap_8 FILLER_19_593 ();
 sg13g2_decap_8 FILLER_19_600 ();
 sg13g2_decap_8 FILLER_19_607 ();
 sg13g2_decap_8 FILLER_19_614 ();
 sg13g2_decap_8 FILLER_19_621 ();
 sg13g2_decap_8 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_635 ();
 sg13g2_decap_8 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_649 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_decap_8 FILLER_19_663 ();
 sg13g2_decap_8 FILLER_19_670 ();
 sg13g2_decap_8 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_684 ();
 sg13g2_decap_8 FILLER_19_691 ();
 sg13g2_decap_8 FILLER_19_698 ();
 sg13g2_decap_8 FILLER_19_705 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_719 ();
 sg13g2_decap_8 FILLER_19_726 ();
 sg13g2_decap_8 FILLER_19_733 ();
 sg13g2_decap_8 FILLER_19_740 ();
 sg13g2_decap_8 FILLER_19_747 ();
 sg13g2_decap_8 FILLER_19_754 ();
 sg13g2_decap_8 FILLER_19_761 ();
 sg13g2_decap_8 FILLER_19_768 ();
 sg13g2_decap_8 FILLER_19_775 ();
 sg13g2_decap_8 FILLER_19_782 ();
 sg13g2_decap_8 FILLER_19_789 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_decap_8 FILLER_19_824 ();
 sg13g2_decap_8 FILLER_19_831 ();
 sg13g2_decap_8 FILLER_19_838 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_fill_2 FILLER_19_859 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_17 ();
 sg13g2_decap_4 FILLER_20_24 ();
 sg13g2_fill_2 FILLER_20_94 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_decap_4 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_decap_4 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_4 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_4 FILLER_20_253 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_294 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_fill_1 FILLER_20_340 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_fill_2 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_371 ();
 sg13g2_fill_2 FILLER_20_389 ();
 sg13g2_fill_1 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_412 ();
 sg13g2_fill_2 FILLER_20_419 ();
 sg13g2_fill_1 FILLER_20_421 ();
 sg13g2_decap_4 FILLER_20_436 ();
 sg13g2_fill_2 FILLER_20_440 ();
 sg13g2_fill_1 FILLER_20_451 ();
 sg13g2_decap_8 FILLER_20_461 ();
 sg13g2_fill_1 FILLER_20_468 ();
 sg13g2_decap_8 FILLER_20_478 ();
 sg13g2_decap_8 FILLER_20_485 ();
 sg13g2_decap_8 FILLER_20_492 ();
 sg13g2_decap_8 FILLER_20_508 ();
 sg13g2_fill_2 FILLER_20_524 ();
 sg13g2_fill_1 FILLER_20_526 ();
 sg13g2_fill_1 FILLER_20_549 ();
 sg13g2_fill_2 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_589 ();
 sg13g2_decap_8 FILLER_20_596 ();
 sg13g2_decap_8 FILLER_20_603 ();
 sg13g2_decap_8 FILLER_20_610 ();
 sg13g2_decap_8 FILLER_20_617 ();
 sg13g2_decap_8 FILLER_20_624 ();
 sg13g2_decap_8 FILLER_20_631 ();
 sg13g2_decap_8 FILLER_20_638 ();
 sg13g2_decap_8 FILLER_20_645 ();
 sg13g2_decap_8 FILLER_20_652 ();
 sg13g2_decap_8 FILLER_20_659 ();
 sg13g2_decap_8 FILLER_20_666 ();
 sg13g2_decap_8 FILLER_20_673 ();
 sg13g2_decap_8 FILLER_20_680 ();
 sg13g2_decap_8 FILLER_20_687 ();
 sg13g2_decap_8 FILLER_20_694 ();
 sg13g2_decap_8 FILLER_20_701 ();
 sg13g2_decap_8 FILLER_20_708 ();
 sg13g2_decap_8 FILLER_20_715 ();
 sg13g2_decap_8 FILLER_20_722 ();
 sg13g2_decap_8 FILLER_20_729 ();
 sg13g2_decap_8 FILLER_20_736 ();
 sg13g2_decap_8 FILLER_20_743 ();
 sg13g2_decap_8 FILLER_20_750 ();
 sg13g2_decap_8 FILLER_20_757 ();
 sg13g2_decap_8 FILLER_20_764 ();
 sg13g2_decap_8 FILLER_20_771 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_decap_8 FILLER_20_785 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_8 FILLER_20_799 ();
 sg13g2_decap_8 FILLER_20_806 ();
 sg13g2_decap_8 FILLER_20_813 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_decap_8 FILLER_20_848 ();
 sg13g2_decap_8 FILLER_20_855 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_41 ();
 sg13g2_fill_2 FILLER_21_45 ();
 sg13g2_decap_8 FILLER_21_51 ();
 sg13g2_decap_4 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_62 ();
 sg13g2_fill_2 FILLER_21_110 ();
 sg13g2_decap_8 FILLER_21_135 ();
 sg13g2_decap_4 FILLER_21_142 ();
 sg13g2_fill_2 FILLER_21_146 ();
 sg13g2_decap_4 FILLER_21_153 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_180 ();
 sg13g2_decap_8 FILLER_21_187 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_4 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_decap_4 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_4 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_decap_4 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_329 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_fill_2 FILLER_21_398 ();
 sg13g2_fill_2 FILLER_21_410 ();
 sg13g2_fill_1 FILLER_21_412 ();
 sg13g2_fill_1 FILLER_21_418 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_fill_2 FILLER_21_430 ();
 sg13g2_decap_4 FILLER_21_468 ();
 sg13g2_fill_2 FILLER_21_472 ();
 sg13g2_decap_4 FILLER_21_518 ();
 sg13g2_fill_2 FILLER_21_534 ();
 sg13g2_fill_1 FILLER_21_570 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_63 ();
 sg13g2_decap_4 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_138 ();
 sg13g2_decap_4 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_166 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_4 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_fill_2 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_451 ();
 sg13g2_decap_8 FILLER_22_516 ();
 sg13g2_decap_4 FILLER_22_523 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_4 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_611 ();
 sg13g2_decap_8 FILLER_22_618 ();
 sg13g2_decap_8 FILLER_22_625 ();
 sg13g2_decap_8 FILLER_22_632 ();
 sg13g2_decap_8 FILLER_22_639 ();
 sg13g2_decap_8 FILLER_22_646 ();
 sg13g2_decap_8 FILLER_22_653 ();
 sg13g2_decap_8 FILLER_22_660 ();
 sg13g2_decap_8 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_674 ();
 sg13g2_decap_8 FILLER_22_681 ();
 sg13g2_decap_8 FILLER_22_688 ();
 sg13g2_decap_8 FILLER_22_695 ();
 sg13g2_decap_8 FILLER_22_702 ();
 sg13g2_decap_8 FILLER_22_709 ();
 sg13g2_decap_8 FILLER_22_716 ();
 sg13g2_decap_8 FILLER_22_723 ();
 sg13g2_decap_8 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_744 ();
 sg13g2_decap_8 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_758 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_decap_8 FILLER_22_779 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_793 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_decap_8 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_842 ();
 sg13g2_decap_8 FILLER_22_849 ();
 sg13g2_decap_4 FILLER_22_856 ();
 sg13g2_fill_2 FILLER_22_860 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_89 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_4 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_4 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_251 ();
 sg13g2_decap_4 FILLER_23_255 ();
 sg13g2_decap_4 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_272 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_decap_4 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_317 ();
 sg13g2_fill_2 FILLER_23_331 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_fill_2 FILLER_23_393 ();
 sg13g2_decap_4 FILLER_23_415 ();
 sg13g2_fill_2 FILLER_23_447 ();
 sg13g2_fill_1 FILLER_23_449 ();
 sg13g2_fill_1 FILLER_23_495 ();
 sg13g2_decap_4 FILLER_23_530 ();
 sg13g2_fill_1 FILLER_23_534 ();
 sg13g2_fill_2 FILLER_23_601 ();
 sg13g2_decap_8 FILLER_23_612 ();
 sg13g2_decap_8 FILLER_23_619 ();
 sg13g2_decap_8 FILLER_23_626 ();
 sg13g2_decap_8 FILLER_23_633 ();
 sg13g2_decap_8 FILLER_23_640 ();
 sg13g2_decap_8 FILLER_23_647 ();
 sg13g2_decap_8 FILLER_23_654 ();
 sg13g2_decap_8 FILLER_23_661 ();
 sg13g2_decap_8 FILLER_23_668 ();
 sg13g2_decap_8 FILLER_23_675 ();
 sg13g2_decap_8 FILLER_23_682 ();
 sg13g2_decap_8 FILLER_23_689 ();
 sg13g2_decap_8 FILLER_23_696 ();
 sg13g2_decap_8 FILLER_23_703 ();
 sg13g2_decap_8 FILLER_23_710 ();
 sg13g2_decap_8 FILLER_23_717 ();
 sg13g2_decap_8 FILLER_23_724 ();
 sg13g2_decap_8 FILLER_23_731 ();
 sg13g2_decap_8 FILLER_23_738 ();
 sg13g2_decap_8 FILLER_23_745 ();
 sg13g2_decap_8 FILLER_23_752 ();
 sg13g2_decap_8 FILLER_23_759 ();
 sg13g2_decap_8 FILLER_23_766 ();
 sg13g2_decap_8 FILLER_23_773 ();
 sg13g2_decap_8 FILLER_23_780 ();
 sg13g2_decap_8 FILLER_23_787 ();
 sg13g2_decap_8 FILLER_23_794 ();
 sg13g2_decap_8 FILLER_23_801 ();
 sg13g2_decap_8 FILLER_23_808 ();
 sg13g2_decap_8 FILLER_23_815 ();
 sg13g2_decap_8 FILLER_23_822 ();
 sg13g2_decap_8 FILLER_23_829 ();
 sg13g2_decap_8 FILLER_23_836 ();
 sg13g2_decap_8 FILLER_23_843 ();
 sg13g2_decap_8 FILLER_23_850 ();
 sg13g2_decap_4 FILLER_23_857 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_69 ();
 sg13g2_fill_1 FILLER_24_71 ();
 sg13g2_decap_4 FILLER_24_92 ();
 sg13g2_fill_1 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_121 ();
 sg13g2_decap_8 FILLER_24_136 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_decap_4 FILLER_24_150 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_181 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_216 ();
 sg13g2_decap_8 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_fill_2 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_424 ();
 sg13g2_fill_1 FILLER_24_478 ();
 sg13g2_fill_2 FILLER_24_489 ();
 sg13g2_fill_1 FILLER_24_491 ();
 sg13g2_fill_1 FILLER_24_499 ();
 sg13g2_decap_8 FILLER_24_520 ();
 sg13g2_fill_1 FILLER_24_527 ();
 sg13g2_decap_4 FILLER_24_541 ();
 sg13g2_fill_1 FILLER_24_545 ();
 sg13g2_fill_1 FILLER_24_555 ();
 sg13g2_fill_2 FILLER_24_580 ();
 sg13g2_decap_4 FILLER_24_587 ();
 sg13g2_fill_1 FILLER_24_591 ();
 sg13g2_decap_8 FILLER_24_618 ();
 sg13g2_decap_8 FILLER_24_625 ();
 sg13g2_decap_8 FILLER_24_632 ();
 sg13g2_decap_8 FILLER_24_639 ();
 sg13g2_decap_8 FILLER_24_646 ();
 sg13g2_decap_8 FILLER_24_653 ();
 sg13g2_decap_8 FILLER_24_660 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_decap_8 FILLER_24_674 ();
 sg13g2_decap_8 FILLER_24_681 ();
 sg13g2_decap_8 FILLER_24_688 ();
 sg13g2_decap_8 FILLER_24_695 ();
 sg13g2_decap_8 FILLER_24_702 ();
 sg13g2_decap_8 FILLER_24_709 ();
 sg13g2_decap_8 FILLER_24_716 ();
 sg13g2_decap_8 FILLER_24_723 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_decap_8 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_744 ();
 sg13g2_decap_8 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_758 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_786 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_842 ();
 sg13g2_decap_8 FILLER_24_849 ();
 sg13g2_decap_4 FILLER_24_856 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_fill_1 FILLER_25_53 ();
 sg13g2_decap_4 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_62 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_4 FILLER_25_117 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_fill_2 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_4 FILLER_25_422 ();
 sg13g2_decap_4 FILLER_25_460 ();
 sg13g2_decap_4 FILLER_25_499 ();
 sg13g2_decap_8 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_fill_2 FILLER_25_550 ();
 sg13g2_fill_1 FILLER_25_552 ();
 sg13g2_fill_1 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_585 ();
 sg13g2_fill_2 FILLER_25_592 ();
 sg13g2_fill_1 FILLER_25_594 ();
 sg13g2_decap_8 FILLER_25_604 ();
 sg13g2_decap_8 FILLER_25_611 ();
 sg13g2_decap_8 FILLER_25_618 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_decap_8 FILLER_25_660 ();
 sg13g2_decap_8 FILLER_25_667 ();
 sg13g2_decap_8 FILLER_25_674 ();
 sg13g2_decap_8 FILLER_25_681 ();
 sg13g2_decap_8 FILLER_25_688 ();
 sg13g2_decap_8 FILLER_25_695 ();
 sg13g2_decap_8 FILLER_25_702 ();
 sg13g2_decap_8 FILLER_25_709 ();
 sg13g2_decap_8 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_737 ();
 sg13g2_decap_8 FILLER_25_744 ();
 sg13g2_decap_8 FILLER_25_751 ();
 sg13g2_decap_8 FILLER_25_758 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_4 FILLER_25_856 ();
 sg13g2_fill_2 FILLER_25_860 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_23 ();
 sg13g2_fill_1 FILLER_26_44 ();
 sg13g2_decap_8 FILLER_26_71 ();
 sg13g2_decap_4 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_94 ();
 sg13g2_decap_4 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_4 FILLER_26_271 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_4 FILLER_26_324 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_4 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_fill_2 FILLER_26_443 ();
 sg13g2_fill_1 FILLER_26_445 ();
 sg13g2_fill_1 FILLER_26_455 ();
 sg13g2_fill_2 FILLER_26_482 ();
 sg13g2_fill_1 FILLER_26_484 ();
 sg13g2_fill_1 FILLER_26_494 ();
 sg13g2_decap_4 FILLER_26_504 ();
 sg13g2_fill_1 FILLER_26_526 ();
 sg13g2_decap_8 FILLER_26_610 ();
 sg13g2_decap_8 FILLER_26_617 ();
 sg13g2_decap_4 FILLER_26_624 ();
 sg13g2_decap_8 FILLER_26_632 ();
 sg13g2_decap_8 FILLER_26_639 ();
 sg13g2_decap_8 FILLER_26_646 ();
 sg13g2_decap_8 FILLER_26_653 ();
 sg13g2_decap_8 FILLER_26_660 ();
 sg13g2_decap_8 FILLER_26_667 ();
 sg13g2_decap_8 FILLER_26_674 ();
 sg13g2_decap_8 FILLER_26_681 ();
 sg13g2_decap_8 FILLER_26_688 ();
 sg13g2_decap_8 FILLER_26_695 ();
 sg13g2_decap_8 FILLER_26_702 ();
 sg13g2_decap_8 FILLER_26_709 ();
 sg13g2_decap_8 FILLER_26_716 ();
 sg13g2_decap_8 FILLER_26_723 ();
 sg13g2_decap_8 FILLER_26_730 ();
 sg13g2_decap_8 FILLER_26_737 ();
 sg13g2_decap_8 FILLER_26_744 ();
 sg13g2_decap_8 FILLER_26_751 ();
 sg13g2_decap_8 FILLER_26_758 ();
 sg13g2_decap_8 FILLER_26_765 ();
 sg13g2_decap_8 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_779 ();
 sg13g2_decap_8 FILLER_26_786 ();
 sg13g2_decap_8 FILLER_26_793 ();
 sg13g2_decap_8 FILLER_26_800 ();
 sg13g2_decap_8 FILLER_26_807 ();
 sg13g2_decap_8 FILLER_26_814 ();
 sg13g2_decap_8 FILLER_26_821 ();
 sg13g2_decap_8 FILLER_26_828 ();
 sg13g2_decap_8 FILLER_26_835 ();
 sg13g2_decap_8 FILLER_26_842 ();
 sg13g2_decap_8 FILLER_26_849 ();
 sg13g2_decap_4 FILLER_26_856 ();
 sg13g2_fill_2 FILLER_26_860 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_66 ();
 sg13g2_decap_4 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_104 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_2 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_decap_4 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_fill_1 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_4 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_decap_4 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_fill_2 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_decap_4 FILLER_27_437 ();
 sg13g2_decap_4 FILLER_27_446 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_fill_1 FILLER_27_467 ();
 sg13g2_fill_2 FILLER_27_482 ();
 sg13g2_fill_1 FILLER_27_484 ();
 sg13g2_decap_8 FILLER_27_528 ();
 sg13g2_decap_8 FILLER_27_535 ();
 sg13g2_fill_1 FILLER_27_542 ();
 sg13g2_decap_8 FILLER_27_552 ();
 sg13g2_decap_4 FILLER_27_559 ();
 sg13g2_fill_2 FILLER_27_563 ();
 sg13g2_decap_4 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_decap_8 FILLER_27_606 ();
 sg13g2_decap_4 FILLER_27_613 ();
 sg13g2_fill_2 FILLER_27_617 ();
 sg13g2_decap_4 FILLER_27_652 ();
 sg13g2_fill_2 FILLER_27_656 ();
 sg13g2_decap_8 FILLER_27_684 ();
 sg13g2_decap_8 FILLER_27_691 ();
 sg13g2_fill_2 FILLER_27_698 ();
 sg13g2_fill_1 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_4 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_734 ();
 sg13g2_decap_8 FILLER_27_741 ();
 sg13g2_decap_8 FILLER_27_748 ();
 sg13g2_decap_8 FILLER_27_755 ();
 sg13g2_decap_8 FILLER_27_762 ();
 sg13g2_decap_8 FILLER_27_769 ();
 sg13g2_decap_8 FILLER_27_776 ();
 sg13g2_decap_8 FILLER_27_783 ();
 sg13g2_decap_8 FILLER_27_790 ();
 sg13g2_decap_8 FILLER_27_797 ();
 sg13g2_decap_8 FILLER_27_804 ();
 sg13g2_decap_8 FILLER_27_811 ();
 sg13g2_decap_8 FILLER_27_818 ();
 sg13g2_decap_8 FILLER_27_825 ();
 sg13g2_decap_8 FILLER_27_832 ();
 sg13g2_decap_8 FILLER_27_839 ();
 sg13g2_decap_8 FILLER_27_846 ();
 sg13g2_decap_8 FILLER_27_853 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_20 ();
 sg13g2_fill_2 FILLER_28_31 ();
 sg13g2_fill_1 FILLER_28_33 ();
 sg13g2_decap_8 FILLER_28_69 ();
 sg13g2_decap_4 FILLER_28_76 ();
 sg13g2_fill_1 FILLER_28_80 ();
 sg13g2_fill_2 FILLER_28_93 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_189 ();
 sg13g2_fill_1 FILLER_28_191 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_245 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_decap_4 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_decap_4 FILLER_28_323 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_decap_4 FILLER_28_340 ();
 sg13g2_decap_4 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_fill_2 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_fill_1 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_461 ();
 sg13g2_decap_8 FILLER_28_468 ();
 sg13g2_fill_2 FILLER_28_475 ();
 sg13g2_fill_1 FILLER_28_477 ();
 sg13g2_decap_8 FILLER_28_492 ();
 sg13g2_decap_4 FILLER_28_504 ();
 sg13g2_fill_1 FILLER_28_508 ();
 sg13g2_decap_4 FILLER_28_535 ();
 sg13g2_fill_2 FILLER_28_539 ();
 sg13g2_decap_4 FILLER_28_619 ();
 sg13g2_fill_1 FILLER_28_623 ();
 sg13g2_fill_2 FILLER_28_641 ();
 sg13g2_fill_2 FILLER_28_666 ();
 sg13g2_decap_4 FILLER_28_680 ();
 sg13g2_decap_4 FILLER_28_688 ();
 sg13g2_decap_8 FILLER_28_738 ();
 sg13g2_decap_8 FILLER_28_745 ();
 sg13g2_decap_8 FILLER_28_752 ();
 sg13g2_decap_8 FILLER_28_759 ();
 sg13g2_decap_8 FILLER_28_766 ();
 sg13g2_decap_8 FILLER_28_773 ();
 sg13g2_decap_8 FILLER_28_780 ();
 sg13g2_decap_8 FILLER_28_787 ();
 sg13g2_decap_8 FILLER_28_794 ();
 sg13g2_decap_8 FILLER_28_801 ();
 sg13g2_decap_8 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_815 ();
 sg13g2_decap_8 FILLER_28_822 ();
 sg13g2_decap_8 FILLER_28_829 ();
 sg13g2_decap_8 FILLER_28_836 ();
 sg13g2_decap_8 FILLER_28_843 ();
 sg13g2_decap_8 FILLER_28_850 ();
 sg13g2_decap_4 FILLER_28_857 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_54 ();
 sg13g2_decap_8 FILLER_29_61 ();
 sg13g2_decap_8 FILLER_29_68 ();
 sg13g2_decap_4 FILLER_29_75 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_decap_4 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_decap_4 FILLER_29_174 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_decap_4 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_271 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_324 ();
 sg13g2_decap_4 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_fill_2 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_29_426 ();
 sg13g2_fill_2 FILLER_29_527 ();
 sg13g2_decap_4 FILLER_29_538 ();
 sg13g2_fill_1 FILLER_29_542 ();
 sg13g2_fill_2 FILLER_29_552 ();
 sg13g2_decap_8 FILLER_29_568 ();
 sg13g2_fill_2 FILLER_29_575 ();
 sg13g2_decap_8 FILLER_29_603 ();
 sg13g2_decap_4 FILLER_29_610 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_decap_8 FILLER_29_629 ();
 sg13g2_fill_2 FILLER_29_636 ();
 sg13g2_fill_2 FILLER_29_643 ();
 sg13g2_fill_1 FILLER_29_645 ();
 sg13g2_decap_8 FILLER_29_655 ();
 sg13g2_fill_2 FILLER_29_662 ();
 sg13g2_fill_2 FILLER_29_699 ();
 sg13g2_decap_8 FILLER_29_711 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_decap_8 FILLER_29_746 ();
 sg13g2_decap_8 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_decap_8 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_4 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_decap_8 FILLER_30_86 ();
 sg13g2_decap_8 FILLER_30_93 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_decap_8 FILLER_30_145 ();
 sg13g2_decap_4 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_decap_4 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_decap_4 FILLER_30_205 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_242 ();
 sg13g2_decap_4 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_decap_4 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_4 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_decap_4 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_378 ();
 sg13g2_fill_1 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_459 ();
 sg13g2_decap_8 FILLER_30_466 ();
 sg13g2_decap_4 FILLER_30_473 ();
 sg13g2_fill_2 FILLER_30_477 ();
 sg13g2_fill_2 FILLER_30_487 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_4 FILLER_30_525 ();
 sg13g2_decap_4 FILLER_30_559 ();
 sg13g2_fill_2 FILLER_30_568 ();
 sg13g2_fill_1 FILLER_30_570 ();
 sg13g2_fill_2 FILLER_30_599 ();
 sg13g2_decap_4 FILLER_30_627 ();
 sg13g2_fill_1 FILLER_30_661 ();
 sg13g2_decap_8 FILLER_30_681 ();
 sg13g2_fill_1 FILLER_30_688 ();
 sg13g2_fill_2 FILLER_30_692 ();
 sg13g2_fill_2 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_8 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_decap_8 FILLER_31_156 ();
 sg13g2_decap_4 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_172 ();
 sg13g2_fill_2 FILLER_31_178 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_decap_4 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_236 ();
 sg13g2_decap_8 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_decap_4 FILLER_31_395 ();
 sg13g2_fill_2 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_476 ();
 sg13g2_fill_2 FILLER_31_501 ();
 sg13g2_fill_1 FILLER_31_503 ();
 sg13g2_decap_4 FILLER_31_519 ();
 sg13g2_fill_1 FILLER_31_537 ();
 sg13g2_fill_2 FILLER_31_578 ();
 sg13g2_decap_8 FILLER_31_635 ();
 sg13g2_fill_1 FILLER_31_642 ();
 sg13g2_decap_4 FILLER_31_652 ();
 sg13g2_fill_1 FILLER_31_656 ();
 sg13g2_decap_4 FILLER_31_677 ();
 sg13g2_fill_2 FILLER_31_681 ();
 sg13g2_fill_2 FILLER_31_691 ();
 sg13g2_fill_1 FILLER_31_707 ();
 sg13g2_fill_2 FILLER_31_718 ();
 sg13g2_fill_1 FILLER_31_720 ();
 sg13g2_fill_2 FILLER_31_733 ();
 sg13g2_fill_1 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_745 ();
 sg13g2_decap_8 FILLER_31_752 ();
 sg13g2_decap_8 FILLER_31_759 ();
 sg13g2_decap_8 FILLER_31_766 ();
 sg13g2_decap_8 FILLER_31_773 ();
 sg13g2_decap_8 FILLER_31_780 ();
 sg13g2_decap_8 FILLER_31_787 ();
 sg13g2_decap_8 FILLER_31_794 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_4 FILLER_31_857 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_85 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_257 ();
 sg13g2_decap_8 FILLER_32_264 ();
 sg13g2_fill_2 FILLER_32_271 ();
 sg13g2_fill_1 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_281 ();
 sg13g2_decap_4 FILLER_32_288 ();
 sg13g2_decap_8 FILLER_32_303 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_decap_4 FILLER_32_367 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_fill_1 FILLER_32_423 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_fill_1 FILLER_32_476 ();
 sg13g2_fill_2 FILLER_32_503 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_fill_1 FILLER_32_520 ();
 sg13g2_decap_4 FILLER_32_526 ();
 sg13g2_decap_4 FILLER_32_538 ();
 sg13g2_decap_4 FILLER_32_546 ();
 sg13g2_decap_4 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_569 ();
 sg13g2_decap_4 FILLER_32_576 ();
 sg13g2_fill_1 FILLER_32_599 ();
 sg13g2_decap_4 FILLER_32_621 ();
 sg13g2_fill_2 FILLER_32_632 ();
 sg13g2_decap_8 FILLER_32_660 ();
 sg13g2_decap_8 FILLER_32_667 ();
 sg13g2_decap_8 FILLER_32_674 ();
 sg13g2_decap_4 FILLER_32_681 ();
 sg13g2_fill_1 FILLER_32_685 ();
 sg13g2_fill_2 FILLER_32_719 ();
 sg13g2_decap_8 FILLER_32_747 ();
 sg13g2_decap_8 FILLER_32_754 ();
 sg13g2_decap_8 FILLER_32_761 ();
 sg13g2_decap_8 FILLER_32_768 ();
 sg13g2_decap_8 FILLER_32_775 ();
 sg13g2_decap_8 FILLER_32_782 ();
 sg13g2_decap_8 FILLER_32_789 ();
 sg13g2_decap_8 FILLER_32_796 ();
 sg13g2_decap_8 FILLER_32_803 ();
 sg13g2_decap_8 FILLER_32_810 ();
 sg13g2_decap_8 FILLER_32_817 ();
 sg13g2_decap_8 FILLER_32_824 ();
 sg13g2_decap_8 FILLER_32_831 ();
 sg13g2_decap_8 FILLER_32_838 ();
 sg13g2_decap_8 FILLER_32_845 ();
 sg13g2_decap_8 FILLER_32_852 ();
 sg13g2_fill_2 FILLER_32_859 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_123 ();
 sg13g2_decap_4 FILLER_33_134 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_decap_4 FILLER_33_167 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_4 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_2 FILLER_33_235 ();
 sg13g2_decap_4 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_fill_2 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_489 ();
 sg13g2_fill_2 FILLER_33_496 ();
 sg13g2_fill_1 FILLER_33_498 ();
 sg13g2_fill_2 FILLER_33_549 ();
 sg13g2_fill_1 FILLER_33_551 ();
 sg13g2_decap_4 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_565 ();
 sg13g2_fill_1 FILLER_33_592 ();
 sg13g2_decap_8 FILLER_33_619 ();
 sg13g2_fill_1 FILLER_33_631 ();
 sg13g2_fill_2 FILLER_33_635 ();
 sg13g2_fill_1 FILLER_33_637 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_1 FILLER_33_656 ();
 sg13g2_fill_2 FILLER_33_665 ();
 sg13g2_fill_2 FILLER_33_703 ();
 sg13g2_fill_1 FILLER_33_724 ();
 sg13g2_decap_8 FILLER_33_751 ();
 sg13g2_decap_8 FILLER_33_758 ();
 sg13g2_decap_8 FILLER_33_765 ();
 sg13g2_decap_8 FILLER_33_772 ();
 sg13g2_decap_8 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_decap_8 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_33_828 ();
 sg13g2_decap_8 FILLER_33_835 ();
 sg13g2_decap_8 FILLER_33_842 ();
 sg13g2_decap_8 FILLER_33_849 ();
 sg13g2_decap_4 FILLER_33_856 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_fill_2 FILLER_34_68 ();
 sg13g2_fill_1 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_294 ();
 sg13g2_fill_1 FILLER_34_296 ();
 sg13g2_decap_4 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_fill_1 FILLER_34_390 ();
 sg13g2_fill_2 FILLER_34_396 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_34_442 ();
 sg13g2_fill_1 FILLER_34_449 ();
 sg13g2_decap_8 FILLER_34_488 ();
 sg13g2_decap_8 FILLER_34_513 ();
 sg13g2_decap_4 FILLER_34_520 ();
 sg13g2_fill_2 FILLER_34_524 ();
 sg13g2_fill_2 FILLER_34_582 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_decap_4 FILLER_34_614 ();
 sg13g2_decap_8 FILLER_34_638 ();
 sg13g2_decap_8 FILLER_34_645 ();
 sg13g2_decap_4 FILLER_34_652 ();
 sg13g2_fill_1 FILLER_34_656 ();
 sg13g2_fill_2 FILLER_34_665 ();
 sg13g2_fill_1 FILLER_34_667 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_fill_2 FILLER_34_691 ();
 sg13g2_decap_4 FILLER_34_698 ();
 sg13g2_fill_2 FILLER_34_717 ();
 sg13g2_fill_2 FILLER_34_723 ();
 sg13g2_fill_2 FILLER_34_734 ();
 sg13g2_decap_8 FILLER_34_745 ();
 sg13g2_decap_8 FILLER_34_752 ();
 sg13g2_decap_8 FILLER_34_759 ();
 sg13g2_decap_8 FILLER_34_766 ();
 sg13g2_decap_8 FILLER_34_773 ();
 sg13g2_decap_8 FILLER_34_780 ();
 sg13g2_decap_8 FILLER_34_787 ();
 sg13g2_decap_8 FILLER_34_794 ();
 sg13g2_decap_8 FILLER_34_801 ();
 sg13g2_decap_8 FILLER_34_808 ();
 sg13g2_decap_8 FILLER_34_815 ();
 sg13g2_decap_8 FILLER_34_822 ();
 sg13g2_decap_8 FILLER_34_829 ();
 sg13g2_decap_8 FILLER_34_836 ();
 sg13g2_decap_8 FILLER_34_843 ();
 sg13g2_decap_8 FILLER_34_850 ();
 sg13g2_decap_4 FILLER_34_857 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_decap_4 FILLER_35_113 ();
 sg13g2_fill_2 FILLER_35_117 ();
 sg13g2_fill_2 FILLER_35_129 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_decap_4 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_181 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_decap_4 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_decap_8 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_257 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_fill_2 FILLER_35_285 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_decap_8 FILLER_35_306 ();
 sg13g2_decap_4 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_334 ();
 sg13g2_decap_8 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_fill_2 FILLER_35_359 ();
 sg13g2_fill_2 FILLER_35_417 ();
 sg13g2_fill_1 FILLER_35_419 ();
 sg13g2_fill_2 FILLER_35_472 ();
 sg13g2_fill_1 FILLER_35_474 ();
 sg13g2_fill_1 FILLER_35_493 ();
 sg13g2_decap_8 FILLER_35_502 ();
 sg13g2_decap_8 FILLER_35_509 ();
 sg13g2_decap_8 FILLER_35_516 ();
 sg13g2_decap_8 FILLER_35_523 ();
 sg13g2_fill_2 FILLER_35_530 ();
 sg13g2_decap_4 FILLER_35_540 ();
 sg13g2_fill_1 FILLER_35_553 ();
 sg13g2_fill_2 FILLER_35_559 ();
 sg13g2_fill_1 FILLER_35_561 ();
 sg13g2_decap_4 FILLER_35_587 ();
 sg13g2_fill_1 FILLER_35_599 ();
 sg13g2_decap_4 FILLER_35_624 ();
 sg13g2_fill_2 FILLER_35_628 ();
 sg13g2_decap_8 FILLER_35_656 ();
 sg13g2_decap_4 FILLER_35_663 ();
 sg13g2_fill_2 FILLER_35_667 ();
 sg13g2_decap_8 FILLER_35_678 ();
 sg13g2_fill_2 FILLER_35_685 ();
 sg13g2_fill_2 FILLER_35_708 ();
 sg13g2_fill_1 FILLER_35_736 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_4 FILLER_36_172 ();
 sg13g2_decap_4 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_270 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_decap_4 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_383 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_36_436 ();
 sg13g2_decap_8 FILLER_36_443 ();
 sg13g2_fill_2 FILLER_36_450 ();
 sg13g2_decap_4 FILLER_36_467 ();
 sg13g2_fill_1 FILLER_36_471 ();
 sg13g2_decap_4 FILLER_36_477 ();
 sg13g2_fill_2 FILLER_36_481 ();
 sg13g2_fill_1 FILLER_36_568 ();
 sg13g2_decap_4 FILLER_36_595 ();
 sg13g2_fill_1 FILLER_36_599 ();
 sg13g2_fill_1 FILLER_36_617 ();
 sg13g2_decap_4 FILLER_36_644 ();
 sg13g2_fill_1 FILLER_36_648 ();
 sg13g2_decap_4 FILLER_36_685 ();
 sg13g2_fill_2 FILLER_36_689 ();
 sg13g2_decap_8 FILLER_36_696 ();
 sg13g2_decap_8 FILLER_36_703 ();
 sg13g2_decap_8 FILLER_36_710 ();
 sg13g2_decap_8 FILLER_36_717 ();
 sg13g2_decap_8 FILLER_36_724 ();
 sg13g2_fill_1 FILLER_36_746 ();
 sg13g2_decap_8 FILLER_36_761 ();
 sg13g2_decap_8 FILLER_36_768 ();
 sg13g2_decap_8 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_782 ();
 sg13g2_decap_8 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_93 ();
 sg13g2_decap_4 FILLER_37_100 ();
 sg13g2_fill_2 FILLER_37_104 ();
 sg13g2_decap_8 FILLER_37_110 ();
 sg13g2_decap_8 FILLER_37_117 ();
 sg13g2_decap_4 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_190 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_204 ();
 sg13g2_decap_4 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_236 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_decap_4 FILLER_37_250 ();
 sg13g2_fill_2 FILLER_37_254 ();
 sg13g2_fill_1 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_8 FILLER_37_278 ();
 sg13g2_decap_4 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_decap_8 FILLER_37_321 ();
 sg13g2_fill_2 FILLER_37_328 ();
 sg13g2_fill_2 FILLER_37_366 ();
 sg13g2_fill_2 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_decap_8 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_37_457 ();
 sg13g2_decap_8 FILLER_37_464 ();
 sg13g2_decap_4 FILLER_37_471 ();
 sg13g2_fill_1 FILLER_37_475 ();
 sg13g2_fill_1 FILLER_37_487 ();
 sg13g2_decap_8 FILLER_37_512 ();
 sg13g2_decap_8 FILLER_37_519 ();
 sg13g2_decap_4 FILLER_37_526 ();
 sg13g2_fill_1 FILLER_37_530 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_2 FILLER_37_553 ();
 sg13g2_fill_1 FILLER_37_555 ();
 sg13g2_fill_2 FILLER_37_562 ();
 sg13g2_fill_1 FILLER_37_573 ();
 sg13g2_fill_2 FILLER_37_583 ();
 sg13g2_fill_1 FILLER_37_585 ();
 sg13g2_fill_2 FILLER_37_617 ();
 sg13g2_decap_8 FILLER_37_628 ();
 sg13g2_decap_4 FILLER_37_635 ();
 sg13g2_fill_1 FILLER_37_639 ();
 sg13g2_decap_8 FILLER_37_659 ();
 sg13g2_decap_8 FILLER_37_666 ();
 sg13g2_fill_2 FILLER_37_673 ();
 sg13g2_fill_2 FILLER_37_680 ();
 sg13g2_fill_2 FILLER_37_687 ();
 sg13g2_fill_1 FILLER_37_720 ();
 sg13g2_fill_1 FILLER_37_736 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_807 ();
 sg13g2_decap_8 FILLER_37_814 ();
 sg13g2_decap_8 FILLER_37_821 ();
 sg13g2_decap_8 FILLER_37_828 ();
 sg13g2_decap_8 FILLER_37_835 ();
 sg13g2_decap_8 FILLER_37_842 ();
 sg13g2_decap_8 FILLER_37_849 ();
 sg13g2_decap_4 FILLER_37_856 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_4 FILLER_38_98 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_decap_4 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_decap_4 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_decap_4 FILLER_38_171 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_2 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_237 ();
 sg13g2_decap_4 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_273 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_4 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_4 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_434 ();
 sg13g2_fill_1 FILLER_38_449 ();
 sg13g2_fill_1 FILLER_38_476 ();
 sg13g2_fill_1 FILLER_38_495 ();
 sg13g2_fill_2 FILLER_38_531 ();
 sg13g2_fill_1 FILLER_38_533 ();
 sg13g2_decap_8 FILLER_38_591 ();
 sg13g2_fill_1 FILLER_38_598 ();
 sg13g2_fill_2 FILLER_38_634 ();
 sg13g2_fill_1 FILLER_38_662 ();
 sg13g2_decap_4 FILLER_38_686 ();
 sg13g2_decap_4 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_721 ();
 sg13g2_fill_2 FILLER_38_741 ();
 sg13g2_fill_1 FILLER_38_743 ();
 sg13g2_decap_4 FILLER_38_765 ();
 sg13g2_fill_2 FILLER_38_769 ();
 sg13g2_decap_8 FILLER_38_775 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_810 ();
 sg13g2_decap_8 FILLER_38_817 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_8 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_838 ();
 sg13g2_decap_8 FILLER_38_845 ();
 sg13g2_decap_8 FILLER_38_852 ();
 sg13g2_fill_2 FILLER_38_859 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_4 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_60 ();
 sg13g2_fill_2 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_80 ();
 sg13g2_decap_8 FILLER_39_143 ();
 sg13g2_decap_8 FILLER_39_150 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_fill_2 FILLER_39_175 ();
 sg13g2_fill_1 FILLER_39_177 ();
 sg13g2_fill_2 FILLER_39_200 ();
 sg13g2_fill_2 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_decap_8 FILLER_39_215 ();
 sg13g2_decap_4 FILLER_39_222 ();
 sg13g2_fill_1 FILLER_39_226 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_275 ();
 sg13g2_fill_1 FILLER_39_277 ();
 sg13g2_fill_2 FILLER_39_286 ();
 sg13g2_fill_1 FILLER_39_288 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_fill_2 FILLER_39_301 ();
 sg13g2_fill_2 FILLER_39_347 ();
 sg13g2_fill_1 FILLER_39_349 ();
 sg13g2_fill_1 FILLER_39_394 ();
 sg13g2_decap_4 FILLER_39_410 ();
 sg13g2_fill_2 FILLER_39_414 ();
 sg13g2_decap_4 FILLER_39_420 ();
 sg13g2_fill_1 FILLER_39_424 ();
 sg13g2_fill_2 FILLER_39_434 ();
 sg13g2_decap_4 FILLER_39_467 ();
 sg13g2_fill_1 FILLER_39_471 ();
 sg13g2_decap_4 FILLER_39_484 ();
 sg13g2_fill_1 FILLER_39_488 ();
 sg13g2_decap_4 FILLER_39_510 ();
 sg13g2_fill_2 FILLER_39_514 ();
 sg13g2_decap_8 FILLER_39_520 ();
 sg13g2_decap_4 FILLER_39_572 ();
 sg13g2_fill_2 FILLER_39_580 ();
 sg13g2_decap_4 FILLER_39_586 ();
 sg13g2_fill_1 FILLER_39_590 ();
 sg13g2_fill_2 FILLER_39_616 ();
 sg13g2_fill_1 FILLER_39_618 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_fill_2 FILLER_39_630 ();
 sg13g2_decap_4 FILLER_39_656 ();
 sg13g2_fill_1 FILLER_39_660 ();
 sg13g2_decap_8 FILLER_39_666 ();
 sg13g2_fill_1 FILLER_39_673 ();
 sg13g2_fill_2 FILLER_39_678 ();
 sg13g2_fill_1 FILLER_39_680 ();
 sg13g2_fill_2 FILLER_39_685 ();
 sg13g2_fill_1 FILLER_39_687 ();
 sg13g2_fill_2 FILLER_39_698 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_4 FILLER_39_721 ();
 sg13g2_fill_2 FILLER_39_725 ();
 sg13g2_fill_1 FILLER_39_732 ();
 sg13g2_fill_2 FILLER_39_739 ();
 sg13g2_fill_1 FILLER_39_741 ();
 sg13g2_decap_8 FILLER_39_759 ();
 sg13g2_decap_4 FILLER_39_766 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_4 FILLER_40_42 ();
 sg13g2_fill_1 FILLER_40_46 ();
 sg13g2_decap_8 FILLER_40_89 ();
 sg13g2_decap_4 FILLER_40_96 ();
 sg13g2_fill_1 FILLER_40_100 ();
 sg13g2_decap_8 FILLER_40_110 ();
 sg13g2_decap_8 FILLER_40_117 ();
 sg13g2_decap_4 FILLER_40_124 ();
 sg13g2_decap_8 FILLER_40_132 ();
 sg13g2_fill_2 FILLER_40_139 ();
 sg13g2_decap_8 FILLER_40_220 ();
 sg13g2_decap_4 FILLER_40_227 ();
 sg13g2_fill_2 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_fill_2 FILLER_40_291 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_fill_1 FILLER_40_378 ();
 sg13g2_decap_4 FILLER_40_391 ();
 sg13g2_fill_2 FILLER_40_395 ();
 sg13g2_fill_2 FILLER_40_405 ();
 sg13g2_fill_2 FILLER_40_441 ();
 sg13g2_fill_1 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_482 ();
 sg13g2_fill_2 FILLER_40_489 ();
 sg13g2_fill_1 FILLER_40_491 ();
 sg13g2_decap_8 FILLER_40_500 ();
 sg13g2_fill_1 FILLER_40_507 ();
 sg13g2_decap_8 FILLER_40_516 ();
 sg13g2_decap_8 FILLER_40_523 ();
 sg13g2_fill_1 FILLER_40_530 ();
 sg13g2_fill_1 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_568 ();
 sg13g2_decap_4 FILLER_40_575 ();
 sg13g2_fill_2 FILLER_40_579 ();
 sg13g2_decap_8 FILLER_40_585 ();
 sg13g2_fill_2 FILLER_40_592 ();
 sg13g2_fill_1 FILLER_40_594 ();
 sg13g2_fill_2 FILLER_40_604 ();
 sg13g2_fill_1 FILLER_40_606 ();
 sg13g2_decap_4 FILLER_40_624 ();
 sg13g2_fill_1 FILLER_40_628 ();
 sg13g2_decap_4 FILLER_40_651 ();
 sg13g2_fill_2 FILLER_40_655 ();
 sg13g2_decap_4 FILLER_40_661 ();
 sg13g2_fill_1 FILLER_40_665 ();
 sg13g2_fill_1 FILLER_40_684 ();
 sg13g2_fill_2 FILLER_40_714 ();
 sg13g2_fill_1 FILLER_40_733 ();
 sg13g2_decap_8 FILLER_40_773 ();
 sg13g2_decap_8 FILLER_40_780 ();
 sg13g2_decap_8 FILLER_40_787 ();
 sg13g2_decap_8 FILLER_40_794 ();
 sg13g2_decap_8 FILLER_40_801 ();
 sg13g2_decap_8 FILLER_40_808 ();
 sg13g2_decap_8 FILLER_40_815 ();
 sg13g2_decap_8 FILLER_40_822 ();
 sg13g2_decap_8 FILLER_40_829 ();
 sg13g2_decap_8 FILLER_40_836 ();
 sg13g2_decap_8 FILLER_40_843 ();
 sg13g2_decap_8 FILLER_40_850 ();
 sg13g2_decap_4 FILLER_40_857 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_4 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_78 ();
 sg13g2_fill_2 FILLER_41_116 ();
 sg13g2_fill_1 FILLER_41_118 ();
 sg13g2_decap_4 FILLER_41_137 ();
 sg13g2_fill_2 FILLER_41_141 ();
 sg13g2_decap_4 FILLER_41_147 ();
 sg13g2_fill_1 FILLER_41_156 ();
 sg13g2_fill_2 FILLER_41_162 ();
 sg13g2_fill_1 FILLER_41_164 ();
 sg13g2_decap_4 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_178 ();
 sg13g2_fill_1 FILLER_41_185 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_4 FILLER_41_210 ();
 sg13g2_fill_2 FILLER_41_214 ();
 sg13g2_decap_8 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_272 ();
 sg13g2_decap_4 FILLER_41_279 ();
 sg13g2_decap_4 FILLER_41_300 ();
 sg13g2_decap_8 FILLER_41_312 ();
 sg13g2_decap_4 FILLER_41_319 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_decap_8 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_347 ();
 sg13g2_fill_1 FILLER_41_354 ();
 sg13g2_decap_4 FILLER_41_360 ();
 sg13g2_fill_2 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_384 ();
 sg13g2_decap_4 FILLER_41_391 ();
 sg13g2_fill_2 FILLER_41_395 ();
 sg13g2_decap_8 FILLER_41_402 ();
 sg13g2_decap_8 FILLER_41_409 ();
 sg13g2_decap_4 FILLER_41_420 ();
 sg13g2_fill_1 FILLER_41_424 ();
 sg13g2_fill_2 FILLER_41_429 ();
 sg13g2_decap_4 FILLER_41_440 ();
 sg13g2_decap_4 FILLER_41_448 ();
 sg13g2_fill_1 FILLER_41_452 ();
 sg13g2_decap_8 FILLER_41_457 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_decap_4 FILLER_41_478 ();
 sg13g2_fill_1 FILLER_41_482 ();
 sg13g2_fill_2 FILLER_41_499 ();
 sg13g2_fill_2 FILLER_41_515 ();
 sg13g2_fill_1 FILLER_41_517 ();
 sg13g2_fill_2 FILLER_41_526 ();
 sg13g2_fill_1 FILLER_41_528 ();
 sg13g2_fill_2 FILLER_41_572 ();
 sg13g2_fill_1 FILLER_41_574 ();
 sg13g2_decap_4 FILLER_41_595 ();
 sg13g2_fill_1 FILLER_41_599 ();
 sg13g2_decap_4 FILLER_41_634 ();
 sg13g2_fill_1 FILLER_41_638 ();
 sg13g2_decap_8 FILLER_41_643 ();
 sg13g2_fill_2 FILLER_41_650 ();
 sg13g2_decap_4 FILLER_41_696 ();
 sg13g2_fill_2 FILLER_41_700 ();
 sg13g2_decap_4 FILLER_41_715 ();
 sg13g2_fill_2 FILLER_41_719 ();
 sg13g2_decap_4 FILLER_41_731 ();
 sg13g2_fill_2 FILLER_41_735 ();
 sg13g2_fill_1 FILLER_41_747 ();
 sg13g2_fill_2 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_4 FILLER_42_63 ();
 sg13g2_fill_2 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_83 ();
 sg13g2_decap_4 FILLER_42_90 ();
 sg13g2_fill_2 FILLER_42_94 ();
 sg13g2_fill_2 FILLER_42_109 ();
 sg13g2_decap_8 FILLER_42_164 ();
 sg13g2_fill_1 FILLER_42_171 ();
 sg13g2_fill_1 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_282 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_decap_8 FILLER_42_320 ();
 sg13g2_fill_2 FILLER_42_327 ();
 sg13g2_decap_8 FILLER_42_337 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_fill_1 FILLER_42_346 ();
 sg13g2_decap_4 FILLER_42_386 ();
 sg13g2_decap_4 FILLER_42_413 ();
 sg13g2_fill_1 FILLER_42_417 ();
 sg13g2_fill_2 FILLER_42_422 ();
 sg13g2_decap_8 FILLER_42_458 ();
 sg13g2_fill_2 FILLER_42_465 ();
 sg13g2_fill_1 FILLER_42_467 ();
 sg13g2_decap_4 FILLER_42_480 ();
 sg13g2_fill_1 FILLER_42_507 ();
 sg13g2_decap_8 FILLER_42_517 ();
 sg13g2_fill_2 FILLER_42_524 ();
 sg13g2_fill_2 FILLER_42_535 ();
 sg13g2_fill_1 FILLER_42_537 ();
 sg13g2_fill_2 FILLER_42_549 ();
 sg13g2_fill_1 FILLER_42_551 ();
 sg13g2_decap_8 FILLER_42_565 ();
 sg13g2_decap_4 FILLER_42_580 ();
 sg13g2_fill_2 FILLER_42_584 ();
 sg13g2_decap_8 FILLER_42_607 ();
 sg13g2_decap_4 FILLER_42_614 ();
 sg13g2_decap_8 FILLER_42_627 ();
 sg13g2_fill_2 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_655 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_4 FILLER_42_669 ();
 sg13g2_fill_2 FILLER_42_673 ();
 sg13g2_fill_1 FILLER_42_680 ();
 sg13g2_decap_4 FILLER_42_699 ();
 sg13g2_fill_1 FILLER_42_703 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_fill_2 FILLER_42_727 ();
 sg13g2_fill_1 FILLER_42_729 ();
 sg13g2_fill_2 FILLER_42_744 ();
 sg13g2_fill_1 FILLER_42_746 ();
 sg13g2_decap_8 FILLER_42_779 ();
 sg13g2_decap_8 FILLER_42_786 ();
 sg13g2_decap_8 FILLER_42_793 ();
 sg13g2_decap_8 FILLER_42_800 ();
 sg13g2_decap_8 FILLER_42_807 ();
 sg13g2_decap_8 FILLER_42_814 ();
 sg13g2_decap_8 FILLER_42_821 ();
 sg13g2_decap_8 FILLER_42_828 ();
 sg13g2_decap_8 FILLER_42_835 ();
 sg13g2_decap_8 FILLER_42_842 ();
 sg13g2_decap_8 FILLER_42_849 ();
 sg13g2_decap_4 FILLER_42_856 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_4 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_67 ();
 sg13g2_decap_4 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_95 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_124 ();
 sg13g2_fill_1 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_4 FILLER_43_140 ();
 sg13g2_fill_1 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_166 ();
 sg13g2_fill_2 FILLER_43_212 ();
 sg13g2_fill_1 FILLER_43_214 ();
 sg13g2_decap_4 FILLER_43_264 ();
 sg13g2_decap_4 FILLER_43_295 ();
 sg13g2_fill_2 FILLER_43_322 ();
 sg13g2_decap_4 FILLER_43_341 ();
 sg13g2_fill_2 FILLER_43_345 ();
 sg13g2_decap_8 FILLER_43_355 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_369 ();
 sg13g2_fill_2 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_4 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_43_430 ();
 sg13g2_fill_1 FILLER_43_437 ();
 sg13g2_decap_4 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_456 ();
 sg13g2_decap_4 FILLER_43_463 ();
 sg13g2_fill_1 FILLER_43_467 ();
 sg13g2_fill_2 FILLER_43_477 ();
 sg13g2_fill_1 FILLER_43_479 ();
 sg13g2_fill_2 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_521 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_8 FILLER_43_544 ();
 sg13g2_decap_8 FILLER_43_557 ();
 sg13g2_decap_4 FILLER_43_564 ();
 sg13g2_fill_2 FILLER_43_568 ();
 sg13g2_decap_8 FILLER_43_586 ();
 sg13g2_decap_8 FILLER_43_593 ();
 sg13g2_fill_2 FILLER_43_614 ();
 sg13g2_fill_1 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_648 ();
 sg13g2_fill_2 FILLER_43_665 ();
 sg13g2_fill_2 FILLER_43_720 ();
 sg13g2_fill_1 FILLER_43_722 ();
 sg13g2_decap_4 FILLER_43_736 ();
 sg13g2_fill_1 FILLER_43_740 ();
 sg13g2_fill_2 FILLER_43_759 ();
 sg13g2_fill_1 FILLER_43_761 ();
 sg13g2_decap_8 FILLER_43_771 ();
 sg13g2_decap_8 FILLER_43_778 ();
 sg13g2_decap_8 FILLER_43_785 ();
 sg13g2_decap_8 FILLER_43_792 ();
 sg13g2_decap_8 FILLER_43_799 ();
 sg13g2_decap_8 FILLER_43_806 ();
 sg13g2_decap_8 FILLER_43_813 ();
 sg13g2_decap_8 FILLER_43_820 ();
 sg13g2_decap_8 FILLER_43_827 ();
 sg13g2_decap_8 FILLER_43_834 ();
 sg13g2_decap_8 FILLER_43_841 ();
 sg13g2_decap_8 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_855 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_fill_2 FILLER_44_21 ();
 sg13g2_fill_2 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_51 ();
 sg13g2_fill_1 FILLER_44_74 ();
 sg13g2_decap_8 FILLER_44_80 ();
 sg13g2_decap_8 FILLER_44_87 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_fill_2 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_122 ();
 sg13g2_decap_8 FILLER_44_129 ();
 sg13g2_decap_4 FILLER_44_136 ();
 sg13g2_decap_4 FILLER_44_156 ();
 sg13g2_decap_8 FILLER_44_180 ();
 sg13g2_decap_4 FILLER_44_187 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_201 ();
 sg13g2_decap_8 FILLER_44_208 ();
 sg13g2_decap_4 FILLER_44_219 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_fill_1 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_265 ();
 sg13g2_decap_8 FILLER_44_272 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_decap_4 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_302 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_decap_4 FILLER_44_340 ();
 sg13g2_decap_4 FILLER_44_368 ();
 sg13g2_fill_2 FILLER_44_372 ();
 sg13g2_decap_4 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_410 ();
 sg13g2_decap_8 FILLER_44_419 ();
 sg13g2_decap_8 FILLER_44_426 ();
 sg13g2_fill_2 FILLER_44_433 ();
 sg13g2_decap_8 FILLER_44_472 ();
 sg13g2_decap_8 FILLER_44_479 ();
 sg13g2_fill_1 FILLER_44_486 ();
 sg13g2_decap_8 FILLER_44_495 ();
 sg13g2_decap_4 FILLER_44_502 ();
 sg13g2_fill_2 FILLER_44_506 ();
 sg13g2_fill_2 FILLER_44_533 ();
 sg13g2_decap_4 FILLER_44_540 ();
 sg13g2_decap_4 FILLER_44_580 ();
 sg13g2_fill_1 FILLER_44_584 ();
 sg13g2_decap_8 FILLER_44_611 ();
 sg13g2_decap_8 FILLER_44_618 ();
 sg13g2_fill_2 FILLER_44_625 ();
 sg13g2_fill_1 FILLER_44_627 ();
 sg13g2_fill_2 FILLER_44_632 ();
 sg13g2_fill_1 FILLER_44_643 ();
 sg13g2_fill_2 FILLER_44_649 ();
 sg13g2_decap_4 FILLER_44_670 ();
 sg13g2_fill_1 FILLER_44_674 ();
 sg13g2_fill_2 FILLER_44_678 ();
 sg13g2_fill_1 FILLER_44_680 ();
 sg13g2_decap_4 FILLER_44_695 ();
 sg13g2_fill_1 FILLER_44_699 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_decap_8 FILLER_44_711 ();
 sg13g2_decap_8 FILLER_44_718 ();
 sg13g2_decap_4 FILLER_44_725 ();
 sg13g2_fill_2 FILLER_44_734 ();
 sg13g2_decap_8 FILLER_44_771 ();
 sg13g2_decap_8 FILLER_44_778 ();
 sg13g2_decap_8 FILLER_44_785 ();
 sg13g2_decap_8 FILLER_44_792 ();
 sg13g2_decap_8 FILLER_44_799 ();
 sg13g2_decap_8 FILLER_44_806 ();
 sg13g2_decap_8 FILLER_44_813 ();
 sg13g2_decap_8 FILLER_44_820 ();
 sg13g2_decap_8 FILLER_44_827 ();
 sg13g2_decap_8 FILLER_44_834 ();
 sg13g2_decap_8 FILLER_44_841 ();
 sg13g2_decap_8 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_855 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_fill_1 FILLER_45_18 ();
 sg13g2_fill_1 FILLER_45_28 ();
 sg13g2_fill_2 FILLER_45_38 ();
 sg13g2_fill_1 FILLER_45_40 ();
 sg13g2_decap_8 FILLER_45_50 ();
 sg13g2_fill_1 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_111 ();
 sg13g2_fill_1 FILLER_45_124 ();
 sg13g2_decap_8 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_143 ();
 sg13g2_fill_1 FILLER_45_145 ();
 sg13g2_fill_2 FILLER_45_160 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_decap_8 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_184 ();
 sg13g2_fill_2 FILLER_45_216 ();
 sg13g2_decap_4 FILLER_45_268 ();
 sg13g2_fill_2 FILLER_45_272 ();
 sg13g2_decap_8 FILLER_45_298 ();
 sg13g2_fill_2 FILLER_45_305 ();
 sg13g2_decap_8 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_362 ();
 sg13g2_fill_2 FILLER_45_369 ();
 sg13g2_fill_1 FILLER_45_371 ();
 sg13g2_decap_4 FILLER_45_393 ();
 sg13g2_fill_1 FILLER_45_406 ();
 sg13g2_decap_4 FILLER_45_456 ();
 sg13g2_fill_2 FILLER_45_480 ();
 sg13g2_decap_4 FILLER_45_490 ();
 sg13g2_fill_1 FILLER_45_494 ();
 sg13g2_decap_8 FILLER_45_524 ();
 sg13g2_fill_1 FILLER_45_531 ();
 sg13g2_decap_8 FILLER_45_551 ();
 sg13g2_fill_2 FILLER_45_571 ();
 sg13g2_decap_8 FILLER_45_577 ();
 sg13g2_decap_8 FILLER_45_584 ();
 sg13g2_fill_2 FILLER_45_591 ();
 sg13g2_fill_1 FILLER_45_688 ();
 sg13g2_decap_8 FILLER_45_699 ();
 sg13g2_fill_2 FILLER_45_706 ();
 sg13g2_fill_1 FILLER_45_708 ();
 sg13g2_decap_8 FILLER_45_743 ();
 sg13g2_decap_8 FILLER_45_750 ();
 sg13g2_decap_8 FILLER_45_757 ();
 sg13g2_decap_8 FILLER_45_764 ();
 sg13g2_decap_8 FILLER_45_771 ();
 sg13g2_decap_8 FILLER_45_778 ();
 sg13g2_decap_8 FILLER_45_785 ();
 sg13g2_decap_8 FILLER_45_792 ();
 sg13g2_decap_8 FILLER_45_799 ();
 sg13g2_decap_8 FILLER_45_806 ();
 sg13g2_decap_8 FILLER_45_813 ();
 sg13g2_decap_8 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_827 ();
 sg13g2_decap_8 FILLER_45_834 ();
 sg13g2_decap_8 FILLER_45_841 ();
 sg13g2_decap_8 FILLER_45_848 ();
 sg13g2_decap_8 FILLER_45_855 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_14 ();
 sg13g2_fill_2 FILLER_46_31 ();
 sg13g2_fill_2 FILLER_46_59 ();
 sg13g2_fill_1 FILLER_46_61 ();
 sg13g2_decap_8 FILLER_46_66 ();
 sg13g2_decap_4 FILLER_46_73 ();
 sg13g2_fill_1 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_82 ();
 sg13g2_decap_4 FILLER_46_89 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_4 FILLER_46_112 ();
 sg13g2_fill_2 FILLER_46_116 ();
 sg13g2_fill_2 FILLER_46_126 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_decap_4 FILLER_46_146 ();
 sg13g2_fill_1 FILLER_46_150 ();
 sg13g2_decap_8 FILLER_46_156 ();
 sg13g2_decap_4 FILLER_46_163 ();
 sg13g2_decap_4 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_240 ();
 sg13g2_decap_4 FILLER_46_247 ();
 sg13g2_decap_4 FILLER_46_272 ();
 sg13g2_fill_2 FILLER_46_276 ();
 sg13g2_fill_2 FILLER_46_290 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_decap_8 FILLER_46_316 ();
 sg13g2_fill_1 FILLER_46_323 ();
 sg13g2_decap_4 FILLER_46_340 ();
 sg13g2_fill_2 FILLER_46_344 ();
 sg13g2_decap_8 FILLER_46_411 ();
 sg13g2_fill_2 FILLER_46_418 ();
 sg13g2_decap_8 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_440 ();
 sg13g2_fill_1 FILLER_46_442 ();
 sg13g2_fill_2 FILLER_46_458 ();
 sg13g2_decap_8 FILLER_46_470 ();
 sg13g2_fill_1 FILLER_46_477 ();
 sg13g2_decap_8 FILLER_46_496 ();
 sg13g2_fill_2 FILLER_46_503 ();
 sg13g2_decap_8 FILLER_46_509 ();
 sg13g2_decap_8 FILLER_46_516 ();
 sg13g2_decap_8 FILLER_46_523 ();
 sg13g2_decap_8 FILLER_46_530 ();
 sg13g2_fill_1 FILLER_46_541 ();
 sg13g2_decap_8 FILLER_46_547 ();
 sg13g2_decap_4 FILLER_46_554 ();
 sg13g2_fill_1 FILLER_46_558 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_4 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_4 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_633 ();
 sg13g2_decap_8 FILLER_46_640 ();
 sg13g2_fill_1 FILLER_46_651 ();
 sg13g2_decap_4 FILLER_46_661 ();
 sg13g2_fill_2 FILLER_46_670 ();
 sg13g2_fill_1 FILLER_46_685 ();
 sg13g2_fill_1 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_734 ();
 sg13g2_decap_8 FILLER_46_741 ();
 sg13g2_decap_8 FILLER_46_748 ();
 sg13g2_decap_8 FILLER_46_755 ();
 sg13g2_decap_8 FILLER_46_762 ();
 sg13g2_decap_8 FILLER_46_769 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_decap_8 FILLER_46_783 ();
 sg13g2_decap_8 FILLER_46_790 ();
 sg13g2_decap_8 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_804 ();
 sg13g2_decap_8 FILLER_46_811 ();
 sg13g2_decap_8 FILLER_46_818 ();
 sg13g2_decap_8 FILLER_46_825 ();
 sg13g2_decap_8 FILLER_46_832 ();
 sg13g2_decap_8 FILLER_46_839 ();
 sg13g2_decap_8 FILLER_46_846 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_18 ();
 sg13g2_fill_2 FILLER_47_22 ();
 sg13g2_fill_1 FILLER_47_42 ();
 sg13g2_decap_4 FILLER_47_59 ();
 sg13g2_fill_2 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_78 ();
 sg13g2_decap_8 FILLER_47_108 ();
 sg13g2_decap_8 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_122 ();
 sg13g2_decap_4 FILLER_47_158 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_4 FILLER_47_189 ();
 sg13g2_fill_1 FILLER_47_193 ();
 sg13g2_decap_4 FILLER_47_217 ();
 sg13g2_decap_4 FILLER_47_227 ();
 sg13g2_fill_2 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_264 ();
 sg13g2_decap_8 FILLER_47_271 ();
 sg13g2_decap_4 FILLER_47_278 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_decap_8 FILLER_47_289 ();
 sg13g2_decap_4 FILLER_47_296 ();
 sg13g2_fill_1 FILLER_47_300 ();
 sg13g2_decap_8 FILLER_47_309 ();
 sg13g2_decap_8 FILLER_47_316 ();
 sg13g2_decap_8 FILLER_47_323 ();
 sg13g2_fill_2 FILLER_47_330 ();
 sg13g2_fill_1 FILLER_47_332 ();
 sg13g2_fill_2 FILLER_47_359 ();
 sg13g2_fill_1 FILLER_47_361 ();
 sg13g2_decap_8 FILLER_47_366 ();
 sg13g2_fill_2 FILLER_47_373 ();
 sg13g2_decap_4 FILLER_47_380 ();
 sg13g2_fill_2 FILLER_47_393 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_2 FILLER_47_421 ();
 sg13g2_fill_1 FILLER_47_423 ();
 sg13g2_decap_4 FILLER_47_427 ();
 sg13g2_fill_1 FILLER_47_431 ();
 sg13g2_decap_4 FILLER_47_444 ();
 sg13g2_fill_1 FILLER_47_448 ();
 sg13g2_decap_4 FILLER_47_454 ();
 sg13g2_fill_1 FILLER_47_458 ();
 sg13g2_fill_2 FILLER_47_464 ();
 sg13g2_fill_1 FILLER_47_480 ();
 sg13g2_decap_8 FILLER_47_486 ();
 sg13g2_decap_4 FILLER_47_493 ();
 sg13g2_fill_1 FILLER_47_497 ();
 sg13g2_fill_2 FILLER_47_511 ();
 sg13g2_fill_1 FILLER_47_513 ();
 sg13g2_fill_2 FILLER_47_555 ();
 sg13g2_fill_1 FILLER_47_557 ();
 sg13g2_fill_2 FILLER_47_563 ();
 sg13g2_decap_4 FILLER_47_570 ();
 sg13g2_fill_1 FILLER_47_574 ();
 sg13g2_decap_4 FILLER_47_584 ();
 sg13g2_fill_2 FILLER_47_620 ();
 sg13g2_fill_1 FILLER_47_622 ();
 sg13g2_decap_8 FILLER_47_654 ();
 sg13g2_fill_2 FILLER_47_661 ();
 sg13g2_fill_1 FILLER_47_663 ();
 sg13g2_fill_1 FILLER_47_680 ();
 sg13g2_fill_1 FILLER_47_686 ();
 sg13g2_fill_2 FILLER_47_695 ();
 sg13g2_fill_1 FILLER_47_697 ();
 sg13g2_fill_2 FILLER_47_703 ();
 sg13g2_fill_1 FILLER_47_705 ();
 sg13g2_fill_1 FILLER_47_719 ();
 sg13g2_decap_4 FILLER_47_727 ();
 sg13g2_decap_8 FILLER_47_744 ();
 sg13g2_decap_8 FILLER_47_751 ();
 sg13g2_decap_8 FILLER_47_758 ();
 sg13g2_decap_8 FILLER_47_765 ();
 sg13g2_decap_8 FILLER_47_772 ();
 sg13g2_decap_8 FILLER_47_779 ();
 sg13g2_decap_8 FILLER_47_786 ();
 sg13g2_decap_8 FILLER_47_793 ();
 sg13g2_decap_8 FILLER_47_800 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_decap_8 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_821 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_835 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_decap_4 FILLER_47_856 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_35 ();
 sg13g2_fill_2 FILLER_48_41 ();
 sg13g2_fill_1 FILLER_48_43 ();
 sg13g2_fill_1 FILLER_48_53 ();
 sg13g2_decap_8 FILLER_48_67 ();
 sg13g2_fill_1 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_88 ();
 sg13g2_fill_2 FILLER_48_93 ();
 sg13g2_fill_1 FILLER_48_118 ();
 sg13g2_decap_8 FILLER_48_131 ();
 sg13g2_decap_8 FILLER_48_138 ();
 sg13g2_decap_4 FILLER_48_145 ();
 sg13g2_fill_1 FILLER_48_149 ();
 sg13g2_decap_8 FILLER_48_158 ();
 sg13g2_decap_8 FILLER_48_178 ();
 sg13g2_fill_1 FILLER_48_185 ();
 sg13g2_decap_8 FILLER_48_220 ();
 sg13g2_fill_2 FILLER_48_227 ();
 sg13g2_decap_4 FILLER_48_250 ();
 sg13g2_fill_1 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_266 ();
 sg13g2_decap_4 FILLER_48_289 ();
 sg13g2_fill_2 FILLER_48_311 ();
 sg13g2_fill_1 FILLER_48_313 ();
 sg13g2_fill_2 FILLER_48_370 ();
 sg13g2_decap_4 FILLER_48_375 ();
 sg13g2_fill_1 FILLER_48_379 ();
 sg13g2_decap_4 FILLER_48_393 ();
 sg13g2_fill_1 FILLER_48_397 ();
 sg13g2_fill_2 FILLER_48_424 ();
 sg13g2_fill_1 FILLER_48_426 ();
 sg13g2_decap_4 FILLER_48_441 ();
 sg13g2_fill_1 FILLER_48_445 ();
 sg13g2_decap_4 FILLER_48_454 ();
 sg13g2_fill_1 FILLER_48_458 ();
 sg13g2_fill_2 FILLER_48_493 ();
 sg13g2_fill_1 FILLER_48_495 ();
 sg13g2_decap_8 FILLER_48_516 ();
 sg13g2_fill_2 FILLER_48_523 ();
 sg13g2_fill_2 FILLER_48_529 ();
 sg13g2_fill_1 FILLER_48_540 ();
 sg13g2_fill_2 FILLER_48_560 ();
 sg13g2_fill_1 FILLER_48_562 ();
 sg13g2_decap_4 FILLER_48_592 ();
 sg13g2_fill_1 FILLER_48_596 ();
 sg13g2_fill_2 FILLER_48_601 ();
 sg13g2_fill_1 FILLER_48_603 ();
 sg13g2_decap_8 FILLER_48_625 ();
 sg13g2_fill_2 FILLER_48_632 ();
 sg13g2_fill_1 FILLER_48_638 ();
 sg13g2_decap_4 FILLER_48_656 ();
 sg13g2_fill_2 FILLER_48_660 ();
 sg13g2_fill_1 FILLER_48_670 ();
 sg13g2_fill_1 FILLER_48_689 ();
 sg13g2_decap_4 FILLER_48_703 ();
 sg13g2_fill_1 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_747 ();
 sg13g2_decap_8 FILLER_48_754 ();
 sg13g2_decap_8 FILLER_48_761 ();
 sg13g2_decap_8 FILLER_48_768 ();
 sg13g2_decap_8 FILLER_48_775 ();
 sg13g2_decap_8 FILLER_48_782 ();
 sg13g2_decap_8 FILLER_48_789 ();
 sg13g2_decap_8 FILLER_48_796 ();
 sg13g2_decap_8 FILLER_48_803 ();
 sg13g2_decap_8 FILLER_48_810 ();
 sg13g2_decap_8 FILLER_48_817 ();
 sg13g2_decap_8 FILLER_48_824 ();
 sg13g2_decap_8 FILLER_48_831 ();
 sg13g2_decap_8 FILLER_48_838 ();
 sg13g2_decap_8 FILLER_48_845 ();
 sg13g2_decap_8 FILLER_48_852 ();
 sg13g2_fill_2 FILLER_48_859 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_fill_2 FILLER_49_48 ();
 sg13g2_fill_1 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_55 ();
 sg13g2_decap_8 FILLER_49_69 ();
 sg13g2_decap_4 FILLER_49_76 ();
 sg13g2_decap_8 FILLER_49_83 ();
 sg13g2_decap_8 FILLER_49_90 ();
 sg13g2_fill_2 FILLER_49_97 ();
 sg13g2_decap_8 FILLER_49_107 ();
 sg13g2_fill_2 FILLER_49_114 ();
 sg13g2_fill_2 FILLER_49_121 ();
 sg13g2_fill_2 FILLER_49_127 ();
 sg13g2_decap_8 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_decap_4 FILLER_49_150 ();
 sg13g2_fill_2 FILLER_49_154 ();
 sg13g2_fill_2 FILLER_49_188 ();
 sg13g2_decap_8 FILLER_49_211 ();
 sg13g2_decap_4 FILLER_49_218 ();
 sg13g2_fill_1 FILLER_49_222 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_248 ();
 sg13g2_fill_2 FILLER_49_255 ();
 sg13g2_decap_8 FILLER_49_281 ();
 sg13g2_decap_8 FILLER_49_288 ();
 sg13g2_fill_2 FILLER_49_299 ();
 sg13g2_fill_1 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_decap_4 FILLER_49_324 ();
 sg13g2_fill_2 FILLER_49_376 ();
 sg13g2_fill_1 FILLER_49_378 ();
 sg13g2_fill_1 FILLER_49_384 ();
 sg13g2_decap_4 FILLER_49_398 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_4 FILLER_49_425 ();
 sg13g2_fill_1 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_449 ();
 sg13g2_fill_2 FILLER_49_456 ();
 sg13g2_fill_1 FILLER_49_458 ();
 sg13g2_decap_8 FILLER_49_472 ();
 sg13g2_fill_2 FILLER_49_479 ();
 sg13g2_decap_8 FILLER_49_493 ();
 sg13g2_decap_8 FILLER_49_500 ();
 sg13g2_fill_2 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_fill_2 FILLER_49_539 ();
 sg13g2_fill_2 FILLER_49_552 ();
 sg13g2_fill_1 FILLER_49_554 ();
 sg13g2_decap_4 FILLER_49_563 ();
 sg13g2_decap_8 FILLER_49_572 ();
 sg13g2_decap_8 FILLER_49_579 ();
 sg13g2_fill_1 FILLER_49_586 ();
 sg13g2_decap_8 FILLER_49_605 ();
 sg13g2_decap_8 FILLER_49_617 ();
 sg13g2_decap_8 FILLER_49_624 ();
 sg13g2_decap_4 FILLER_49_631 ();
 sg13g2_decap_8 FILLER_49_643 ();
 sg13g2_decap_8 FILLER_49_650 ();
 sg13g2_decap_8 FILLER_49_657 ();
 sg13g2_decap_4 FILLER_49_664 ();
 sg13g2_fill_2 FILLER_49_668 ();
 sg13g2_fill_2 FILLER_49_678 ();
 sg13g2_fill_1 FILLER_49_680 ();
 sg13g2_decap_4 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_698 ();
 sg13g2_fill_2 FILLER_49_705 ();
 sg13g2_decap_8 FILLER_49_719 ();
 sg13g2_decap_8 FILLER_49_726 ();
 sg13g2_decap_8 FILLER_49_733 ();
 sg13g2_decap_8 FILLER_49_740 ();
 sg13g2_decap_8 FILLER_49_747 ();
 sg13g2_decap_8 FILLER_49_754 ();
 sg13g2_decap_8 FILLER_49_761 ();
 sg13g2_decap_8 FILLER_49_768 ();
 sg13g2_decap_8 FILLER_49_775 ();
 sg13g2_decap_8 FILLER_49_782 ();
 sg13g2_decap_8 FILLER_49_789 ();
 sg13g2_decap_8 FILLER_49_796 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_810 ();
 sg13g2_decap_8 FILLER_49_817 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_decap_8 FILLER_49_838 ();
 sg13g2_decap_8 FILLER_49_845 ();
 sg13g2_decap_8 FILLER_49_852 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_fill_1 FILLER_50_26 ();
 sg13g2_fill_2 FILLER_50_46 ();
 sg13g2_fill_1 FILLER_50_65 ();
 sg13g2_fill_2 FILLER_50_84 ();
 sg13g2_decap_4 FILLER_50_103 ();
 sg13g2_fill_1 FILLER_50_107 ();
 sg13g2_decap_8 FILLER_50_120 ();
 sg13g2_fill_1 FILLER_50_127 ();
 sg13g2_decap_8 FILLER_50_150 ();
 sg13g2_decap_4 FILLER_50_161 ();
 sg13g2_fill_1 FILLER_50_165 ();
 sg13g2_fill_2 FILLER_50_180 ();
 sg13g2_fill_2 FILLER_50_196 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_decap_4 FILLER_50_233 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_263 ();
 sg13g2_fill_1 FILLER_50_290 ();
 sg13g2_decap_8 FILLER_50_304 ();
 sg13g2_decap_4 FILLER_50_311 ();
 sg13g2_fill_2 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_372 ();
 sg13g2_decap_8 FILLER_50_379 ();
 sg13g2_decap_4 FILLER_50_386 ();
 sg13g2_fill_2 FILLER_50_390 ();
 sg13g2_fill_2 FILLER_50_426 ();
 sg13g2_fill_1 FILLER_50_428 ();
 sg13g2_fill_1 FILLER_50_454 ();
 sg13g2_fill_2 FILLER_50_482 ();
 sg13g2_fill_2 FILLER_50_505 ();
 sg13g2_fill_1 FILLER_50_507 ();
 sg13g2_decap_4 FILLER_50_529 ();
 sg13g2_fill_1 FILLER_50_533 ();
 sg13g2_fill_1 FILLER_50_553 ();
 sg13g2_fill_2 FILLER_50_604 ();
 sg13g2_fill_2 FILLER_50_614 ();
 sg13g2_fill_1 FILLER_50_616 ();
 sg13g2_fill_2 FILLER_50_625 ();
 sg13g2_fill_1 FILLER_50_627 ();
 sg13g2_decap_8 FILLER_50_645 ();
 sg13g2_decap_8 FILLER_50_652 ();
 sg13g2_decap_4 FILLER_50_672 ();
 sg13g2_decap_4 FILLER_50_688 ();
 sg13g2_fill_1 FILLER_50_692 ();
 sg13g2_decap_4 FILLER_50_722 ();
 sg13g2_fill_1 FILLER_50_726 ();
 sg13g2_decap_8 FILLER_50_737 ();
 sg13g2_decap_8 FILLER_50_744 ();
 sg13g2_decap_8 FILLER_50_751 ();
 sg13g2_decap_8 FILLER_50_758 ();
 sg13g2_decap_8 FILLER_50_765 ();
 sg13g2_decap_8 FILLER_50_772 ();
 sg13g2_decap_8 FILLER_50_779 ();
 sg13g2_decap_8 FILLER_50_786 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_decap_8 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_807 ();
 sg13g2_decap_8 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_821 ();
 sg13g2_decap_8 FILLER_50_828 ();
 sg13g2_decap_8 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_842 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_11 ();
 sg13g2_decap_8 FILLER_51_53 ();
 sg13g2_decap_4 FILLER_51_60 ();
 sg13g2_fill_1 FILLER_51_64 ();
 sg13g2_decap_4 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_86 ();
 sg13g2_decap_8 FILLER_51_92 ();
 sg13g2_decap_8 FILLER_51_99 ();
 sg13g2_decap_4 FILLER_51_106 ();
 sg13g2_decap_4 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_157 ();
 sg13g2_fill_2 FILLER_51_203 ();
 sg13g2_fill_1 FILLER_51_205 ();
 sg13g2_decap_4 FILLER_51_219 ();
 sg13g2_fill_2 FILLER_51_223 ();
 sg13g2_fill_2 FILLER_51_234 ();
 sg13g2_fill_1 FILLER_51_236 ();
 sg13g2_decap_4 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_274 ();
 sg13g2_fill_2 FILLER_51_287 ();
 sg13g2_fill_1 FILLER_51_289 ();
 sg13g2_decap_8 FILLER_51_302 ();
 sg13g2_fill_2 FILLER_51_309 ();
 sg13g2_fill_1 FILLER_51_311 ();
 sg13g2_fill_1 FILLER_51_316 ();
 sg13g2_decap_4 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_362 ();
 sg13g2_fill_2 FILLER_51_368 ();
 sg13g2_fill_2 FILLER_51_375 ();
 sg13g2_fill_1 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_397 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_2 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_51_415 ();
 sg13g2_decap_8 FILLER_51_422 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_8 FILLER_51_439 ();
 sg13g2_decap_8 FILLER_51_446 ();
 sg13g2_decap_8 FILLER_51_453 ();
 sg13g2_decap_4 FILLER_51_460 ();
 sg13g2_decap_8 FILLER_51_472 ();
 sg13g2_decap_4 FILLER_51_479 ();
 sg13g2_decap_8 FILLER_51_500 ();
 sg13g2_decap_8 FILLER_51_507 ();
 sg13g2_fill_1 FILLER_51_514 ();
 sg13g2_decap_8 FILLER_51_529 ();
 sg13g2_decap_8 FILLER_51_536 ();
 sg13g2_fill_1 FILLER_51_557 ();
 sg13g2_decap_8 FILLER_51_574 ();
 sg13g2_decap_8 FILLER_51_581 ();
 sg13g2_fill_1 FILLER_51_588 ();
 sg13g2_decap_4 FILLER_51_608 ();
 sg13g2_fill_2 FILLER_51_617 ();
 sg13g2_fill_1 FILLER_51_628 ();
 sg13g2_fill_2 FILLER_51_645 ();
 sg13g2_fill_1 FILLER_51_647 ();
 sg13g2_fill_1 FILLER_51_665 ();
 sg13g2_decap_8 FILLER_51_683 ();
 sg13g2_fill_1 FILLER_51_690 ();
 sg13g2_decap_8 FILLER_51_700 ();
 sg13g2_fill_2 FILLER_51_707 ();
 sg13g2_fill_2 FILLER_51_714 ();
 sg13g2_fill_1 FILLER_51_721 ();
 sg13g2_fill_1 FILLER_51_730 ();
 sg13g2_decap_8 FILLER_51_762 ();
 sg13g2_decap_8 FILLER_51_769 ();
 sg13g2_decap_8 FILLER_51_776 ();
 sg13g2_decap_8 FILLER_51_783 ();
 sg13g2_decap_8 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_797 ();
 sg13g2_decap_8 FILLER_51_804 ();
 sg13g2_decap_8 FILLER_51_811 ();
 sg13g2_decap_8 FILLER_51_818 ();
 sg13g2_decap_8 FILLER_51_825 ();
 sg13g2_decap_8 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_839 ();
 sg13g2_decap_8 FILLER_51_846 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_15 ();
 sg13g2_fill_1 FILLER_52_22 ();
 sg13g2_fill_2 FILLER_52_31 ();
 sg13g2_fill_2 FILLER_52_41 ();
 sg13g2_fill_1 FILLER_52_47 ();
 sg13g2_decap_4 FILLER_52_58 ();
 sg13g2_fill_1 FILLER_52_78 ();
 sg13g2_decap_4 FILLER_52_97 ();
 sg13g2_fill_1 FILLER_52_101 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_4 FILLER_52_140 ();
 sg13g2_fill_1 FILLER_52_163 ();
 sg13g2_decap_8 FILLER_52_256 ();
 sg13g2_decap_4 FILLER_52_263 ();
 sg13g2_fill_1 FILLER_52_267 ();
 sg13g2_decap_8 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_279 ();
 sg13g2_decap_8 FILLER_52_290 ();
 sg13g2_decap_4 FILLER_52_297 ();
 sg13g2_fill_2 FILLER_52_327 ();
 sg13g2_fill_1 FILLER_52_329 ();
 sg13g2_decap_4 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_370 ();
 sg13g2_fill_2 FILLER_52_377 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_fill_2 FILLER_52_391 ();
 sg13g2_fill_1 FILLER_52_393 ();
 sg13g2_decap_4 FILLER_52_398 ();
 sg13g2_fill_2 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_52_418 ();
 sg13g2_decap_8 FILLER_52_425 ();
 sg13g2_fill_2 FILLER_52_432 ();
 sg13g2_decap_4 FILLER_52_439 ();
 sg13g2_fill_2 FILLER_52_451 ();
 sg13g2_decap_8 FILLER_52_458 ();
 sg13g2_decap_8 FILLER_52_465 ();
 sg13g2_fill_2 FILLER_52_480 ();
 sg13g2_fill_1 FILLER_52_482 ();
 sg13g2_decap_8 FILLER_52_494 ();
 sg13g2_decap_4 FILLER_52_507 ();
 sg13g2_fill_1 FILLER_52_511 ();
 sg13g2_decap_8 FILLER_52_530 ();
 sg13g2_fill_2 FILLER_52_537 ();
 sg13g2_fill_1 FILLER_52_544 ();
 sg13g2_fill_1 FILLER_52_549 ();
 sg13g2_fill_1 FILLER_52_559 ();
 sg13g2_fill_2 FILLER_52_575 ();
 sg13g2_fill_1 FILLER_52_577 ();
 sg13g2_fill_2 FILLER_52_599 ();
 sg13g2_fill_2 FILLER_52_619 ();
 sg13g2_fill_1 FILLER_52_621 ();
 sg13g2_decap_4 FILLER_52_626 ();
 sg13g2_decap_8 FILLER_52_638 ();
 sg13g2_fill_2 FILLER_52_645 ();
 sg13g2_decap_4 FILLER_52_658 ();
 sg13g2_decap_4 FILLER_52_670 ();
 sg13g2_fill_2 FILLER_52_674 ();
 sg13g2_fill_2 FILLER_52_689 ();
 sg13g2_fill_1 FILLER_52_717 ();
 sg13g2_fill_1 FILLER_52_746 ();
 sg13g2_decap_8 FILLER_52_751 ();
 sg13g2_decap_8 FILLER_52_758 ();
 sg13g2_decap_8 FILLER_52_765 ();
 sg13g2_decap_8 FILLER_52_772 ();
 sg13g2_decap_8 FILLER_52_779 ();
 sg13g2_decap_8 FILLER_52_786 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_decap_8 FILLER_52_800 ();
 sg13g2_decap_8 FILLER_52_807 ();
 sg13g2_decap_8 FILLER_52_814 ();
 sg13g2_decap_8 FILLER_52_821 ();
 sg13g2_decap_8 FILLER_52_828 ();
 sg13g2_decap_8 FILLER_52_835 ();
 sg13g2_decap_8 FILLER_52_842 ();
 sg13g2_decap_8 FILLER_52_849 ();
 sg13g2_decap_4 FILLER_52_856 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_37 ();
 sg13g2_fill_2 FILLER_53_41 ();
 sg13g2_decap_8 FILLER_53_61 ();
 sg13g2_decap_8 FILLER_53_68 ();
 sg13g2_fill_2 FILLER_53_75 ();
 sg13g2_fill_2 FILLER_53_82 ();
 sg13g2_fill_1 FILLER_53_84 ();
 sg13g2_decap_4 FILLER_53_90 ();
 sg13g2_decap_8 FILLER_53_99 ();
 sg13g2_decap_4 FILLER_53_106 ();
 sg13g2_fill_2 FILLER_53_110 ();
 sg13g2_decap_4 FILLER_53_121 ();
 sg13g2_decap_8 FILLER_53_138 ();
 sg13g2_decap_4 FILLER_53_145 ();
 sg13g2_fill_2 FILLER_53_149 ();
 sg13g2_fill_1 FILLER_53_155 ();
 sg13g2_fill_2 FILLER_53_170 ();
 sg13g2_fill_1 FILLER_53_172 ();
 sg13g2_fill_1 FILLER_53_199 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_224 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_293 ();
 sg13g2_fill_1 FILLER_53_315 ();
 sg13g2_fill_2 FILLER_53_343 ();
 sg13g2_fill_1 FILLER_53_345 ();
 sg13g2_fill_2 FILLER_53_351 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_360 ();
 sg13g2_fill_1 FILLER_53_362 ();
 sg13g2_decap_4 FILLER_53_389 ();
 sg13g2_fill_1 FILLER_53_407 ();
 sg13g2_fill_2 FILLER_53_442 ();
 sg13g2_decap_4 FILLER_53_468 ();
 sg13g2_fill_1 FILLER_53_483 ();
 sg13g2_decap_8 FILLER_53_500 ();
 sg13g2_fill_2 FILLER_53_507 ();
 sg13g2_fill_1 FILLER_53_607 ();
 sg13g2_fill_2 FILLER_53_632 ();
 sg13g2_fill_1 FILLER_53_634 ();
 sg13g2_fill_2 FILLER_53_640 ();
 sg13g2_fill_1 FILLER_53_642 ();
 sg13g2_decap_8 FILLER_53_648 ();
 sg13g2_decap_4 FILLER_53_655 ();
 sg13g2_decap_8 FILLER_53_679 ();
 sg13g2_fill_1 FILLER_53_686 ();
 sg13g2_decap_8 FILLER_53_692 ();
 sg13g2_decap_8 FILLER_53_713 ();
 sg13g2_decap_8 FILLER_53_720 ();
 sg13g2_decap_4 FILLER_53_727 ();
 sg13g2_fill_1 FILLER_53_731 ();
 sg13g2_fill_2 FILLER_53_735 ();
 sg13g2_fill_1 FILLER_53_737 ();
 sg13g2_decap_8 FILLER_53_764 ();
 sg13g2_decap_8 FILLER_53_771 ();
 sg13g2_decap_8 FILLER_53_778 ();
 sg13g2_decap_8 FILLER_53_785 ();
 sg13g2_decap_8 FILLER_53_792 ();
 sg13g2_decap_8 FILLER_53_799 ();
 sg13g2_decap_8 FILLER_53_806 ();
 sg13g2_decap_8 FILLER_53_813 ();
 sg13g2_decap_8 FILLER_53_820 ();
 sg13g2_decap_8 FILLER_53_827 ();
 sg13g2_decap_8 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_841 ();
 sg13g2_decap_8 FILLER_53_848 ();
 sg13g2_decap_8 FILLER_53_855 ();
 sg13g2_fill_2 FILLER_54_26 ();
 sg13g2_fill_1 FILLER_54_48 ();
 sg13g2_decap_8 FILLER_54_66 ();
 sg13g2_fill_1 FILLER_54_73 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_106 ();
 sg13g2_fill_2 FILLER_54_115 ();
 sg13g2_fill_1 FILLER_54_117 ();
 sg13g2_decap_4 FILLER_54_135 ();
 sg13g2_fill_2 FILLER_54_147 ();
 sg13g2_fill_1 FILLER_54_149 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_fill_1 FILLER_54_164 ();
 sg13g2_decap_4 FILLER_54_169 ();
 sg13g2_fill_2 FILLER_54_173 ();
 sg13g2_decap_4 FILLER_54_233 ();
 sg13g2_decap_8 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_249 ();
 sg13g2_fill_2 FILLER_54_257 ();
 sg13g2_decap_8 FILLER_54_264 ();
 sg13g2_decap_8 FILLER_54_271 ();
 sg13g2_decap_4 FILLER_54_278 ();
 sg13g2_decap_4 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_294 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_decap_4 FILLER_54_315 ();
 sg13g2_decap_4 FILLER_54_323 ();
 sg13g2_fill_2 FILLER_54_327 ();
 sg13g2_decap_8 FILLER_54_334 ();
 sg13g2_fill_1 FILLER_54_341 ();
 sg13g2_fill_2 FILLER_54_351 ();
 sg13g2_fill_2 FILLER_54_394 ();
 sg13g2_fill_1 FILLER_54_396 ();
 sg13g2_fill_1 FILLER_54_405 ();
 sg13g2_decap_8 FILLER_54_410 ();
 sg13g2_fill_2 FILLER_54_422 ();
 sg13g2_decap_8 FILLER_54_446 ();
 sg13g2_decap_8 FILLER_54_453 ();
 sg13g2_fill_1 FILLER_54_460 ();
 sg13g2_decap_8 FILLER_54_466 ();
 sg13g2_decap_8 FILLER_54_473 ();
 sg13g2_decap_8 FILLER_54_480 ();
 sg13g2_decap_8 FILLER_54_498 ();
 sg13g2_decap_8 FILLER_54_505 ();
 sg13g2_decap_8 FILLER_54_524 ();
 sg13g2_decap_8 FILLER_54_531 ();
 sg13g2_fill_1 FILLER_54_538 ();
 sg13g2_decap_4 FILLER_54_551 ();
 sg13g2_decap_4 FILLER_54_570 ();
 sg13g2_fill_1 FILLER_54_574 ();
 sg13g2_decap_8 FILLER_54_579 ();
 sg13g2_fill_2 FILLER_54_586 ();
 sg13g2_fill_2 FILLER_54_610 ();
 sg13g2_fill_2 FILLER_54_626 ();
 sg13g2_decap_8 FILLER_54_650 ();
 sg13g2_fill_1 FILLER_54_657 ();
 sg13g2_decap_8 FILLER_54_675 ();
 sg13g2_fill_2 FILLER_54_682 ();
 sg13g2_fill_1 FILLER_54_684 ();
 sg13g2_fill_2 FILLER_54_704 ();
 sg13g2_decap_8 FILLER_54_755 ();
 sg13g2_decap_8 FILLER_54_762 ();
 sg13g2_decap_8 FILLER_54_769 ();
 sg13g2_decap_8 FILLER_54_776 ();
 sg13g2_decap_8 FILLER_54_783 ();
 sg13g2_decap_8 FILLER_54_790 ();
 sg13g2_decap_8 FILLER_54_797 ();
 sg13g2_decap_8 FILLER_54_804 ();
 sg13g2_decap_8 FILLER_54_811 ();
 sg13g2_decap_8 FILLER_54_818 ();
 sg13g2_decap_8 FILLER_54_825 ();
 sg13g2_decap_8 FILLER_54_832 ();
 sg13g2_decap_8 FILLER_54_839 ();
 sg13g2_decap_8 FILLER_54_846 ();
 sg13g2_decap_8 FILLER_54_853 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_27 ();
 sg13g2_fill_1 FILLER_55_35 ();
 sg13g2_fill_1 FILLER_55_48 ();
 sg13g2_fill_2 FILLER_55_54 ();
 sg13g2_decap_4 FILLER_55_60 ();
 sg13g2_fill_1 FILLER_55_64 ();
 sg13g2_decap_8 FILLER_55_73 ();
 sg13g2_decap_8 FILLER_55_80 ();
 sg13g2_decap_4 FILLER_55_87 ();
 sg13g2_fill_2 FILLER_55_96 ();
 sg13g2_fill_2 FILLER_55_103 ();
 sg13g2_decap_8 FILLER_55_110 ();
 sg13g2_decap_4 FILLER_55_117 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_fill_1 FILLER_55_131 ();
 sg13g2_fill_2 FILLER_55_137 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_2 FILLER_55_157 ();
 sg13g2_decap_8 FILLER_55_181 ();
 sg13g2_decap_4 FILLER_55_188 ();
 sg13g2_fill_1 FILLER_55_192 ();
 sg13g2_decap_8 FILLER_55_206 ();
 sg13g2_decap_8 FILLER_55_213 ();
 sg13g2_decap_8 FILLER_55_220 ();
 sg13g2_decap_8 FILLER_55_227 ();
 sg13g2_decap_8 FILLER_55_234 ();
 sg13g2_fill_2 FILLER_55_254 ();
 sg13g2_fill_2 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_344 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_fill_1 FILLER_55_404 ();
 sg13g2_decap_4 FILLER_55_477 ();
 sg13g2_fill_1 FILLER_55_481 ();
 sg13g2_decap_8 FILLER_55_499 ();
 sg13g2_fill_2 FILLER_55_506 ();
 sg13g2_decap_4 FILLER_55_529 ();
 sg13g2_fill_2 FILLER_55_533 ();
 sg13g2_fill_1 FILLER_55_561 ();
 sg13g2_fill_2 FILLER_55_600 ();
 sg13g2_decap_8 FILLER_55_628 ();
 sg13g2_fill_2 FILLER_55_651 ();
 sg13g2_decap_8 FILLER_55_661 ();
 sg13g2_decap_8 FILLER_55_668 ();
 sg13g2_decap_8 FILLER_55_675 ();
 sg13g2_fill_1 FILLER_55_694 ();
 sg13g2_decap_8 FILLER_55_708 ();
 sg13g2_decap_8 FILLER_55_715 ();
 sg13g2_decap_4 FILLER_55_722 ();
 sg13g2_fill_1 FILLER_55_726 ();
 sg13g2_fill_2 FILLER_55_740 ();
 sg13g2_decap_8 FILLER_55_755 ();
 sg13g2_decap_8 FILLER_55_762 ();
 sg13g2_decap_8 FILLER_55_769 ();
 sg13g2_decap_8 FILLER_55_776 ();
 sg13g2_decap_8 FILLER_55_783 ();
 sg13g2_decap_8 FILLER_55_790 ();
 sg13g2_decap_8 FILLER_55_797 ();
 sg13g2_decap_8 FILLER_55_804 ();
 sg13g2_decap_8 FILLER_55_811 ();
 sg13g2_decap_8 FILLER_55_818 ();
 sg13g2_decap_8 FILLER_55_825 ();
 sg13g2_decap_8 FILLER_55_832 ();
 sg13g2_decap_8 FILLER_55_839 ();
 sg13g2_decap_8 FILLER_55_846 ();
 sg13g2_decap_8 FILLER_55_853 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_fill_2 FILLER_56_26 ();
 sg13g2_decap_8 FILLER_56_40 ();
 sg13g2_decap_4 FILLER_56_47 ();
 sg13g2_decap_4 FILLER_56_85 ();
 sg13g2_fill_2 FILLER_56_97 ();
 sg13g2_fill_1 FILLER_56_104 ();
 sg13g2_fill_1 FILLER_56_118 ();
 sg13g2_decap_8 FILLER_56_127 ();
 sg13g2_fill_1 FILLER_56_142 ();
 sg13g2_decap_8 FILLER_56_146 ();
 sg13g2_decap_8 FILLER_56_153 ();
 sg13g2_fill_2 FILLER_56_160 ();
 sg13g2_decap_4 FILLER_56_202 ();
 sg13g2_fill_2 FILLER_56_220 ();
 sg13g2_decap_8 FILLER_56_261 ();
 sg13g2_decap_8 FILLER_56_268 ();
 sg13g2_decap_4 FILLER_56_275 ();
 sg13g2_fill_1 FILLER_56_279 ();
 sg13g2_fill_1 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_302 ();
 sg13g2_decap_8 FILLER_56_308 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_decap_4 FILLER_56_329 ();
 sg13g2_fill_1 FILLER_56_348 ();
 sg13g2_fill_2 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_423 ();
 sg13g2_decap_8 FILLER_56_439 ();
 sg13g2_decap_8 FILLER_56_446 ();
 sg13g2_decap_8 FILLER_56_453 ();
 sg13g2_decap_4 FILLER_56_460 ();
 sg13g2_decap_8 FILLER_56_478 ();
 sg13g2_decap_4 FILLER_56_501 ();
 sg13g2_fill_2 FILLER_56_505 ();
 sg13g2_decap_4 FILLER_56_529 ();
 sg13g2_fill_1 FILLER_56_533 ();
 sg13g2_fill_2 FILLER_56_544 ();
 sg13g2_fill_1 FILLER_56_550 ();
 sg13g2_decap_8 FILLER_56_564 ();
 sg13g2_decap_4 FILLER_56_571 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_decap_8 FILLER_56_580 ();
 sg13g2_decap_4 FILLER_56_587 ();
 sg13g2_fill_2 FILLER_56_611 ();
 sg13g2_decap_8 FILLER_56_630 ();
 sg13g2_decap_4 FILLER_56_637 ();
 sg13g2_fill_1 FILLER_56_641 ();
 sg13g2_fill_2 FILLER_56_652 ();
 sg13g2_fill_1 FILLER_56_654 ();
 sg13g2_decap_8 FILLER_56_672 ();
 sg13g2_fill_2 FILLER_56_679 ();
 sg13g2_fill_1 FILLER_56_681 ();
 sg13g2_decap_8 FILLER_56_686 ();
 sg13g2_decap_8 FILLER_56_693 ();
 sg13g2_decap_4 FILLER_56_700 ();
 sg13g2_fill_2 FILLER_56_721 ();
 sg13g2_decap_8 FILLER_56_728 ();
 sg13g2_fill_2 FILLER_56_735 ();
 sg13g2_fill_2 FILLER_56_740 ();
 sg13g2_fill_1 FILLER_56_742 ();
 sg13g2_decap_8 FILLER_56_769 ();
 sg13g2_decap_8 FILLER_56_776 ();
 sg13g2_decap_8 FILLER_56_783 ();
 sg13g2_decap_8 FILLER_56_790 ();
 sg13g2_decap_8 FILLER_56_797 ();
 sg13g2_decap_8 FILLER_56_804 ();
 sg13g2_decap_8 FILLER_56_811 ();
 sg13g2_decap_8 FILLER_56_818 ();
 sg13g2_decap_8 FILLER_56_825 ();
 sg13g2_decap_8 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_839 ();
 sg13g2_decap_8 FILLER_56_846 ();
 sg13g2_decap_8 FILLER_56_853 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_15 ();
 sg13g2_fill_1 FILLER_57_27 ();
 sg13g2_decap_4 FILLER_57_58 ();
 sg13g2_fill_2 FILLER_57_62 ();
 sg13g2_decap_4 FILLER_57_68 ();
 sg13g2_fill_2 FILLER_57_72 ();
 sg13g2_decap_4 FILLER_57_80 ();
 sg13g2_decap_8 FILLER_57_89 ();
 sg13g2_fill_2 FILLER_57_96 ();
 sg13g2_decap_8 FILLER_57_103 ();
 sg13g2_decap_8 FILLER_57_110 ();
 sg13g2_decap_8 FILLER_57_117 ();
 sg13g2_decap_8 FILLER_57_124 ();
 sg13g2_decap_4 FILLER_57_131 ();
 sg13g2_fill_2 FILLER_57_152 ();
 sg13g2_fill_1 FILLER_57_154 ();
 sg13g2_decap_4 FILLER_57_164 ();
 sg13g2_fill_1 FILLER_57_168 ();
 sg13g2_fill_2 FILLER_57_178 ();
 sg13g2_fill_1 FILLER_57_180 ();
 sg13g2_decap_8 FILLER_57_186 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_fill_2 FILLER_57_255 ();
 sg13g2_decap_8 FILLER_57_275 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_fill_2 FILLER_57_307 ();
 sg13g2_fill_1 FILLER_57_309 ();
 sg13g2_fill_2 FILLER_57_320 ();
 sg13g2_decap_8 FILLER_57_327 ();
 sg13g2_decap_4 FILLER_57_334 ();
 sg13g2_fill_2 FILLER_57_338 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_2 FILLER_57_366 ();
 sg13g2_fill_1 FILLER_57_382 ();
 sg13g2_fill_2 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_410 ();
 sg13g2_fill_1 FILLER_57_425 ();
 sg13g2_decap_4 FILLER_57_460 ();
 sg13g2_decap_8 FILLER_57_474 ();
 sg13g2_decap_8 FILLER_57_481 ();
 sg13g2_decap_4 FILLER_57_503 ();
 sg13g2_fill_2 FILLER_57_507 ();
 sg13g2_decap_8 FILLER_57_532 ();
 sg13g2_fill_2 FILLER_57_539 ();
 sg13g2_fill_1 FILLER_57_541 ();
 sg13g2_fill_2 FILLER_57_568 ();
 sg13g2_fill_1 FILLER_57_570 ();
 sg13g2_fill_1 FILLER_57_606 ();
 sg13g2_fill_1 FILLER_57_641 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_fill_2 FILLER_57_668 ();
 sg13g2_fill_1 FILLER_57_670 ();
 sg13g2_decap_8 FILLER_57_697 ();
 sg13g2_decap_4 FILLER_57_704 ();
 sg13g2_fill_1 FILLER_57_708 ();
 sg13g2_decap_4 FILLER_57_730 ();
 sg13g2_fill_1 FILLER_57_734 ();
 sg13g2_fill_2 FILLER_57_749 ();
 sg13g2_fill_1 FILLER_57_751 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_793 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_decap_8 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_decap_8 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_842 ();
 sg13g2_decap_8 FILLER_57_849 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_15 ();
 sg13g2_fill_2 FILLER_58_19 ();
 sg13g2_fill_1 FILLER_58_33 ();
 sg13g2_fill_2 FILLER_58_55 ();
 sg13g2_fill_1 FILLER_58_57 ();
 sg13g2_decap_4 FILLER_58_71 ();
 sg13g2_decap_8 FILLER_58_100 ();
 sg13g2_fill_2 FILLER_58_128 ();
 sg13g2_fill_2 FILLER_58_134 ();
 sg13g2_fill_1 FILLER_58_136 ();
 sg13g2_decap_8 FILLER_58_150 ();
 sg13g2_decap_4 FILLER_58_157 ();
 sg13g2_fill_2 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_4 FILLER_58_186 ();
 sg13g2_fill_1 FILLER_58_190 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_fill_1 FILLER_58_234 ();
 sg13g2_fill_2 FILLER_58_240 ();
 sg13g2_decap_4 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_341 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_decap_8 FILLER_58_369 ();
 sg13g2_fill_1 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_417 ();
 sg13g2_fill_1 FILLER_58_419 ();
 sg13g2_decap_4 FILLER_58_438 ();
 sg13g2_fill_2 FILLER_58_442 ();
 sg13g2_fill_2 FILLER_58_449 ();
 sg13g2_fill_1 FILLER_58_451 ();
 sg13g2_fill_2 FILLER_58_461 ();
 sg13g2_fill_1 FILLER_58_463 ();
 sg13g2_decap_8 FILLER_58_477 ();
 sg13g2_decap_4 FILLER_58_484 ();
 sg13g2_fill_1 FILLER_58_488 ();
 sg13g2_decap_8 FILLER_58_503 ();
 sg13g2_decap_4 FILLER_58_510 ();
 sg13g2_fill_1 FILLER_58_514 ();
 sg13g2_decap_8 FILLER_58_523 ();
 sg13g2_fill_2 FILLER_58_530 ();
 sg13g2_decap_8 FILLER_58_546 ();
 sg13g2_decap_4 FILLER_58_562 ();
 sg13g2_fill_1 FILLER_58_581 ();
 sg13g2_decap_8 FILLER_58_613 ();
 sg13g2_decap_8 FILLER_58_620 ();
 sg13g2_fill_1 FILLER_58_635 ();
 sg13g2_decap_8 FILLER_58_666 ();
 sg13g2_fill_2 FILLER_58_673 ();
 sg13g2_decap_4 FILLER_58_708 ();
 sg13g2_fill_2 FILLER_58_712 ();
 sg13g2_decap_8 FILLER_58_723 ();
 sg13g2_decap_8 FILLER_58_730 ();
 sg13g2_decap_8 FILLER_58_737 ();
 sg13g2_fill_2 FILLER_58_744 ();
 sg13g2_decap_4 FILLER_58_756 ();
 sg13g2_decap_8 FILLER_58_786 ();
 sg13g2_decap_8 FILLER_58_793 ();
 sg13g2_decap_8 FILLER_58_800 ();
 sg13g2_decap_8 FILLER_58_807 ();
 sg13g2_decap_8 FILLER_58_814 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_fill_2 FILLER_59_34 ();
 sg13g2_decap_8 FILLER_59_76 ();
 sg13g2_decap_4 FILLER_59_83 ();
 sg13g2_fill_1 FILLER_59_87 ();
 sg13g2_fill_2 FILLER_59_92 ();
 sg13g2_fill_1 FILLER_59_94 ();
 sg13g2_decap_8 FILLER_59_100 ();
 sg13g2_decap_4 FILLER_59_107 ();
 sg13g2_fill_1 FILLER_59_111 ();
 sg13g2_fill_2 FILLER_59_124 ();
 sg13g2_fill_1 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_145 ();
 sg13g2_fill_2 FILLER_59_152 ();
 sg13g2_fill_2 FILLER_59_166 ();
 sg13g2_fill_1 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_207 ();
 sg13g2_fill_1 FILLER_59_214 ();
 sg13g2_decap_8 FILLER_59_227 ();
 sg13g2_decap_4 FILLER_59_234 ();
 sg13g2_fill_2 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_256 ();
 sg13g2_fill_2 FILLER_59_263 ();
 sg13g2_decap_4 FILLER_59_269 ();
 sg13g2_fill_2 FILLER_59_273 ();
 sg13g2_fill_2 FILLER_59_289 ();
 sg13g2_fill_1 FILLER_59_291 ();
 sg13g2_decap_8 FILLER_59_311 ();
 sg13g2_decap_4 FILLER_59_318 ();
 sg13g2_decap_8 FILLER_59_331 ();
 sg13g2_decap_4 FILLER_59_338 ();
 sg13g2_fill_1 FILLER_59_342 ();
 sg13g2_decap_8 FILLER_59_368 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_decap_4 FILLER_59_382 ();
 sg13g2_fill_1 FILLER_59_386 ();
 sg13g2_fill_1 FILLER_59_401 ();
 sg13g2_fill_2 FILLER_59_454 ();
 sg13g2_fill_2 FILLER_59_483 ();
 sg13g2_fill_1 FILLER_59_507 ();
 sg13g2_fill_2 FILLER_59_521 ();
 sg13g2_decap_4 FILLER_59_532 ();
 sg13g2_fill_2 FILLER_59_536 ();
 sg13g2_fill_1 FILLER_59_568 ();
 sg13g2_decap_8 FILLER_59_573 ();
 sg13g2_fill_2 FILLER_59_611 ();
 sg13g2_fill_1 FILLER_59_613 ();
 sg13g2_fill_1 FILLER_59_618 ();
 sg13g2_decap_4 FILLER_59_627 ();
 sg13g2_fill_1 FILLER_59_649 ();
 sg13g2_decap_8 FILLER_59_678 ();
 sg13g2_fill_1 FILLER_59_685 ();
 sg13g2_decap_8 FILLER_59_702 ();
 sg13g2_decap_4 FILLER_59_709 ();
 sg13g2_fill_2 FILLER_59_739 ();
 sg13g2_decap_8 FILLER_59_767 ();
 sg13g2_decap_8 FILLER_59_774 ();
 sg13g2_decap_8 FILLER_59_781 ();
 sg13g2_decap_8 FILLER_59_788 ();
 sg13g2_decap_8 FILLER_59_795 ();
 sg13g2_decap_8 FILLER_59_802 ();
 sg13g2_decap_8 FILLER_59_809 ();
 sg13g2_decap_8 FILLER_59_816 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_decap_8 FILLER_59_830 ();
 sg13g2_decap_8 FILLER_59_837 ();
 sg13g2_decap_8 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_851 ();
 sg13g2_decap_4 FILLER_59_858 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_fill_2 FILLER_60_14 ();
 sg13g2_fill_1 FILLER_60_25 ();
 sg13g2_fill_1 FILLER_60_46 ();
 sg13g2_fill_1 FILLER_60_51 ();
 sg13g2_fill_1 FILLER_60_61 ();
 sg13g2_decap_4 FILLER_60_76 ();
 sg13g2_fill_2 FILLER_60_80 ();
 sg13g2_fill_2 FILLER_60_90 ();
 sg13g2_decap_8 FILLER_60_100 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_decap_4 FILLER_60_120 ();
 sg13g2_fill_1 FILLER_60_128 ();
 sg13g2_fill_1 FILLER_60_144 ();
 sg13g2_decap_8 FILLER_60_151 ();
 sg13g2_fill_2 FILLER_60_158 ();
 sg13g2_fill_1 FILLER_60_160 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_4 FILLER_60_196 ();
 sg13g2_fill_1 FILLER_60_200 ();
 sg13g2_decap_8 FILLER_60_206 ();
 sg13g2_decap_4 FILLER_60_213 ();
 sg13g2_fill_1 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_227 ();
 sg13g2_fill_1 FILLER_60_229 ();
 sg13g2_fill_1 FILLER_60_240 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_fill_1 FILLER_60_256 ();
 sg13g2_decap_8 FILLER_60_276 ();
 sg13g2_decap_4 FILLER_60_308 ();
 sg13g2_fill_2 FILLER_60_312 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_decap_8 FILLER_60_341 ();
 sg13g2_decap_4 FILLER_60_348 ();
 sg13g2_decap_8 FILLER_60_362 ();
 sg13g2_decap_8 FILLER_60_369 ();
 sg13g2_fill_2 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_384 ();
 sg13g2_fill_2 FILLER_60_391 ();
 sg13g2_fill_1 FILLER_60_393 ();
 sg13g2_fill_2 FILLER_60_425 ();
 sg13g2_fill_1 FILLER_60_427 ();
 sg13g2_decap_8 FILLER_60_454 ();
 sg13g2_decap_4 FILLER_60_461 ();
 sg13g2_fill_2 FILLER_60_474 ();
 sg13g2_decap_8 FILLER_60_479 ();
 sg13g2_decap_4 FILLER_60_486 ();
 sg13g2_fill_1 FILLER_60_490 ();
 sg13g2_fill_1 FILLER_60_495 ();
 sg13g2_decap_8 FILLER_60_506 ();
 sg13g2_decap_4 FILLER_60_513 ();
 sg13g2_fill_2 FILLER_60_537 ();
 sg13g2_fill_1 FILLER_60_539 ();
 sg13g2_fill_2 FILLER_60_561 ();
 sg13g2_fill_2 FILLER_60_573 ();
 sg13g2_fill_1 FILLER_60_575 ();
 sg13g2_fill_1 FILLER_60_602 ();
 sg13g2_fill_2 FILLER_60_629 ();
 sg13g2_fill_2 FILLER_60_663 ();
 sg13g2_decap_4 FILLER_60_677 ();
 sg13g2_fill_2 FILLER_60_681 ();
 sg13g2_fill_2 FILLER_60_694 ();
 sg13g2_fill_1 FILLER_60_696 ();
 sg13g2_fill_2 FILLER_60_701 ();
 sg13g2_decap_8 FILLER_60_720 ();
 sg13g2_fill_2 FILLER_60_727 ();
 sg13g2_fill_1 FILLER_60_729 ();
 sg13g2_fill_2 FILLER_60_737 ();
 sg13g2_fill_1 FILLER_60_739 ();
 sg13g2_decap_8 FILLER_60_758 ();
 sg13g2_decap_4 FILLER_60_765 ();
 sg13g2_decap_8 FILLER_60_782 ();
 sg13g2_decap_8 FILLER_60_789 ();
 sg13g2_decap_8 FILLER_60_796 ();
 sg13g2_decap_8 FILLER_60_803 ();
 sg13g2_decap_8 FILLER_60_810 ();
 sg13g2_decap_8 FILLER_60_817 ();
 sg13g2_decap_8 FILLER_60_824 ();
 sg13g2_decap_8 FILLER_60_831 ();
 sg13g2_decap_8 FILLER_60_838 ();
 sg13g2_decap_8 FILLER_60_845 ();
 sg13g2_decap_8 FILLER_60_852 ();
 sg13g2_fill_2 FILLER_60_859 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_4 FILLER_61_39 ();
 sg13g2_fill_2 FILLER_61_43 ();
 sg13g2_decap_4 FILLER_61_57 ();
 sg13g2_decap_4 FILLER_61_69 ();
 sg13g2_fill_1 FILLER_61_73 ();
 sg13g2_decap_4 FILLER_61_87 ();
 sg13g2_fill_1 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_96 ();
 sg13g2_decap_4 FILLER_61_103 ();
 sg13g2_fill_2 FILLER_61_107 ();
 sg13g2_fill_2 FILLER_61_124 ();
 sg13g2_fill_2 FILLER_61_139 ();
 sg13g2_fill_1 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_152 ();
 sg13g2_fill_2 FILLER_61_162 ();
 sg13g2_decap_4 FILLER_61_189 ();
 sg13g2_fill_1 FILLER_61_193 ();
 sg13g2_decap_4 FILLER_61_206 ();
 sg13g2_fill_2 FILLER_61_210 ();
 sg13g2_decap_4 FILLER_61_239 ();
 sg13g2_fill_2 FILLER_61_243 ();
 sg13g2_decap_8 FILLER_61_253 ();
 sg13g2_fill_2 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_262 ();
 sg13g2_decap_8 FILLER_61_279 ();
 sg13g2_decap_8 FILLER_61_286 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_4 FILLER_61_308 ();
 sg13g2_fill_2 FILLER_61_312 ();
 sg13g2_decap_8 FILLER_61_335 ();
 sg13g2_fill_2 FILLER_61_342 ();
 sg13g2_fill_2 FILLER_61_397 ();
 sg13g2_fill_1 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_408 ();
 sg13g2_fill_2 FILLER_61_415 ();
 sg13g2_fill_1 FILLER_61_417 ();
 sg13g2_fill_2 FILLER_61_423 ();
 sg13g2_fill_1 FILLER_61_425 ();
 sg13g2_decap_8 FILLER_61_444 ();
 sg13g2_decap_8 FILLER_61_451 ();
 sg13g2_decap_8 FILLER_61_458 ();
 sg13g2_decap_4 FILLER_61_465 ();
 sg13g2_fill_1 FILLER_61_469 ();
 sg13g2_decap_4 FILLER_61_475 ();
 sg13g2_fill_2 FILLER_61_479 ();
 sg13g2_decap_8 FILLER_61_507 ();
 sg13g2_decap_4 FILLER_61_514 ();
 sg13g2_fill_2 FILLER_61_518 ();
 sg13g2_decap_8 FILLER_61_533 ();
 sg13g2_decap_4 FILLER_61_540 ();
 sg13g2_fill_2 FILLER_61_544 ();
 sg13g2_fill_1 FILLER_61_585 ();
 sg13g2_fill_2 FILLER_61_599 ();
 sg13g2_decap_8 FILLER_61_609 ();
 sg13g2_fill_2 FILLER_61_616 ();
 sg13g2_fill_2 FILLER_61_626 ();
 sg13g2_fill_1 FILLER_61_628 ();
 sg13g2_fill_1 FILLER_61_647 ();
 sg13g2_fill_1 FILLER_61_664 ();
 sg13g2_decap_8 FILLER_61_669 ();
 sg13g2_decap_4 FILLER_61_676 ();
 sg13g2_fill_1 FILLER_61_701 ();
 sg13g2_decap_4 FILLER_61_715 ();
 sg13g2_fill_1 FILLER_61_736 ();
 sg13g2_fill_1 FILLER_61_747 ();
 sg13g2_fill_1 FILLER_61_761 ();
 sg13g2_decap_8 FILLER_61_788 ();
 sg13g2_decap_8 FILLER_61_795 ();
 sg13g2_decap_8 FILLER_61_802 ();
 sg13g2_decap_8 FILLER_61_809 ();
 sg13g2_decap_8 FILLER_61_816 ();
 sg13g2_decap_8 FILLER_61_823 ();
 sg13g2_decap_8 FILLER_61_830 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_4 FILLER_61_858 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_9 ();
 sg13g2_fill_2 FILLER_62_23 ();
 sg13g2_decap_4 FILLER_62_33 ();
 sg13g2_fill_1 FILLER_62_37 ();
 sg13g2_decap_4 FILLER_62_55 ();
 sg13g2_fill_2 FILLER_62_59 ();
 sg13g2_decap_8 FILLER_62_82 ();
 sg13g2_fill_2 FILLER_62_89 ();
 sg13g2_fill_1 FILLER_62_91 ();
 sg13g2_decap_4 FILLER_62_111 ();
 sg13g2_fill_2 FILLER_62_115 ();
 sg13g2_fill_2 FILLER_62_122 ();
 sg13g2_decap_8 FILLER_62_148 ();
 sg13g2_decap_8 FILLER_62_155 ();
 sg13g2_fill_2 FILLER_62_178 ();
 sg13g2_fill_1 FILLER_62_180 ();
 sg13g2_decap_4 FILLER_62_186 ();
 sg13g2_fill_1 FILLER_62_190 ();
 sg13g2_fill_2 FILLER_62_213 ();
 sg13g2_decap_4 FILLER_62_224 ();
 sg13g2_fill_2 FILLER_62_238 ();
 sg13g2_decap_4 FILLER_62_253 ();
 sg13g2_decap_8 FILLER_62_274 ();
 sg13g2_decap_8 FILLER_62_281 ();
 sg13g2_fill_2 FILLER_62_288 ();
 sg13g2_decap_8 FILLER_62_302 ();
 sg13g2_fill_2 FILLER_62_309 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_decap_4 FILLER_62_345 ();
 sg13g2_fill_1 FILLER_62_349 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_4 FILLER_62_380 ();
 sg13g2_fill_1 FILLER_62_384 ();
 sg13g2_fill_2 FILLER_62_393 ();
 sg13g2_fill_1 FILLER_62_395 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_4 FILLER_62_417 ();
 sg13g2_fill_1 FILLER_62_440 ();
 sg13g2_fill_2 FILLER_62_453 ();
 sg13g2_fill_1 FILLER_62_455 ();
 sg13g2_decap_8 FILLER_62_481 ();
 sg13g2_decap_8 FILLER_62_488 ();
 sg13g2_fill_2 FILLER_62_495 ();
 sg13g2_decap_8 FILLER_62_517 ();
 sg13g2_decap_8 FILLER_62_524 ();
 sg13g2_fill_2 FILLER_62_531 ();
 sg13g2_fill_1 FILLER_62_533 ();
 sg13g2_fill_2 FILLER_62_546 ();
 sg13g2_fill_1 FILLER_62_560 ();
 sg13g2_fill_2 FILLER_62_569 ();
 sg13g2_fill_1 FILLER_62_571 ();
 sg13g2_decap_4 FILLER_62_577 ();
 sg13g2_fill_1 FILLER_62_581 ();
 sg13g2_decap_8 FILLER_62_586 ();
 sg13g2_decap_8 FILLER_62_593 ();
 sg13g2_fill_1 FILLER_62_600 ();
 sg13g2_fill_2 FILLER_62_627 ();
 sg13g2_fill_1 FILLER_62_629 ();
 sg13g2_decap_8 FILLER_62_665 ();
 sg13g2_fill_2 FILLER_62_672 ();
 sg13g2_fill_1 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_711 ();
 sg13g2_fill_2 FILLER_62_721 ();
 sg13g2_fill_1 FILLER_62_723 ();
 sg13g2_fill_1 FILLER_62_733 ();
 sg13g2_fill_2 FILLER_62_738 ();
 sg13g2_fill_2 FILLER_62_758 ();
 sg13g2_decap_8 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_798 ();
 sg13g2_decap_8 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_fill_1 FILLER_63_26 ();
 sg13g2_fill_2 FILLER_63_40 ();
 sg13g2_decap_8 FILLER_63_46 ();
 sg13g2_fill_2 FILLER_63_53 ();
 sg13g2_decap_8 FILLER_63_72 ();
 sg13g2_fill_1 FILLER_63_79 ();
 sg13g2_decap_4 FILLER_63_85 ();
 sg13g2_decap_8 FILLER_63_97 ();
 sg13g2_decap_4 FILLER_63_124 ();
 sg13g2_fill_2 FILLER_63_128 ();
 sg13g2_fill_1 FILLER_63_159 ();
 sg13g2_decap_4 FILLER_63_168 ();
 sg13g2_fill_1 FILLER_63_172 ();
 sg13g2_fill_1 FILLER_63_178 ();
 sg13g2_decap_4 FILLER_63_184 ();
 sg13g2_fill_2 FILLER_63_188 ();
 sg13g2_decap_8 FILLER_63_195 ();
 sg13g2_decap_8 FILLER_63_202 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_fill_2 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_220 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_fill_1 FILLER_63_233 ();
 sg13g2_decap_8 FILLER_63_242 ();
 sg13g2_fill_2 FILLER_63_249 ();
 sg13g2_fill_1 FILLER_63_258 ();
 sg13g2_fill_2 FILLER_63_264 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_fill_2 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_285 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_fill_2 FILLER_63_322 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_decap_4 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_fill_1 FILLER_63_344 ();
 sg13g2_decap_4 FILLER_63_371 ();
 sg13g2_fill_2 FILLER_63_375 ();
 sg13g2_fill_2 FILLER_63_398 ();
 sg13g2_fill_1 FILLER_63_400 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_4 FILLER_63_420 ();
 sg13g2_fill_2 FILLER_63_438 ();
 sg13g2_fill_1 FILLER_63_440 ();
 sg13g2_decap_4 FILLER_63_453 ();
 sg13g2_decap_8 FILLER_63_476 ();
 sg13g2_fill_2 FILLER_63_483 ();
 sg13g2_fill_1 FILLER_63_485 ();
 sg13g2_decap_8 FILLER_63_498 ();
 sg13g2_fill_1 FILLER_63_505 ();
 sg13g2_fill_2 FILLER_63_514 ();
 sg13g2_fill_1 FILLER_63_516 ();
 sg13g2_decap_8 FILLER_63_530 ();
 sg13g2_fill_1 FILLER_63_537 ();
 sg13g2_decap_4 FILLER_63_553 ();
 sg13g2_fill_1 FILLER_63_565 ();
 sg13g2_decap_8 FILLER_63_639 ();
 sg13g2_decap_4 FILLER_63_646 ();
 sg13g2_decap_8 FILLER_63_654 ();
 sg13g2_fill_2 FILLER_63_661 ();
 sg13g2_fill_2 FILLER_63_715 ();
 sg13g2_fill_2 FILLER_63_735 ();
 sg13g2_fill_1 FILLER_63_737 ();
 sg13g2_fill_1 FILLER_63_747 ();
 sg13g2_decap_8 FILLER_63_774 ();
 sg13g2_decap_8 FILLER_63_781 ();
 sg13g2_decap_8 FILLER_63_788 ();
 sg13g2_decap_8 FILLER_63_795 ();
 sg13g2_decap_8 FILLER_63_802 ();
 sg13g2_decap_8 FILLER_63_809 ();
 sg13g2_decap_8 FILLER_63_816 ();
 sg13g2_decap_8 FILLER_63_823 ();
 sg13g2_decap_8 FILLER_63_830 ();
 sg13g2_decap_8 FILLER_63_837 ();
 sg13g2_decap_8 FILLER_63_844 ();
 sg13g2_decap_8 FILLER_63_851 ();
 sg13g2_decap_4 FILLER_63_858 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_15 ();
 sg13g2_fill_2 FILLER_64_34 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_4 FILLER_64_63 ();
 sg13g2_fill_1 FILLER_64_67 ();
 sg13g2_decap_4 FILLER_64_72 ();
 sg13g2_fill_2 FILLER_64_79 ();
 sg13g2_fill_1 FILLER_64_81 ();
 sg13g2_decap_8 FILLER_64_87 ();
 sg13g2_fill_2 FILLER_64_102 ();
 sg13g2_decap_8 FILLER_64_131 ();
 sg13g2_fill_2 FILLER_64_138 ();
 sg13g2_decap_4 FILLER_64_153 ();
 sg13g2_decap_4 FILLER_64_166 ();
 sg13g2_fill_2 FILLER_64_180 ();
 sg13g2_fill_1 FILLER_64_182 ();
 sg13g2_fill_1 FILLER_64_206 ();
 sg13g2_decap_8 FILLER_64_223 ();
 sg13g2_decap_4 FILLER_64_230 ();
 sg13g2_fill_2 FILLER_64_234 ();
 sg13g2_decap_8 FILLER_64_251 ();
 sg13g2_decap_4 FILLER_64_258 ();
 sg13g2_fill_2 FILLER_64_267 ();
 sg13g2_fill_1 FILLER_64_269 ();
 sg13g2_decap_8 FILLER_64_281 ();
 sg13g2_decap_4 FILLER_64_288 ();
 sg13g2_fill_1 FILLER_64_292 ();
 sg13g2_fill_1 FILLER_64_297 ();
 sg13g2_decap_4 FILLER_64_306 ();
 sg13g2_fill_2 FILLER_64_314 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_decap_8 FILLER_64_345 ();
 sg13g2_fill_2 FILLER_64_352 ();
 sg13g2_decap_4 FILLER_64_379 ();
 sg13g2_decap_4 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_403 ();
 sg13g2_decap_8 FILLER_64_418 ();
 sg13g2_decap_8 FILLER_64_425 ();
 sg13g2_fill_1 FILLER_64_432 ();
 sg13g2_decap_4 FILLER_64_441 ();
 sg13g2_decap_4 FILLER_64_456 ();
 sg13g2_decap_4 FILLER_64_471 ();
 sg13g2_fill_2 FILLER_64_475 ();
 sg13g2_decap_8 FILLER_64_503 ();
 sg13g2_fill_1 FILLER_64_522 ();
 sg13g2_decap_8 FILLER_64_549 ();
 sg13g2_decap_8 FILLER_64_556 ();
 sg13g2_fill_2 FILLER_64_563 ();
 sg13g2_decap_8 FILLER_64_570 ();
 sg13g2_decap_8 FILLER_64_577 ();
 sg13g2_fill_2 FILLER_64_611 ();
 sg13g2_fill_1 FILLER_64_613 ();
 sg13g2_fill_2 FILLER_64_640 ();
 sg13g2_fill_1 FILLER_64_642 ();
 sg13g2_decap_8 FILLER_64_646 ();
 sg13g2_fill_2 FILLER_64_653 ();
 sg13g2_fill_1 FILLER_64_655 ();
 sg13g2_decap_8 FILLER_64_660 ();
 sg13g2_decap_8 FILLER_64_667 ();
 sg13g2_decap_4 FILLER_64_674 ();
 sg13g2_fill_2 FILLER_64_678 ();
 sg13g2_fill_2 FILLER_64_685 ();
 sg13g2_fill_2 FILLER_64_696 ();
 sg13g2_decap_8 FILLER_64_715 ();
 sg13g2_fill_1 FILLER_64_722 ();
 sg13g2_decap_4 FILLER_64_753 ();
 sg13g2_fill_2 FILLER_64_757 ();
 sg13g2_decap_8 FILLER_64_768 ();
 sg13g2_decap_8 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_782 ();
 sg13g2_decap_8 FILLER_64_789 ();
 sg13g2_decap_8 FILLER_64_796 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_decap_8 FILLER_64_810 ();
 sg13g2_decap_8 FILLER_64_817 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_15 ();
 sg13g2_fill_2 FILLER_65_25 ();
 sg13g2_fill_1 FILLER_65_27 ();
 sg13g2_fill_1 FILLER_65_38 ();
 sg13g2_decap_4 FILLER_65_101 ();
 sg13g2_decap_4 FILLER_65_110 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_decap_8 FILLER_65_125 ();
 sg13g2_decap_8 FILLER_65_132 ();
 sg13g2_fill_2 FILLER_65_139 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_2 FILLER_65_157 ();
 sg13g2_fill_1 FILLER_65_159 ();
 sg13g2_decap_4 FILLER_65_165 ();
 sg13g2_fill_1 FILLER_65_174 ();
 sg13g2_decap_8 FILLER_65_183 ();
 sg13g2_decap_8 FILLER_65_190 ();
 sg13g2_decap_4 FILLER_65_197 ();
 sg13g2_fill_2 FILLER_65_201 ();
 sg13g2_decap_4 FILLER_65_208 ();
 sg13g2_decap_8 FILLER_65_219 ();
 sg13g2_decap_4 FILLER_65_226 ();
 sg13g2_fill_1 FILLER_65_230 ();
 sg13g2_decap_8 FILLER_65_240 ();
 sg13g2_decap_8 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_284 ();
 sg13g2_fill_2 FILLER_65_291 ();
 sg13g2_fill_1 FILLER_65_293 ();
 sg13g2_decap_4 FILLER_65_302 ();
 sg13g2_fill_1 FILLER_65_314 ();
 sg13g2_decap_8 FILLER_65_324 ();
 sg13g2_fill_2 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_337 ();
 sg13g2_decap_8 FILLER_65_352 ();
 sg13g2_decap_4 FILLER_65_359 ();
 sg13g2_fill_1 FILLER_65_363 ();
 sg13g2_decap_4 FILLER_65_372 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_4 FILLER_65_399 ();
 sg13g2_fill_1 FILLER_65_403 ();
 sg13g2_fill_1 FILLER_65_427 ();
 sg13g2_fill_2 FILLER_65_433 ();
 sg13g2_fill_1 FILLER_65_435 ();
 sg13g2_decap_4 FILLER_65_450 ();
 sg13g2_decap_8 FILLER_65_475 ();
 sg13g2_fill_2 FILLER_65_482 ();
 sg13g2_fill_1 FILLER_65_484 ();
 sg13g2_decap_4 FILLER_65_489 ();
 sg13g2_decap_8 FILLER_65_501 ();
 sg13g2_decap_8 FILLER_65_508 ();
 sg13g2_decap_8 FILLER_65_515 ();
 sg13g2_decap_4 FILLER_65_527 ();
 sg13g2_decap_8 FILLER_65_536 ();
 sg13g2_decap_8 FILLER_65_543 ();
 sg13g2_fill_1 FILLER_65_555 ();
 sg13g2_fill_1 FILLER_65_595 ();
 sg13g2_fill_2 FILLER_65_625 ();
 sg13g2_fill_1 FILLER_65_627 ();
 sg13g2_fill_2 FILLER_65_643 ();
 sg13g2_decap_4 FILLER_65_671 ();
 sg13g2_fill_2 FILLER_65_680 ();
 sg13g2_fill_1 FILLER_65_698 ();
 sg13g2_decap_8 FILLER_65_739 ();
 sg13g2_decap_8 FILLER_65_746 ();
 sg13g2_decap_8 FILLER_65_753 ();
 sg13g2_decap_8 FILLER_65_760 ();
 sg13g2_decap_8 FILLER_65_767 ();
 sg13g2_decap_8 FILLER_65_774 ();
 sg13g2_decap_8 FILLER_65_781 ();
 sg13g2_decap_8 FILLER_65_788 ();
 sg13g2_decap_8 FILLER_65_795 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_decap_8 FILLER_65_809 ();
 sg13g2_decap_8 FILLER_65_816 ();
 sg13g2_decap_8 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_830 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_fill_1 FILLER_66_40 ();
 sg13g2_decap_8 FILLER_66_57 ();
 sg13g2_decap_8 FILLER_66_64 ();
 sg13g2_decap_8 FILLER_66_71 ();
 sg13g2_fill_1 FILLER_66_78 ();
 sg13g2_decap_8 FILLER_66_102 ();
 sg13g2_decap_8 FILLER_66_109 ();
 sg13g2_fill_2 FILLER_66_141 ();
 sg13g2_fill_1 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_152 ();
 sg13g2_fill_1 FILLER_66_159 ();
 sg13g2_decap_4 FILLER_66_177 ();
 sg13g2_fill_1 FILLER_66_181 ();
 sg13g2_fill_1 FILLER_66_193 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_decap_8 FILLER_66_221 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_fill_1 FILLER_66_230 ();
 sg13g2_decap_4 FILLER_66_276 ();
 sg13g2_fill_2 FILLER_66_280 ();
 sg13g2_fill_1 FILLER_66_295 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_fill_2 FILLER_66_332 ();
 sg13g2_fill_1 FILLER_66_334 ();
 sg13g2_decap_8 FILLER_66_351 ();
 sg13g2_decap_4 FILLER_66_358 ();
 sg13g2_decap_8 FILLER_66_367 ();
 sg13g2_decap_4 FILLER_66_374 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_fill_1 FILLER_66_387 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_66_421 ();
 sg13g2_fill_1 FILLER_66_423 ();
 sg13g2_fill_2 FILLER_66_435 ();
 sg13g2_fill_1 FILLER_66_437 ();
 sg13g2_decap_8 FILLER_66_443 ();
 sg13g2_decap_8 FILLER_66_450 ();
 sg13g2_decap_4 FILLER_66_457 ();
 sg13g2_fill_2 FILLER_66_465 ();
 sg13g2_decap_8 FILLER_66_484 ();
 sg13g2_fill_1 FILLER_66_491 ();
 sg13g2_decap_4 FILLER_66_508 ();
 sg13g2_fill_1 FILLER_66_512 ();
 sg13g2_decap_4 FILLER_66_540 ();
 sg13g2_decap_8 FILLER_66_558 ();
 sg13g2_fill_2 FILLER_66_565 ();
 sg13g2_fill_2 FILLER_66_580 ();
 sg13g2_decap_4 FILLER_66_592 ();
 sg13g2_fill_1 FILLER_66_596 ();
 sg13g2_fill_2 FILLER_66_617 ();
 sg13g2_fill_1 FILLER_66_627 ();
 sg13g2_decap_8 FILLER_66_634 ();
 sg13g2_fill_1 FILLER_66_641 ();
 sg13g2_decap_4 FILLER_66_651 ();
 sg13g2_decap_8 FILLER_66_681 ();
 sg13g2_decap_4 FILLER_66_688 ();
 sg13g2_decap_4 FILLER_66_705 ();
 sg13g2_fill_1 FILLER_66_709 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_decap_4 FILLER_66_721 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_37 ();
 sg13g2_fill_2 FILLER_67_69 ();
 sg13g2_decap_4 FILLER_67_74 ();
 sg13g2_fill_1 FILLER_67_78 ();
 sg13g2_fill_1 FILLER_67_100 ();
 sg13g2_fill_2 FILLER_67_110 ();
 sg13g2_decap_8 FILLER_67_124 ();
 sg13g2_fill_2 FILLER_67_131 ();
 sg13g2_fill_1 FILLER_67_133 ();
 sg13g2_decap_4 FILLER_67_138 ();
 sg13g2_fill_2 FILLER_67_146 ();
 sg13g2_decap_4 FILLER_67_156 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_fill_1 FILLER_67_182 ();
 sg13g2_decap_4 FILLER_67_187 ();
 sg13g2_decap_8 FILLER_67_199 ();
 sg13g2_fill_2 FILLER_67_206 ();
 sg13g2_decap_4 FILLER_67_221 ();
 sg13g2_fill_1 FILLER_67_225 ();
 sg13g2_fill_1 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_244 ();
 sg13g2_fill_2 FILLER_67_251 ();
 sg13g2_decap_4 FILLER_67_277 ();
 sg13g2_fill_1 FILLER_67_281 ();
 sg13g2_fill_2 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_299 ();
 sg13g2_fill_2 FILLER_67_310 ();
 sg13g2_fill_1 FILLER_67_312 ();
 sg13g2_fill_1 FILLER_67_326 ();
 sg13g2_decap_8 FILLER_67_337 ();
 sg13g2_decap_8 FILLER_67_344 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_decap_8 FILLER_67_379 ();
 sg13g2_decap_4 FILLER_67_386 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_fill_1 FILLER_67_414 ();
 sg13g2_decap_8 FILLER_67_423 ();
 sg13g2_decap_4 FILLER_67_430 ();
 sg13g2_fill_1 FILLER_67_434 ();
 sg13g2_decap_4 FILLER_67_441 ();
 sg13g2_fill_1 FILLER_67_445 ();
 sg13g2_decap_8 FILLER_67_462 ();
 sg13g2_fill_1 FILLER_67_469 ();
 sg13g2_fill_2 FILLER_67_486 ();
 sg13g2_fill_1 FILLER_67_488 ();
 sg13g2_decap_4 FILLER_67_515 ();
 sg13g2_fill_2 FILLER_67_519 ();
 sg13g2_decap_8 FILLER_67_529 ();
 sg13g2_decap_8 FILLER_67_536 ();
 sg13g2_fill_2 FILLER_67_543 ();
 sg13g2_fill_1 FILLER_67_545 ();
 sg13g2_decap_4 FILLER_67_559 ();
 sg13g2_decap_4 FILLER_67_589 ();
 sg13g2_fill_1 FILLER_67_593 ();
 sg13g2_decap_8 FILLER_67_606 ();
 sg13g2_decap_4 FILLER_67_613 ();
 sg13g2_fill_2 FILLER_67_617 ();
 sg13g2_decap_8 FILLER_67_624 ();
 sg13g2_fill_2 FILLER_67_631 ();
 sg13g2_decap_4 FILLER_67_643 ();
 sg13g2_fill_1 FILLER_67_647 ();
 sg13g2_fill_2 FILLER_67_663 ();
 sg13g2_fill_1 FILLER_67_665 ();
 sg13g2_fill_1 FILLER_67_705 ();
 sg13g2_decap_8 FILLER_67_739 ();
 sg13g2_decap_8 FILLER_67_746 ();
 sg13g2_decap_8 FILLER_67_753 ();
 sg13g2_decap_8 FILLER_67_760 ();
 sg13g2_decap_8 FILLER_67_767 ();
 sg13g2_decap_8 FILLER_67_774 ();
 sg13g2_decap_8 FILLER_67_781 ();
 sg13g2_decap_8 FILLER_67_788 ();
 sg13g2_decap_8 FILLER_67_795 ();
 sg13g2_decap_8 FILLER_67_802 ();
 sg13g2_decap_8 FILLER_67_809 ();
 sg13g2_decap_8 FILLER_67_816 ();
 sg13g2_decap_8 FILLER_67_823 ();
 sg13g2_decap_8 FILLER_67_830 ();
 sg13g2_decap_8 FILLER_67_837 ();
 sg13g2_decap_8 FILLER_67_844 ();
 sg13g2_decap_8 FILLER_67_851 ();
 sg13g2_decap_4 FILLER_67_858 ();
 sg13g2_fill_2 FILLER_68_40 ();
 sg13g2_decap_4 FILLER_68_55 ();
 sg13g2_fill_2 FILLER_68_59 ();
 sg13g2_decap_8 FILLER_68_118 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_fill_2 FILLER_68_144 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_163 ();
 sg13g2_decap_8 FILLER_68_191 ();
 sg13g2_decap_8 FILLER_68_198 ();
 sg13g2_decap_4 FILLER_68_205 ();
 sg13g2_fill_2 FILLER_68_209 ();
 sg13g2_decap_8 FILLER_68_221 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_243 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_252 ();
 sg13g2_decap_8 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_276 ();
 sg13g2_decap_8 FILLER_68_283 ();
 sg13g2_decap_4 FILLER_68_290 ();
 sg13g2_fill_2 FILLER_68_294 ();
 sg13g2_fill_2 FILLER_68_309 ();
 sg13g2_decap_8 FILLER_68_326 ();
 sg13g2_fill_1 FILLER_68_333 ();
 sg13g2_decap_4 FILLER_68_339 ();
 sg13g2_fill_2 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_351 ();
 sg13g2_decap_4 FILLER_68_358 ();
 sg13g2_fill_2 FILLER_68_390 ();
 sg13g2_fill_1 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_406 ();
 sg13g2_fill_2 FILLER_68_413 ();
 sg13g2_decap_8 FILLER_68_421 ();
 sg13g2_decap_4 FILLER_68_428 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_decap_4 FILLER_68_459 ();
 sg13g2_fill_1 FILLER_68_463 ();
 sg13g2_decap_8 FILLER_68_473 ();
 sg13g2_decap_8 FILLER_68_480 ();
 sg13g2_decap_8 FILLER_68_487 ();
 sg13g2_decap_8 FILLER_68_507 ();
 sg13g2_decap_8 FILLER_68_514 ();
 sg13g2_decap_8 FILLER_68_521 ();
 sg13g2_decap_8 FILLER_68_528 ();
 sg13g2_decap_4 FILLER_68_535 ();
 sg13g2_fill_2 FILLER_68_543 ();
 sg13g2_fill_1 FILLER_68_545 ();
 sg13g2_fill_1 FILLER_68_551 ();
 sg13g2_decap_8 FILLER_68_565 ();
 sg13g2_fill_1 FILLER_68_572 ();
 sg13g2_fill_2 FILLER_68_582 ();
 sg13g2_fill_2 FILLER_68_626 ();
 sg13g2_decap_4 FILLER_68_633 ();
 sg13g2_decap_8 FILLER_68_641 ();
 sg13g2_decap_8 FILLER_68_648 ();
 sg13g2_decap_4 FILLER_68_655 ();
 sg13g2_fill_1 FILLER_68_659 ();
 sg13g2_decap_8 FILLER_68_675 ();
 sg13g2_decap_4 FILLER_68_682 ();
 sg13g2_fill_2 FILLER_68_691 ();
 sg13g2_fill_1 FILLER_68_693 ();
 sg13g2_decap_8 FILLER_68_702 ();
 sg13g2_decap_8 FILLER_68_709 ();
 sg13g2_decap_8 FILLER_68_716 ();
 sg13g2_decap_8 FILLER_68_736 ();
 sg13g2_decap_8 FILLER_68_743 ();
 sg13g2_decap_8 FILLER_68_750 ();
 sg13g2_decap_8 FILLER_68_757 ();
 sg13g2_decap_8 FILLER_68_764 ();
 sg13g2_decap_8 FILLER_68_771 ();
 sg13g2_decap_8 FILLER_68_778 ();
 sg13g2_decap_8 FILLER_68_785 ();
 sg13g2_decap_8 FILLER_68_792 ();
 sg13g2_decap_8 FILLER_68_799 ();
 sg13g2_decap_8 FILLER_68_806 ();
 sg13g2_decap_8 FILLER_68_813 ();
 sg13g2_decap_8 FILLER_68_820 ();
 sg13g2_decap_8 FILLER_68_827 ();
 sg13g2_decap_8 FILLER_68_834 ();
 sg13g2_decap_8 FILLER_68_841 ();
 sg13g2_decap_8 FILLER_68_848 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_decap_4 FILLER_69_15 ();
 sg13g2_fill_2 FILLER_69_19 ();
 sg13g2_fill_1 FILLER_69_39 ();
 sg13g2_decap_4 FILLER_69_49 ();
 sg13g2_fill_1 FILLER_69_53 ();
 sg13g2_decap_4 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_79 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_decap_8 FILLER_69_99 ();
 sg13g2_decap_8 FILLER_69_106 ();
 sg13g2_decap_4 FILLER_69_113 ();
 sg13g2_fill_2 FILLER_69_117 ();
 sg13g2_decap_8 FILLER_69_129 ();
 sg13g2_decap_4 FILLER_69_136 ();
 sg13g2_decap_8 FILLER_69_156 ();
 sg13g2_decap_4 FILLER_69_163 ();
 sg13g2_decap_8 FILLER_69_186 ();
 sg13g2_decap_4 FILLER_69_193 ();
 sg13g2_decap_8 FILLER_69_222 ();
 sg13g2_fill_1 FILLER_69_229 ();
 sg13g2_decap_8 FILLER_69_239 ();
 sg13g2_fill_2 FILLER_69_257 ();
 sg13g2_fill_1 FILLER_69_259 ();
 sg13g2_fill_2 FILLER_69_269 ();
 sg13g2_fill_2 FILLER_69_302 ();
 sg13g2_decap_8 FILLER_69_312 ();
 sg13g2_fill_2 FILLER_69_329 ();
 sg13g2_fill_1 FILLER_69_331 ();
 sg13g2_decap_8 FILLER_69_360 ();
 sg13g2_decap_4 FILLER_69_367 ();
 sg13g2_fill_1 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_decap_4 FILLER_69_408 ();
 sg13g2_fill_1 FILLER_69_433 ();
 sg13g2_decap_8 FILLER_69_453 ();
 sg13g2_decap_8 FILLER_69_478 ();
 sg13g2_fill_2 FILLER_69_495 ();
 sg13g2_fill_2 FILLER_69_502 ();
 sg13g2_fill_1 FILLER_69_504 ();
 sg13g2_fill_1 FILLER_69_511 ();
 sg13g2_fill_2 FILLER_69_526 ();
 sg13g2_decap_8 FILLER_69_558 ();
 sg13g2_decap_8 FILLER_69_565 ();
 sg13g2_fill_2 FILLER_69_572 ();
 sg13g2_fill_1 FILLER_69_582 ();
 sg13g2_decap_4 FILLER_69_592 ();
 sg13g2_decap_4 FILLER_69_601 ();
 sg13g2_fill_1 FILLER_69_605 ();
 sg13g2_decap_4 FILLER_69_615 ();
 sg13g2_fill_1 FILLER_69_619 ();
 sg13g2_fill_1 FILLER_69_646 ();
 sg13g2_fill_2 FILLER_69_656 ();
 sg13g2_fill_2 FILLER_69_663 ();
 sg13g2_fill_1 FILLER_69_665 ();
 sg13g2_decap_8 FILLER_69_671 ();
 sg13g2_decap_8 FILLER_69_678 ();
 sg13g2_fill_2 FILLER_69_685 ();
 sg13g2_fill_2 FILLER_69_704 ();
 sg13g2_decap_4 FILLER_69_732 ();
 sg13g2_fill_2 FILLER_69_736 ();
 sg13g2_decap_8 FILLER_69_750 ();
 sg13g2_decap_8 FILLER_69_757 ();
 sg13g2_decap_8 FILLER_69_764 ();
 sg13g2_decap_8 FILLER_69_771 ();
 sg13g2_decap_8 FILLER_69_778 ();
 sg13g2_decap_8 FILLER_69_785 ();
 sg13g2_decap_8 FILLER_69_792 ();
 sg13g2_decap_8 FILLER_69_799 ();
 sg13g2_decap_8 FILLER_69_806 ();
 sg13g2_decap_8 FILLER_69_813 ();
 sg13g2_decap_8 FILLER_69_820 ();
 sg13g2_decap_8 FILLER_69_827 ();
 sg13g2_decap_8 FILLER_69_834 ();
 sg13g2_decap_8 FILLER_69_841 ();
 sg13g2_decap_8 FILLER_69_848 ();
 sg13g2_decap_8 FILLER_69_855 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_21 ();
 sg13g2_fill_1 FILLER_70_23 ();
 sg13g2_decap_4 FILLER_70_50 ();
 sg13g2_fill_2 FILLER_70_54 ();
 sg13g2_fill_1 FILLER_70_82 ();
 sg13g2_fill_2 FILLER_70_101 ();
 sg13g2_fill_2 FILLER_70_107 ();
 sg13g2_decap_4 FILLER_70_114 ();
 sg13g2_fill_1 FILLER_70_118 ();
 sg13g2_decap_4 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_132 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_fill_2 FILLER_70_168 ();
 sg13g2_fill_2 FILLER_70_200 ();
 sg13g2_fill_1 FILLER_70_202 ();
 sg13g2_fill_2 FILLER_70_208 ();
 sg13g2_decap_4 FILLER_70_215 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_decap_4 FILLER_70_249 ();
 sg13g2_fill_2 FILLER_70_260 ();
 sg13g2_fill_2 FILLER_70_267 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_1 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_303 ();
 sg13g2_fill_1 FILLER_70_305 ();
 sg13g2_decap_8 FILLER_70_325 ();
 sg13g2_fill_1 FILLER_70_332 ();
 sg13g2_decap_4 FILLER_70_338 ();
 sg13g2_decap_8 FILLER_70_346 ();
 sg13g2_decap_8 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_fill_2 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_4 FILLER_70_392 ();
 sg13g2_fill_1 FILLER_70_396 ();
 sg13g2_decap_4 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_70_420 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_442 ();
 sg13g2_decap_8 FILLER_70_449 ();
 sg13g2_decap_4 FILLER_70_456 ();
 sg13g2_fill_2 FILLER_70_460 ();
 sg13g2_decap_8 FILLER_70_472 ();
 sg13g2_decap_8 FILLER_70_479 ();
 sg13g2_fill_1 FILLER_70_486 ();
 sg13g2_decap_4 FILLER_70_499 ();
 sg13g2_decap_4 FILLER_70_508 ();
 sg13g2_fill_1 FILLER_70_512 ();
 sg13g2_decap_4 FILLER_70_517 ();
 sg13g2_fill_1 FILLER_70_521 ();
 sg13g2_fill_1 FILLER_70_529 ();
 sg13g2_decap_8 FILLER_70_535 ();
 sg13g2_decap_4 FILLER_70_542 ();
 sg13g2_fill_1 FILLER_70_546 ();
 sg13g2_fill_1 FILLER_70_564 ();
 sg13g2_fill_1 FILLER_70_569 ();
 sg13g2_decap_8 FILLER_70_593 ();
 sg13g2_decap_4 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_628 ();
 sg13g2_fill_1 FILLER_70_642 ();
 sg13g2_fill_2 FILLER_70_647 ();
 sg13g2_decap_4 FILLER_70_661 ();
 sg13g2_fill_1 FILLER_70_711 ();
 sg13g2_decap_8 FILLER_70_765 ();
 sg13g2_decap_8 FILLER_70_772 ();
 sg13g2_decap_8 FILLER_70_779 ();
 sg13g2_decap_8 FILLER_70_786 ();
 sg13g2_decap_8 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_800 ();
 sg13g2_decap_8 FILLER_70_807 ();
 sg13g2_decap_8 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_821 ();
 sg13g2_decap_8 FILLER_70_828 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_84 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_95 ();
 sg13g2_fill_1 FILLER_71_136 ();
 sg13g2_decap_8 FILLER_71_155 ();
 sg13g2_fill_2 FILLER_71_162 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_decap_4 FILLER_71_172 ();
 sg13g2_fill_2 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_4 FILLER_71_189 ();
 sg13g2_fill_2 FILLER_71_193 ();
 sg13g2_decap_8 FILLER_71_204 ();
 sg13g2_decap_8 FILLER_71_211 ();
 sg13g2_fill_1 FILLER_71_218 ();
 sg13g2_decap_8 FILLER_71_223 ();
 sg13g2_decap_8 FILLER_71_230 ();
 sg13g2_fill_2 FILLER_71_237 ();
 sg13g2_fill_1 FILLER_71_239 ();
 sg13g2_decap_8 FILLER_71_244 ();
 sg13g2_decap_8 FILLER_71_251 ();
 sg13g2_fill_1 FILLER_71_258 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_fill_1 FILLER_71_294 ();
 sg13g2_decap_4 FILLER_71_305 ();
 sg13g2_decap_8 FILLER_71_314 ();
 sg13g2_decap_4 FILLER_71_321 ();
 sg13g2_fill_1 FILLER_71_325 ();
 sg13g2_decap_4 FILLER_71_330 ();
 sg13g2_fill_2 FILLER_71_334 ();
 sg13g2_fill_1 FILLER_71_344 ();
 sg13g2_decap_8 FILLER_71_349 ();
 sg13g2_fill_2 FILLER_71_356 ();
 sg13g2_fill_1 FILLER_71_358 ();
 sg13g2_decap_4 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_386 ();
 sg13g2_fill_2 FILLER_71_393 ();
 sg13g2_fill_1 FILLER_71_395 ();
 sg13g2_decap_4 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_71_411 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_fill_1 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_452 ();
 sg13g2_fill_2 FILLER_71_458 ();
 sg13g2_fill_2 FILLER_71_478 ();
 sg13g2_decap_4 FILLER_71_487 ();
 sg13g2_fill_2 FILLER_71_510 ();
 sg13g2_fill_1 FILLER_71_512 ();
 sg13g2_decap_8 FILLER_71_529 ();
 sg13g2_decap_4 FILLER_71_539 ();
 sg13g2_fill_1 FILLER_71_543 ();
 sg13g2_decap_8 FILLER_71_580 ();
 sg13g2_decap_8 FILLER_71_592 ();
 sg13g2_decap_8 FILLER_71_599 ();
 sg13g2_fill_1 FILLER_71_606 ();
 sg13g2_decap_8 FILLER_71_611 ();
 sg13g2_decap_8 FILLER_71_618 ();
 sg13g2_fill_1 FILLER_71_625 ();
 sg13g2_fill_1 FILLER_71_631 ();
 sg13g2_fill_2 FILLER_71_647 ();
 sg13g2_fill_1 FILLER_71_649 ();
 sg13g2_fill_2 FILLER_71_664 ();
 sg13g2_fill_1 FILLER_71_666 ();
 sg13g2_decap_4 FILLER_71_683 ();
 sg13g2_decap_8 FILLER_71_699 ();
 sg13g2_fill_2 FILLER_71_706 ();
 sg13g2_fill_1 FILLER_71_712 ();
 sg13g2_fill_1 FILLER_71_717 ();
 sg13g2_fill_2 FILLER_71_746 ();
 sg13g2_fill_2 FILLER_71_761 ();
 sg13g2_decap_8 FILLER_71_767 ();
 sg13g2_decap_8 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_781 ();
 sg13g2_decap_8 FILLER_71_788 ();
 sg13g2_decap_8 FILLER_71_795 ();
 sg13g2_decap_8 FILLER_71_802 ();
 sg13g2_decap_8 FILLER_71_809 ();
 sg13g2_decap_8 FILLER_71_816 ();
 sg13g2_decap_8 FILLER_71_823 ();
 sg13g2_decap_8 FILLER_71_830 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_844 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_4 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_84 ();
 sg13g2_decap_4 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_142 ();
 sg13g2_decap_8 FILLER_72_149 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_183 ();
 sg13g2_fill_1 FILLER_72_230 ();
 sg13g2_fill_2 FILLER_72_236 ();
 sg13g2_decap_8 FILLER_72_250 ();
 sg13g2_fill_2 FILLER_72_276 ();
 sg13g2_fill_1 FILLER_72_278 ();
 sg13g2_fill_2 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_287 ();
 sg13g2_decap_4 FILLER_72_309 ();
 sg13g2_fill_2 FILLER_72_313 ();
 sg13g2_fill_1 FILLER_72_320 ();
 sg13g2_fill_1 FILLER_72_328 ();
 sg13g2_fill_2 FILLER_72_350 ();
 sg13g2_decap_4 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_368 ();
 sg13g2_fill_2 FILLER_72_374 ();
 sg13g2_fill_1 FILLER_72_395 ();
 sg13g2_fill_1 FILLER_72_414 ();
 sg13g2_decap_4 FILLER_72_421 ();
 sg13g2_fill_2 FILLER_72_425 ();
 sg13g2_decap_8 FILLER_72_433 ();
 sg13g2_fill_2 FILLER_72_440 ();
 sg13g2_fill_1 FILLER_72_442 ();
 sg13g2_fill_1 FILLER_72_457 ();
 sg13g2_fill_1 FILLER_72_463 ();
 sg13g2_fill_1 FILLER_72_468 ();
 sg13g2_decap_8 FILLER_72_474 ();
 sg13g2_decap_8 FILLER_72_481 ();
 sg13g2_fill_1 FILLER_72_488 ();
 sg13g2_fill_2 FILLER_72_505 ();
 sg13g2_fill_1 FILLER_72_507 ();
 sg13g2_fill_2 FILLER_72_517 ();
 sg13g2_decap_4 FILLER_72_524 ();
 sg13g2_decap_4 FILLER_72_548 ();
 sg13g2_fill_2 FILLER_72_577 ();
 sg13g2_fill_1 FILLER_72_579 ();
 sg13g2_fill_2 FILLER_72_588 ();
 sg13g2_decap_8 FILLER_72_606 ();
 sg13g2_fill_1 FILLER_72_613 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_fill_2 FILLER_72_672 ();
 sg13g2_fill_1 FILLER_72_674 ();
 sg13g2_fill_1 FILLER_72_680 ();
 sg13g2_decap_4 FILLER_72_685 ();
 sg13g2_decap_4 FILLER_72_698 ();
 sg13g2_fill_1 FILLER_72_702 ();
 sg13g2_decap_4 FILLER_72_747 ();
 sg13g2_fill_1 FILLER_72_751 ();
 sg13g2_decap_8 FILLER_72_778 ();
 sg13g2_decap_8 FILLER_72_785 ();
 sg13g2_decap_8 FILLER_72_792 ();
 sg13g2_decap_8 FILLER_72_799 ();
 sg13g2_decap_8 FILLER_72_806 ();
 sg13g2_decap_8 FILLER_72_813 ();
 sg13g2_decap_8 FILLER_72_820 ();
 sg13g2_decap_8 FILLER_72_827 ();
 sg13g2_decap_8 FILLER_72_834 ();
 sg13g2_decap_8 FILLER_72_841 ();
 sg13g2_decap_8 FILLER_72_848 ();
 sg13g2_decap_8 FILLER_72_855 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_4 FILLER_73_91 ();
 sg13g2_fill_2 FILLER_73_95 ();
 sg13g2_decap_8 FILLER_73_106 ();
 sg13g2_decap_8 FILLER_73_113 ();
 sg13g2_decap_4 FILLER_73_120 ();
 sg13g2_fill_2 FILLER_73_124 ();
 sg13g2_decap_8 FILLER_73_139 ();
 sg13g2_decap_8 FILLER_73_146 ();
 sg13g2_fill_2 FILLER_73_153 ();
 sg13g2_fill_1 FILLER_73_155 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_decap_8 FILLER_73_183 ();
 sg13g2_decap_4 FILLER_73_195 ();
 sg13g2_fill_2 FILLER_73_199 ();
 sg13g2_decap_4 FILLER_73_212 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_fill_2 FILLER_73_238 ();
 sg13g2_fill_2 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_fill_2 FILLER_73_263 ();
 sg13g2_decap_4 FILLER_73_270 ();
 sg13g2_decap_4 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_289 ();
 sg13g2_fill_2 FILLER_73_296 ();
 sg13g2_decap_8 FILLER_73_302 ();
 sg13g2_decap_8 FILLER_73_309 ();
 sg13g2_fill_1 FILLER_73_316 ();
 sg13g2_decap_8 FILLER_73_331 ();
 sg13g2_decap_8 FILLER_73_338 ();
 sg13g2_decap_4 FILLER_73_345 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_4 FILLER_73_366 ();
 sg13g2_decap_4 FILLER_73_375 ();
 sg13g2_decap_4 FILLER_73_385 ();
 sg13g2_fill_2 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_73_421 ();
 sg13g2_decap_8 FILLER_73_444 ();
 sg13g2_decap_8 FILLER_73_451 ();
 sg13g2_decap_4 FILLER_73_458 ();
 sg13g2_fill_2 FILLER_73_462 ();
 sg13g2_decap_4 FILLER_73_477 ();
 sg13g2_decap_8 FILLER_73_499 ();
 sg13g2_fill_1 FILLER_73_506 ();
 sg13g2_decap_4 FILLER_73_520 ();
 sg13g2_decap_8 FILLER_73_543 ();
 sg13g2_decap_8 FILLER_73_550 ();
 sg13g2_decap_8 FILLER_73_557 ();
 sg13g2_decap_8 FILLER_73_564 ();
 sg13g2_decap_8 FILLER_73_571 ();
 sg13g2_decap_4 FILLER_73_578 ();
 sg13g2_fill_2 FILLER_73_582 ();
 sg13g2_decap_4 FILLER_73_646 ();
 sg13g2_fill_2 FILLER_73_650 ();
 sg13g2_decap_8 FILLER_73_657 ();
 sg13g2_decap_4 FILLER_73_664 ();
 sg13g2_fill_2 FILLER_73_668 ();
 sg13g2_decap_8 FILLER_73_696 ();
 sg13g2_decap_8 FILLER_73_703 ();
 sg13g2_decap_8 FILLER_73_710 ();
 sg13g2_fill_1 FILLER_73_717 ();
 sg13g2_decap_8 FILLER_73_768 ();
 sg13g2_decap_8 FILLER_73_775 ();
 sg13g2_decap_8 FILLER_73_782 ();
 sg13g2_decap_8 FILLER_73_789 ();
 sg13g2_decap_8 FILLER_73_796 ();
 sg13g2_decap_8 FILLER_73_803 ();
 sg13g2_decap_8 FILLER_73_810 ();
 sg13g2_decap_8 FILLER_73_817 ();
 sg13g2_decap_8 FILLER_73_824 ();
 sg13g2_decap_8 FILLER_73_831 ();
 sg13g2_decap_8 FILLER_73_838 ();
 sg13g2_decap_8 FILLER_73_845 ();
 sg13g2_decap_8 FILLER_73_852 ();
 sg13g2_fill_2 FILLER_73_859 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_fill_1 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_150 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_decap_8 FILLER_74_232 ();
 sg13g2_fill_2 FILLER_74_239 ();
 sg13g2_fill_1 FILLER_74_241 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_fill_1 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_292 ();
 sg13g2_decap_4 FILLER_74_310 ();
 sg13g2_decap_8 FILLER_74_337 ();
 sg13g2_decap_4 FILLER_74_344 ();
 sg13g2_fill_2 FILLER_74_348 ();
 sg13g2_fill_2 FILLER_74_366 ();
 sg13g2_fill_1 FILLER_74_368 ();
 sg13g2_decap_8 FILLER_74_388 ();
 sg13g2_fill_2 FILLER_74_400 ();
 sg13g2_fill_1 FILLER_74_402 ();
 sg13g2_decap_8 FILLER_74_409 ();
 sg13g2_fill_2 FILLER_74_416 ();
 sg13g2_fill_1 FILLER_74_418 ();
 sg13g2_fill_2 FILLER_74_424 ();
 sg13g2_fill_2 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_437 ();
 sg13g2_decap_8 FILLER_74_448 ();
 sg13g2_fill_2 FILLER_74_455 ();
 sg13g2_decap_8 FILLER_74_466 ();
 sg13g2_fill_2 FILLER_74_484 ();
 sg13g2_fill_2 FILLER_74_506 ();
 sg13g2_decap_4 FILLER_74_513 ();
 sg13g2_decap_8 FILLER_74_544 ();
 sg13g2_decap_8 FILLER_74_551 ();
 sg13g2_fill_2 FILLER_74_571 ();
 sg13g2_fill_1 FILLER_74_573 ();
 sg13g2_fill_2 FILLER_74_591 ();
 sg13g2_decap_8 FILLER_74_607 ();
 sg13g2_fill_2 FILLER_74_614 ();
 sg13g2_fill_1 FILLER_74_616 ();
 sg13g2_fill_2 FILLER_74_622 ();
 sg13g2_fill_1 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_678 ();
 sg13g2_decap_8 FILLER_74_688 ();
 sg13g2_decap_8 FILLER_74_695 ();
 sg13g2_decap_8 FILLER_74_702 ();
 sg13g2_decap_8 FILLER_74_709 ();
 sg13g2_decap_8 FILLER_74_716 ();
 sg13g2_decap_8 FILLER_74_758 ();
 sg13g2_decap_8 FILLER_74_765 ();
 sg13g2_decap_8 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_786 ();
 sg13g2_decap_8 FILLER_74_793 ();
 sg13g2_decap_8 FILLER_74_800 ();
 sg13g2_decap_8 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_814 ();
 sg13g2_decap_8 FILLER_74_821 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_decap_8 FILLER_74_835 ();
 sg13g2_decap_8 FILLER_74_842 ();
 sg13g2_decap_8 FILLER_74_849 ();
 sg13g2_decap_4 FILLER_74_856 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_fill_2 FILLER_75_154 ();
 sg13g2_fill_1 FILLER_75_156 ();
 sg13g2_decap_8 FILLER_75_178 ();
 sg13g2_decap_8 FILLER_75_185 ();
 sg13g2_decap_8 FILLER_75_192 ();
 sg13g2_decap_8 FILLER_75_207 ();
 sg13g2_decap_8 FILLER_75_214 ();
 sg13g2_fill_2 FILLER_75_221 ();
 sg13g2_decap_4 FILLER_75_257 ();
 sg13g2_fill_2 FILLER_75_261 ();
 sg13g2_fill_2 FILLER_75_272 ();
 sg13g2_fill_1 FILLER_75_274 ();
 sg13g2_decap_8 FILLER_75_282 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_fill_2 FILLER_75_316 ();
 sg13g2_fill_1 FILLER_75_318 ();
 sg13g2_decap_4 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_339 ();
 sg13g2_fill_2 FILLER_75_346 ();
 sg13g2_decap_4 FILLER_75_351 ();
 sg13g2_decap_4 FILLER_75_358 ();
 sg13g2_fill_2 FILLER_75_362 ();
 sg13g2_decap_4 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_fill_2 FILLER_75_390 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_decap_4 FILLER_75_413 ();
 sg13g2_fill_2 FILLER_75_417 ();
 sg13g2_decap_8 FILLER_75_439 ();
 sg13g2_decap_8 FILLER_75_446 ();
 sg13g2_decap_8 FILLER_75_473 ();
 sg13g2_decap_4 FILLER_75_480 ();
 sg13g2_fill_2 FILLER_75_484 ();
 sg13g2_fill_1 FILLER_75_495 ();
 sg13g2_decap_8 FILLER_75_505 ();
 sg13g2_decap_8 FILLER_75_512 ();
 sg13g2_fill_2 FILLER_75_519 ();
 sg13g2_fill_1 FILLER_75_521 ();
 sg13g2_fill_2 FILLER_75_526 ();
 sg13g2_decap_4 FILLER_75_551 ();
 sg13g2_fill_1 FILLER_75_555 ();
 sg13g2_decap_4 FILLER_75_627 ();
 sg13g2_fill_2 FILLER_75_631 ();
 sg13g2_decap_8 FILLER_75_643 ();
 sg13g2_decap_8 FILLER_75_650 ();
 sg13g2_decap_4 FILLER_75_657 ();
 sg13g2_fill_2 FILLER_75_661 ();
 sg13g2_decap_8 FILLER_75_667 ();
 sg13g2_decap_4 FILLER_75_674 ();
 sg13g2_decap_8 FILLER_75_681 ();
 sg13g2_decap_8 FILLER_75_688 ();
 sg13g2_decap_8 FILLER_75_695 ();
 sg13g2_decap_8 FILLER_75_702 ();
 sg13g2_decap_8 FILLER_75_709 ();
 sg13g2_decap_8 FILLER_75_716 ();
 sg13g2_decap_8 FILLER_75_723 ();
 sg13g2_decap_4 FILLER_75_730 ();
 sg13g2_fill_2 FILLER_75_734 ();
 sg13g2_decap_8 FILLER_75_745 ();
 sg13g2_decap_8 FILLER_75_752 ();
 sg13g2_decap_8 FILLER_75_759 ();
 sg13g2_decap_8 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_773 ();
 sg13g2_decap_8 FILLER_75_780 ();
 sg13g2_decap_8 FILLER_75_787 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_8 FILLER_75_822 ();
 sg13g2_decap_8 FILLER_75_829 ();
 sg13g2_decap_8 FILLER_75_836 ();
 sg13g2_decap_8 FILLER_75_843 ();
 sg13g2_decap_8 FILLER_75_850 ();
 sg13g2_decap_4 FILLER_75_857 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_161 ();
 sg13g2_fill_2 FILLER_76_173 ();
 sg13g2_decap_8 FILLER_76_180 ();
 sg13g2_decap_8 FILLER_76_187 ();
 sg13g2_decap_4 FILLER_76_194 ();
 sg13g2_fill_1 FILLER_76_198 ();
 sg13g2_decap_4 FILLER_76_210 ();
 sg13g2_fill_2 FILLER_76_214 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_4 FILLER_76_231 ();
 sg13g2_fill_1 FILLER_76_243 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_decap_8 FILLER_76_256 ();
 sg13g2_decap_8 FILLER_76_263 ();
 sg13g2_decap_4 FILLER_76_270 ();
 sg13g2_fill_2 FILLER_76_274 ();
 sg13g2_fill_2 FILLER_76_281 ();
 sg13g2_fill_1 FILLER_76_283 ();
 sg13g2_decap_8 FILLER_76_289 ();
 sg13g2_decap_8 FILLER_76_320 ();
 sg13g2_decap_8 FILLER_76_327 ();
 sg13g2_decap_8 FILLER_76_334 ();
 sg13g2_fill_1 FILLER_76_341 ();
 sg13g2_fill_1 FILLER_76_347 ();
 sg13g2_fill_1 FILLER_76_361 ();
 sg13g2_fill_2 FILLER_76_376 ();
 sg13g2_fill_1 FILLER_76_378 ();
 sg13g2_decap_4 FILLER_76_384 ();
 sg13g2_fill_1 FILLER_76_388 ();
 sg13g2_fill_2 FILLER_76_394 ();
 sg13g2_fill_1 FILLER_76_396 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_2 FILLER_76_429 ();
 sg13g2_fill_1 FILLER_76_453 ();
 sg13g2_decap_4 FILLER_76_459 ();
 sg13g2_fill_1 FILLER_76_463 ();
 sg13g2_fill_2 FILLER_76_472 ();
 sg13g2_fill_1 FILLER_76_481 ();
 sg13g2_fill_1 FILLER_76_492 ();
 sg13g2_fill_2 FILLER_76_513 ();
 sg13g2_fill_1 FILLER_76_515 ();
 sg13g2_decap_8 FILLER_76_543 ();
 sg13g2_decap_8 FILLER_76_550 ();
 sg13g2_decap_8 FILLER_76_557 ();
 sg13g2_decap_8 FILLER_76_564 ();
 sg13g2_decap_8 FILLER_76_571 ();
 sg13g2_decap_8 FILLER_76_578 ();
 sg13g2_fill_2 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_591 ();
 sg13g2_decap_8 FILLER_76_598 ();
 sg13g2_decap_8 FILLER_76_618 ();
 sg13g2_decap_8 FILLER_76_625 ();
 sg13g2_decap_8 FILLER_76_632 ();
 sg13g2_decap_8 FILLER_76_639 ();
 sg13g2_decap_8 FILLER_76_646 ();
 sg13g2_decap_8 FILLER_76_653 ();
 sg13g2_decap_8 FILLER_76_660 ();
 sg13g2_decap_8 FILLER_76_667 ();
 sg13g2_decap_8 FILLER_76_674 ();
 sg13g2_decap_8 FILLER_76_681 ();
 sg13g2_decap_8 FILLER_76_688 ();
 sg13g2_decap_8 FILLER_76_695 ();
 sg13g2_decap_8 FILLER_76_702 ();
 sg13g2_decap_8 FILLER_76_709 ();
 sg13g2_decap_8 FILLER_76_716 ();
 sg13g2_decap_8 FILLER_76_723 ();
 sg13g2_decap_8 FILLER_76_730 ();
 sg13g2_decap_8 FILLER_76_737 ();
 sg13g2_decap_8 FILLER_76_744 ();
 sg13g2_decap_8 FILLER_76_751 ();
 sg13g2_decap_8 FILLER_76_758 ();
 sg13g2_decap_8 FILLER_76_765 ();
 sg13g2_decap_8 FILLER_76_772 ();
 sg13g2_decap_8 FILLER_76_779 ();
 sg13g2_decap_8 FILLER_76_786 ();
 sg13g2_decap_8 FILLER_76_793 ();
 sg13g2_decap_8 FILLER_76_800 ();
 sg13g2_decap_8 FILLER_76_807 ();
 sg13g2_decap_8 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_821 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_4 FILLER_76_856 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_fill_2 FILLER_77_154 ();
 sg13g2_fill_1 FILLER_77_156 ();
 sg13g2_fill_1 FILLER_77_183 ();
 sg13g2_fill_2 FILLER_77_205 ();
 sg13g2_fill_2 FILLER_77_228 ();
 sg13g2_decap_4 FILLER_77_252 ();
 sg13g2_decap_4 FILLER_77_296 ();
 sg13g2_fill_1 FILLER_77_300 ();
 sg13g2_decap_4 FILLER_77_305 ();
 sg13g2_decap_8 FILLER_77_313 ();
 sg13g2_decap_8 FILLER_77_320 ();
 sg13g2_decap_8 FILLER_77_327 ();
 sg13g2_decap_4 FILLER_77_334 ();
 sg13g2_fill_2 FILLER_77_338 ();
 sg13g2_decap_8 FILLER_77_356 ();
 sg13g2_decap_8 FILLER_77_363 ();
 sg13g2_decap_4 FILLER_77_370 ();
 sg13g2_fill_1 FILLER_77_374 ();
 sg13g2_fill_2 FILLER_77_405 ();
 sg13g2_fill_1 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_77_426 ();
 sg13g2_decap_4 FILLER_77_433 ();
 sg13g2_fill_2 FILLER_77_437 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_472 ();
 sg13g2_decap_4 FILLER_77_479 ();
 sg13g2_fill_1 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_495 ();
 sg13g2_decap_4 FILLER_77_502 ();
 sg13g2_fill_1 FILLER_77_506 ();
 sg13g2_decap_4 FILLER_77_512 ();
 sg13g2_fill_2 FILLER_77_516 ();
 sg13g2_decap_8 FILLER_77_545 ();
 sg13g2_decap_8 FILLER_77_552 ();
 sg13g2_decap_8 FILLER_77_559 ();
 sg13g2_decap_8 FILLER_77_566 ();
 sg13g2_decap_8 FILLER_77_573 ();
 sg13g2_decap_8 FILLER_77_580 ();
 sg13g2_decap_8 FILLER_77_587 ();
 sg13g2_decap_8 FILLER_77_594 ();
 sg13g2_decap_8 FILLER_77_601 ();
 sg13g2_decap_8 FILLER_77_608 ();
 sg13g2_decap_8 FILLER_77_615 ();
 sg13g2_decap_8 FILLER_77_622 ();
 sg13g2_decap_8 FILLER_77_629 ();
 sg13g2_decap_8 FILLER_77_636 ();
 sg13g2_decap_8 FILLER_77_643 ();
 sg13g2_decap_8 FILLER_77_650 ();
 sg13g2_decap_8 FILLER_77_657 ();
 sg13g2_decap_8 FILLER_77_664 ();
 sg13g2_decap_8 FILLER_77_671 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_decap_8 FILLER_77_685 ();
 sg13g2_decap_8 FILLER_77_692 ();
 sg13g2_decap_8 FILLER_77_699 ();
 sg13g2_decap_8 FILLER_77_706 ();
 sg13g2_decap_8 FILLER_77_713 ();
 sg13g2_decap_8 FILLER_77_720 ();
 sg13g2_decap_8 FILLER_77_727 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_decap_8 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_776 ();
 sg13g2_decap_8 FILLER_77_783 ();
 sg13g2_decap_8 FILLER_77_790 ();
 sg13g2_decap_8 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_decap_8 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_832 ();
 sg13g2_decap_8 FILLER_77_839 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_4 FILLER_78_184 ();
 sg13g2_fill_2 FILLER_78_188 ();
 sg13g2_decap_8 FILLER_78_202 ();
 sg13g2_decap_8 FILLER_78_209 ();
 sg13g2_fill_1 FILLER_78_216 ();
 sg13g2_fill_2 FILLER_78_226 ();
 sg13g2_fill_2 FILLER_78_242 ();
 sg13g2_fill_1 FILLER_78_244 ();
 sg13g2_decap_8 FILLER_78_250 ();
 sg13g2_decap_8 FILLER_78_257 ();
 sg13g2_decap_8 FILLER_78_264 ();
 sg13g2_fill_1 FILLER_78_279 ();
 sg13g2_fill_2 FILLER_78_285 ();
 sg13g2_fill_1 FILLER_78_287 ();
 sg13g2_fill_2 FILLER_78_293 ();
 sg13g2_fill_2 FILLER_78_303 ();
 sg13g2_fill_2 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_4 FILLER_78_357 ();
 sg13g2_fill_2 FILLER_78_361 ();
 sg13g2_decap_4 FILLER_78_378 ();
 sg13g2_fill_1 FILLER_78_382 ();
 sg13g2_fill_2 FILLER_78_388 ();
 sg13g2_fill_1 FILLER_78_390 ();
 sg13g2_decap_4 FILLER_78_397 ();
 sg13g2_fill_2 FILLER_78_401 ();
 sg13g2_decap_4 FILLER_78_422 ();
 sg13g2_decap_4 FILLER_78_434 ();
 sg13g2_fill_2 FILLER_78_438 ();
 sg13g2_decap_4 FILLER_78_445 ();
 sg13g2_fill_1 FILLER_78_449 ();
 sg13g2_decap_4 FILLER_78_455 ();
 sg13g2_fill_1 FILLER_78_470 ();
 sg13g2_decap_4 FILLER_78_484 ();
 sg13g2_fill_2 FILLER_78_495 ();
 sg13g2_fill_1 FILLER_78_497 ();
 sg13g2_fill_2 FILLER_78_503 ();
 sg13g2_decap_8 FILLER_78_535 ();
 sg13g2_decap_8 FILLER_78_542 ();
 sg13g2_decap_8 FILLER_78_549 ();
 sg13g2_decap_8 FILLER_78_556 ();
 sg13g2_decap_8 FILLER_78_563 ();
 sg13g2_decap_8 FILLER_78_570 ();
 sg13g2_decap_8 FILLER_78_577 ();
 sg13g2_decap_8 FILLER_78_584 ();
 sg13g2_decap_8 FILLER_78_591 ();
 sg13g2_decap_8 FILLER_78_598 ();
 sg13g2_decap_8 FILLER_78_605 ();
 sg13g2_decap_8 FILLER_78_612 ();
 sg13g2_decap_8 FILLER_78_619 ();
 sg13g2_decap_8 FILLER_78_626 ();
 sg13g2_decap_8 FILLER_78_633 ();
 sg13g2_decap_8 FILLER_78_640 ();
 sg13g2_decap_8 FILLER_78_647 ();
 sg13g2_decap_8 FILLER_78_654 ();
 sg13g2_decap_8 FILLER_78_661 ();
 sg13g2_decap_8 FILLER_78_668 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_696 ();
 sg13g2_decap_8 FILLER_78_703 ();
 sg13g2_decap_8 FILLER_78_710 ();
 sg13g2_decap_8 FILLER_78_717 ();
 sg13g2_decap_8 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_731 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_752 ();
 sg13g2_decap_8 FILLER_78_759 ();
 sg13g2_decap_8 FILLER_78_766 ();
 sg13g2_decap_8 FILLER_78_773 ();
 sg13g2_decap_8 FILLER_78_780 ();
 sg13g2_decap_8 FILLER_78_787 ();
 sg13g2_decap_8 FILLER_78_794 ();
 sg13g2_decap_8 FILLER_78_801 ();
 sg13g2_decap_8 FILLER_78_808 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_decap_4 FILLER_78_857 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_4 FILLER_79_154 ();
 sg13g2_fill_2 FILLER_79_158 ();
 sg13g2_fill_2 FILLER_79_169 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_1 FILLER_79_176 ();
 sg13g2_fill_2 FILLER_79_182 ();
 sg13g2_fill_1 FILLER_79_184 ();
 sg13g2_fill_1 FILLER_79_189 ();
 sg13g2_fill_1 FILLER_79_216 ();
 sg13g2_fill_2 FILLER_79_274 ();
 sg13g2_fill_2 FILLER_79_289 ();
 sg13g2_fill_1 FILLER_79_291 ();
 sg13g2_decap_4 FILLER_79_297 ();
 sg13g2_fill_2 FILLER_79_314 ();
 sg13g2_decap_8 FILLER_79_320 ();
 sg13g2_fill_1 FILLER_79_327 ();
 sg13g2_decap_4 FILLER_79_332 ();
 sg13g2_fill_2 FILLER_79_362 ();
 sg13g2_fill_1 FILLER_79_364 ();
 sg13g2_decap_4 FILLER_79_373 ();
 sg13g2_fill_2 FILLER_79_399 ();
 sg13g2_fill_1 FILLER_79_448 ();
 sg13g2_fill_1 FILLER_79_461 ();
 sg13g2_fill_2 FILLER_79_467 ();
 sg13g2_fill_1 FILLER_79_469 ();
 sg13g2_fill_2 FILLER_79_475 ();
 sg13g2_decap_4 FILLER_79_510 ();
 sg13g2_decap_8 FILLER_79_526 ();
 sg13g2_decap_8 FILLER_79_533 ();
 sg13g2_decap_8 FILLER_79_540 ();
 sg13g2_decap_8 FILLER_79_547 ();
 sg13g2_decap_8 FILLER_79_554 ();
 sg13g2_decap_8 FILLER_79_561 ();
 sg13g2_decap_8 FILLER_79_568 ();
 sg13g2_decap_8 FILLER_79_575 ();
 sg13g2_decap_8 FILLER_79_582 ();
 sg13g2_decap_8 FILLER_79_589 ();
 sg13g2_decap_8 FILLER_79_596 ();
 sg13g2_decap_8 FILLER_79_603 ();
 sg13g2_decap_8 FILLER_79_610 ();
 sg13g2_decap_8 FILLER_79_617 ();
 sg13g2_decap_8 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_631 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_659 ();
 sg13g2_decap_8 FILLER_79_666 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_687 ();
 sg13g2_decap_8 FILLER_79_694 ();
 sg13g2_decap_8 FILLER_79_701 ();
 sg13g2_decap_8 FILLER_79_708 ();
 sg13g2_decap_8 FILLER_79_715 ();
 sg13g2_decap_8 FILLER_79_722 ();
 sg13g2_decap_8 FILLER_79_729 ();
 sg13g2_decap_8 FILLER_79_736 ();
 sg13g2_decap_8 FILLER_79_743 ();
 sg13g2_decap_8 FILLER_79_750 ();
 sg13g2_decap_8 FILLER_79_757 ();
 sg13g2_decap_8 FILLER_79_764 ();
 sg13g2_decap_8 FILLER_79_771 ();
 sg13g2_decap_8 FILLER_79_778 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_fill_1 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_191 ();
 sg13g2_fill_2 FILLER_80_198 ();
 sg13g2_fill_1 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_205 ();
 sg13g2_decap_8 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_decap_8 FILLER_80_230 ();
 sg13g2_fill_2 FILLER_80_237 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_fill_2 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_270 ();
 sg13g2_fill_2 FILLER_80_277 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_4 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_339 ();
 sg13g2_fill_1 FILLER_80_346 ();
 sg13g2_decap_8 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_358 ();
 sg13g2_fill_2 FILLER_80_364 ();
 sg13g2_fill_1 FILLER_80_366 ();
 sg13g2_fill_2 FILLER_80_377 ();
 sg13g2_fill_1 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_fill_2 FILLER_80_404 ();
 sg13g2_decap_4 FILLER_80_414 ();
 sg13g2_fill_1 FILLER_80_418 ();
 sg13g2_fill_2 FILLER_80_424 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_fill_2 FILLER_80_450 ();
 sg13g2_fill_1 FILLER_80_452 ();
 sg13g2_decap_4 FILLER_80_457 ();
 sg13g2_fill_2 FILLER_80_461 ();
 sg13g2_decap_4 FILLER_80_467 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_4 FILLER_80_493 ();
 sg13g2_fill_2 FILLER_80_497 ();
 sg13g2_decap_8 FILLER_80_509 ();
 sg13g2_decap_8 FILLER_80_516 ();
 sg13g2_decap_8 FILLER_80_523 ();
 sg13g2_decap_8 FILLER_80_530 ();
 sg13g2_decap_8 FILLER_80_537 ();
 sg13g2_decap_8 FILLER_80_544 ();
 sg13g2_decap_8 FILLER_80_551 ();
 sg13g2_decap_8 FILLER_80_558 ();
 sg13g2_decap_8 FILLER_80_565 ();
 sg13g2_decap_8 FILLER_80_572 ();
 sg13g2_decap_8 FILLER_80_579 ();
 sg13g2_decap_8 FILLER_80_586 ();
 sg13g2_decap_8 FILLER_80_593 ();
 sg13g2_decap_8 FILLER_80_600 ();
 sg13g2_decap_8 FILLER_80_607 ();
 sg13g2_decap_8 FILLER_80_614 ();
 sg13g2_decap_8 FILLER_80_621 ();
 sg13g2_decap_8 FILLER_80_628 ();
 sg13g2_decap_8 FILLER_80_635 ();
 sg13g2_decap_8 FILLER_80_642 ();
 sg13g2_decap_8 FILLER_80_649 ();
 sg13g2_decap_8 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_663 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_8 FILLER_80_677 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_decap_8 FILLER_80_691 ();
 sg13g2_decap_8 FILLER_80_698 ();
 sg13g2_decap_8 FILLER_80_705 ();
 sg13g2_decap_8 FILLER_80_712 ();
 sg13g2_decap_8 FILLER_80_719 ();
 sg13g2_decap_8 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_733 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_decap_8 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_754 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_decap_8 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_810 ();
 sg13g2_decap_8 FILLER_80_817 ();
 sg13g2_decap_8 FILLER_80_824 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_fill_2 FILLER_80_859 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net164;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule
