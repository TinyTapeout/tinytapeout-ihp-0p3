module tt_um_arud4172_ROOTS_vga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire clknet_0_clk;
 wire \color_index[0] ;
 wire \color_index[1] ;
 wire \color_index[2] ;
 wire dir_x;
 wire dir_y;
 wire \frame_counter[0] ;
 wire \frame_counter[1] ;
 wire \frame_counter[2] ;
 wire \frame_counter[3] ;
 wire \frame_counter[4] ;
 wire \frame_counter[5] ;
 wire \frame_counter[6] ;
 wire \frame_counter[7] ;
 wire \frame_divider[0] ;
 wire \frame_divider[1] ;
 wire hsync;
 wire \logo_left[0] ;
 wire \logo_left[1] ;
 wire \logo_left[2] ;
 wire \logo_left[3] ;
 wire \logo_left[4] ;
 wire \logo_left[5] ;
 wire \logo_left[6] ;
 wire \logo_left[7] ;
 wire \logo_left[8] ;
 wire \logo_left[9] ;
 wire \logo_top[0] ;
 wire \logo_top[1] ;
 wire \logo_top[2] ;
 wire \logo_top[3] ;
 wire \logo_top[4] ;
 wire \logo_top[5] ;
 wire \logo_top[6] ;
 wire \logo_top[7] ;
 wire \logo_top[8] ;
 wire \logo_top[9] ;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \prev_y[0] ;
 wire \prev_y[1] ;
 wire \prev_y[2] ;
 wire \prev_y[3] ;
 wire \prev_y[4] ;
 wire \prev_y[5] ;
 wire \prev_y[6] ;
 wire \prev_y[7] ;
 wire \prev_y[8] ;
 wire \prev_y[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire \vga_sync_gen.vsync ;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;

 sg13g2_inv_1 _3766_ (.Y(_0636_),
    .A(net141));
 sg13g2_inv_1 _3767_ (.Y(_0647_),
    .A(net96));
 sg13g2_inv_1 _3768_ (.Y(_0658_),
    .A(net2615));
 sg13g2_inv_2 _3769_ (.Y(_0669_),
    .A(net2617));
 sg13g2_inv_1 _3770_ (.Y(_0680_),
    .A(\logo_top[7] ));
 sg13g2_inv_1 _3771_ (.Y(_0691_),
    .A(\logo_top[6] ));
 sg13g2_inv_1 _3772_ (.Y(_0702_),
    .A(\logo_top[5] ));
 sg13g2_inv_1 _3773_ (.Y(_0713_),
    .A(\logo_top[4] ));
 sg13g2_inv_1 _3774_ (.Y(_0724_),
    .A(\logo_top[2] ));
 sg13g2_inv_1 _3775_ (.Y(_0735_),
    .A(\logo_top[0] ));
 sg13g2_inv_1 _3776_ (.Y(_0746_),
    .A(net104));
 sg13g2_inv_1 _3777_ (.Y(_0757_),
    .A(\logo_left[5] ));
 sg13g2_inv_1 _3778_ (.Y(_0768_),
    .A(net106));
 sg13g2_inv_1 _3779_ (.Y(_0779_),
    .A(\pix_x[8] ));
 sg13g2_inv_2 _3780_ (.Y(_0790_),
    .A(\pix_y[8] ));
 sg13g2_inv_1 _3781_ (.Y(_0801_),
    .A(net158));
 sg13g2_inv_2 _3782_ (.Y(_0812_),
    .A(\pix_y[7] ));
 sg13g2_inv_1 _3783_ (.Y(_0823_),
    .A(net2603));
 sg13g2_inv_1 _3784_ (.Y(_0834_),
    .A(net2607));
 sg13g2_inv_1 _3785_ (.Y(_0845_),
    .A(net2610));
 sg13g2_inv_1 _3786_ (.Y(_0856_),
    .A(net2612));
 sg13g2_inv_1 _3787_ (.Y(_0867_),
    .A(net2613));
 sg13g2_inv_1 _3788_ (.Y(_0878_),
    .A(net2628));
 sg13g2_inv_1 _3789_ (.Y(_0889_),
    .A(net123));
 sg13g2_inv_1 _3790_ (.Y(_0900_),
    .A(\prev_y[6] ));
 sg13g2_inv_1 _3791_ (.Y(_0911_),
    .A(\prev_y[8] ));
 sg13g2_inv_1 _3792_ (.Y(_0922_),
    .A(net109));
 sg13g2_inv_1 _3793_ (.Y(_0933_),
    .A(net2));
 sg13g2_inv_1 _3794_ (.Y(_0944_),
    .A(net3));
 sg13g2_inv_1 _3795_ (.Y(_0955_),
    .A(\frame_counter[3] ));
 sg13g2_nand2_1 _3796_ (.Y(_0966_),
    .A(\pix_y[8] ),
    .B(_0801_));
 sg13g2_nand2_1 _3797_ (.Y(_0977_),
    .A(net2608),
    .B(net2612));
 sg13g2_nor4_1 _3798_ (.A(net2607),
    .B(net2610),
    .C(_0966_),
    .D(_0977_),
    .Y(_0988_));
 sg13g2_and4_1 _3799_ (.A(net173),
    .B(net2603),
    .C(net2605),
    .D(_0988_),
    .X(_0001_));
 sg13g2_nand3_1 _3800_ (.B(net163),
    .C(\pix_x[4] ),
    .A(net2620),
    .Y(_1009_));
 sg13g2_nor3_1 _3801_ (.A(net136),
    .B(\pix_x[5] ),
    .C(\pix_x[4] ),
    .Y(_1020_));
 sg13g2_nand4_1 _3802_ (.B(net2619),
    .C(net134),
    .A(_0779_),
    .Y(_1031_),
    .D(_1009_));
 sg13g2_nor2_1 _3803_ (.A(net137),
    .B(_1031_),
    .Y(_0000_));
 sg13g2_nand2b_1 _3804_ (.Y(_1052_),
    .B(\logo_left[0] ),
    .A_N(\pix_x[0] ));
 sg13g2_nor2b_1 _3805_ (.A(\logo_left[1] ),
    .B_N(\pix_x[1] ),
    .Y(_1063_));
 sg13g2_xnor2_1 _3806_ (.Y(_1074_),
    .A(\logo_left[1] ),
    .B(\pix_x[1] ));
 sg13g2_xnor2_1 _3807_ (.Y(_1085_),
    .A(_1052_),
    .B(_1074_));
 sg13g2_nand2_1 _3808_ (.Y(_1096_),
    .A(_0724_),
    .B(net2611));
 sg13g2_xor2_1 _3809_ (.B(net2611),
    .A(\logo_top[2] ),
    .X(_1107_));
 sg13g2_nor2_1 _3810_ (.A(\logo_top[1] ),
    .B(_0856_),
    .Y(_1118_));
 sg13g2_nand2_2 _3811_ (.Y(_1129_),
    .A(\logo_top[0] ),
    .B(_0867_));
 sg13g2_xnor2_1 _3812_ (.Y(_1140_),
    .A(\logo_top[1] ),
    .B(\pix_y[1] ));
 sg13g2_a21oi_2 _3813_ (.B1(_1118_),
    .Y(_1151_),
    .A2(_1140_),
    .A1(_1129_));
 sg13g2_o21ai_1 _3814_ (.B1(_1096_),
    .Y(_1162_),
    .A1(_1107_),
    .A2(_1151_));
 sg13g2_nor2b_1 _3815_ (.A(\logo_top[3] ),
    .B_N(net2609),
    .Y(_1173_));
 sg13g2_xnor2_1 _3816_ (.Y(_1184_),
    .A(\logo_top[3] ),
    .B(net2609));
 sg13g2_xor2_1 _3817_ (.B(_1184_),
    .A(_1162_),
    .X(_1195_));
 sg13g2_xnor2_1 _3818_ (.Y(_1206_),
    .A(_1162_),
    .B(_1184_));
 sg13g2_xor2_1 _3819_ (.B(\pix_y[4] ),
    .A(\logo_top[4] ),
    .X(_1217_));
 sg13g2_a21oi_2 _3820_ (.B1(_1173_),
    .Y(_1228_),
    .A2(_1184_),
    .A1(_1162_));
 sg13g2_nor2_1 _3821_ (.A(_1217_),
    .B(_1228_),
    .Y(_1239_));
 sg13g2_xor2_1 _3822_ (.B(_1228_),
    .A(_1217_),
    .X(_1250_));
 sg13g2_xnor2_1 _3823_ (.Y(_1261_),
    .A(_1217_),
    .B(_1228_));
 sg13g2_xor2_1 _3824_ (.B(_1151_),
    .A(_1107_),
    .X(_1272_));
 sg13g2_xnor2_1 _3825_ (.Y(_1283_),
    .A(_1107_),
    .B(_1151_));
 sg13g2_nand2_2 _3826_ (.Y(_1294_),
    .A(_0735_),
    .B(\pix_y[0] ));
 sg13g2_and2_2 _3827_ (.A(_1129_),
    .B(_1294_),
    .X(_1305_));
 sg13g2_nand2_2 _3828_ (.Y(_1316_),
    .A(_1129_),
    .B(_1294_));
 sg13g2_xor2_1 _3829_ (.B(_1140_),
    .A(_1129_),
    .X(_1327_));
 sg13g2_xnor2_1 _3830_ (.Y(_1338_),
    .A(_1129_),
    .B(_1140_));
 sg13g2_nor2_1 _3831_ (.A(net2559),
    .B(net2538),
    .Y(_1349_));
 sg13g2_nand2_1 _3832_ (.Y(_1360_),
    .A(_1140_),
    .B(net2589));
 sg13g2_nand2_2 _3833_ (.Y(_1371_),
    .A(net2490),
    .B(net2463));
 sg13g2_nand2b_1 _3834_ (.Y(_1382_),
    .B(net2619),
    .A_N(\logo_left[7] ));
 sg13g2_xor2_1 _3835_ (.B(net2619),
    .A(\logo_left[7] ),
    .X(_1393_));
 sg13g2_nor2b_1 _3836_ (.A(\logo_left[6] ),
    .B_N(net2620),
    .Y(_1404_));
 sg13g2_xnor2_1 _3837_ (.Y(_1415_),
    .A(\logo_left[6] ),
    .B(net2620));
 sg13g2_nor2b_1 _3838_ (.A(\logo_left[5] ),
    .B_N(net2621),
    .Y(_1426_));
 sg13g2_xnor2_1 _3839_ (.Y(_1437_),
    .A(\logo_left[5] ),
    .B(net2621));
 sg13g2_nor2b_1 _3840_ (.A(\logo_left[4] ),
    .B_N(\pix_x[4] ),
    .Y(_1448_));
 sg13g2_a21oi_1 _3841_ (.A1(_1052_),
    .A2(_1074_),
    .Y(_1459_),
    .B1(_1063_));
 sg13g2_a21o_1 _3842_ (.A2(_1074_),
    .A1(_1052_),
    .B1(_1063_),
    .X(_1470_));
 sg13g2_nor2b_1 _3843_ (.A(net2618),
    .B_N(\pix_x[3] ),
    .Y(_1481_));
 sg13g2_nand2b_1 _3844_ (.Y(_1492_),
    .B(net2618),
    .A_N(\pix_x[3] ));
 sg13g2_xnor2_1 _3845_ (.Y(_1503_),
    .A(net2618),
    .B(\pix_x[3] ));
 sg13g2_nor2b_1 _3846_ (.A(\logo_left[2] ),
    .B_N(\pix_x[2] ),
    .Y(_1514_));
 sg13g2_xnor2_1 _3847_ (.Y(_1525_),
    .A(\logo_left[2] ),
    .B(\pix_x[2] ));
 sg13g2_nand2_1 _3848_ (.Y(_1536_),
    .A(_1503_),
    .B(_1525_));
 sg13g2_a21oi_1 _3849_ (.A1(_1492_),
    .A2(_1514_),
    .Y(_1547_),
    .B1(_1481_));
 sg13g2_o21ai_1 _3850_ (.B1(_1547_),
    .Y(_1558_),
    .A1(_1459_),
    .A2(_1536_));
 sg13g2_xnor2_1 _3851_ (.Y(_1569_),
    .A(\logo_left[4] ),
    .B(\pix_x[4] ));
 sg13g2_a21oi_1 _3852_ (.A1(_1558_),
    .A2(_1569_),
    .Y(_1580_),
    .B1(_1448_));
 sg13g2_a21o_1 _3853_ (.A2(_1569_),
    .A1(_1558_),
    .B1(_1448_),
    .X(_1591_));
 sg13g2_a21o_2 _3854_ (.A2(_1591_),
    .A1(_1437_),
    .B1(_1426_),
    .X(_1602_));
 sg13g2_a21oi_2 _3855_ (.B1(_1404_),
    .Y(_1613_),
    .A2(_1602_),
    .A1(_1415_));
 sg13g2_or2_1 _3856_ (.X(_1624_),
    .B(_1613_),
    .A(_1393_));
 sg13g2_xor2_1 _3857_ (.B(_1613_),
    .A(_1393_),
    .X(_1635_));
 sg13g2_xnor2_1 _3858_ (.Y(_1646_),
    .A(_1393_),
    .B(_1613_));
 sg13g2_xor2_1 _3859_ (.B(_1569_),
    .A(_1558_),
    .X(_1657_));
 sg13g2_xnor2_1 _3860_ (.Y(_1668_),
    .A(_1558_),
    .B(_1569_));
 sg13g2_a21oi_1 _3861_ (.A1(_1470_),
    .A2(_1525_),
    .Y(_1679_),
    .B1(_1514_));
 sg13g2_xnor2_1 _3862_ (.Y(_1690_),
    .A(_1503_),
    .B(_1679_));
 sg13g2_xor2_1 _3863_ (.B(_1679_),
    .A(_1503_),
    .X(_1701_));
 sg13g2_nor2_2 _3864_ (.A(net2455),
    .B(net2454),
    .Y(_1712_));
 sg13g2_nand2_1 _3865_ (.Y(_1723_),
    .A(net2458),
    .B(net2452));
 sg13g2_xor2_1 _3866_ (.B(_1602_),
    .A(_1415_),
    .X(_1734_));
 sg13g2_xnor2_1 _3867_ (.Y(_1745_),
    .A(_1415_),
    .B(_1602_));
 sg13g2_xnor2_1 _3868_ (.Y(_1756_),
    .A(_1437_),
    .B(_1580_));
 sg13g2_xnor2_1 _3869_ (.Y(_1767_),
    .A(_1437_),
    .B(_1591_));
 sg13g2_nor2_1 _3870_ (.A(net2451),
    .B(net2366),
    .Y(_1778_));
 sg13g2_nand2_1 _3871_ (.Y(_1789_),
    .A(net2453),
    .B(net2360));
 sg13g2_nor2_2 _3872_ (.A(net2269),
    .B(net2249),
    .Y(_1800_));
 sg13g2_nand2_2 _3873_ (.Y(_1811_),
    .A(net2286),
    .B(net2247));
 sg13g2_nor2_1 _3874_ (.A(net2458),
    .B(net2453),
    .Y(_1822_));
 sg13g2_nand2_1 _3875_ (.Y(_1833_),
    .A(net2455),
    .B(net2451));
 sg13g2_nor2_2 _3876_ (.A(net2452),
    .B(net2361),
    .Y(_1844_));
 sg13g2_nand2_2 _3877_ (.Y(_1855_),
    .A(net2454),
    .B(net2368));
 sg13g2_nor2_2 _3878_ (.A(net2375),
    .B(net2249),
    .Y(_1866_));
 sg13g2_o21ai_1 _3879_ (.B1(net2099),
    .Y(_1877_),
    .A1(net2375),
    .A2(_1811_));
 sg13g2_a21oi_2 _3880_ (.B1(net2146),
    .Y(_1888_),
    .A2(net2088),
    .A1(net2373));
 sg13g2_nor2_2 _3881_ (.A(net2453),
    .B(net2369),
    .Y(_1899_));
 sg13g2_nand2_1 _3882_ (.Y(_1910_),
    .A(net2451),
    .B(net2360));
 sg13g2_nor2_2 _3883_ (.A(net2270),
    .B(_1899_),
    .Y(_1921_));
 sg13g2_nand2_2 _3884_ (.Y(_1932_),
    .A(net2275),
    .B(net2241));
 sg13g2_nor2_2 _3885_ (.A(net2455),
    .B(net2451),
    .Y(_1943_));
 sg13g2_nand2_2 _3886_ (.Y(_1954_),
    .A(net2460),
    .B(net2454));
 sg13g2_nor2_1 _3887_ (.A(net2458),
    .B(net2451),
    .Y(_1965_));
 sg13g2_nand2_1 _3888_ (.Y(_1976_),
    .A(net2455),
    .B(net2454));
 sg13g2_xnor2_1 _3889_ (.Y(_1987_),
    .A(net2456),
    .B(net2454));
 sg13g2_xnor2_1 _3890_ (.Y(_1998_),
    .A(net2459),
    .B(net2453));
 sg13g2_nor2_1 _3891_ (.A(net2456),
    .B(net2260),
    .Y(_2009_));
 sg13g2_nand2_1 _3892_ (.Y(_2020_),
    .A(net2458),
    .B(net2277));
 sg13g2_nor2_2 _3893_ (.A(net2251),
    .B(net2362),
    .Y(_2031_));
 sg13g2_nor2_1 _3894_ (.A(net2458),
    .B(net2369),
    .Y(_2042_));
 sg13g2_nand2_1 _3895_ (.Y(_2053_),
    .A(net2456),
    .B(net2360));
 sg13g2_nand2_2 _3896_ (.Y(_2064_),
    .A(net2277),
    .B(net2236));
 sg13g2_nor2_2 _3897_ (.A(net2252),
    .B(net2238),
    .Y(_2075_));
 sg13g2_a21oi_2 _3898_ (.B1(net2090),
    .Y(_2086_),
    .A2(net2079),
    .A1(net2345));
 sg13g2_o21ai_1 _3899_ (.B1(net2137),
    .Y(_2097_),
    .A1(net2349),
    .A2(_2075_));
 sg13g2_nor2_1 _3900_ (.A(net2595),
    .B(net2530),
    .Y(_2108_));
 sg13g2_nand2_2 _3901_ (.Y(_2119_),
    .A(net2571),
    .B(net2549));
 sg13g2_nor2_1 _3902_ (.A(_1140_),
    .B(net2566),
    .Y(_2130_));
 sg13g2_nand2_1 _3903_ (.Y(_2141_),
    .A(net2578),
    .B(net2538));
 sg13g2_nor2_2 _3904_ (.A(net2595),
    .B(net2549),
    .Y(_2152_));
 sg13g2_nand2_1 _3905_ (.Y(_2163_),
    .A(net2564),
    .B(net2526));
 sg13g2_nor2_1 _3906_ (.A(net2478),
    .B(net2445),
    .Y(_2174_));
 sg13g2_nand2_2 _3907_ (.Y(_2185_),
    .A(net2465),
    .B(net2434));
 sg13g2_nor2_1 _3908_ (.A(net2459),
    .B(net2362),
    .Y(_2196_));
 sg13g2_nand2_2 _3909_ (.Y(_2207_),
    .A(_1668_),
    .B(net2370));
 sg13g2_nor2_1 _3910_ (.A(_1712_),
    .B(net2239),
    .Y(_2218_));
 sg13g2_a21oi_2 _3911_ (.B1(net2349),
    .Y(_2229_),
    .A2(net2362),
    .A1(net2455));
 sg13g2_o21ai_1 _3912_ (.B1(net2346),
    .Y(_2240_),
    .A1(net2459),
    .A2(net2366));
 sg13g2_nor2_2 _3913_ (.A(net2274),
    .B(_2240_),
    .Y(_2251_));
 sg13g2_nor2_2 _3914_ (.A(net2459),
    .B(net2256),
    .Y(_2262_));
 sg13g2_nand2_2 _3915_ (.Y(_2273_),
    .A(net2456),
    .B(net2280));
 sg13g2_nor2_1 _3916_ (.A(net2367),
    .B(net2357),
    .Y(_2284_));
 sg13g2_nand2_1 _3917_ (.Y(_2295_),
    .A(net2360),
    .B(net2358));
 sg13g2_nor2_2 _3918_ (.A(net2271),
    .B(net2231),
    .Y(_2306_));
 sg13g2_nand2_2 _3919_ (.Y(_2317_),
    .A(net2280),
    .B(net2232));
 sg13g2_nor3_2 _3920_ (.A(net2097),
    .B(_2251_),
    .C(_2306_),
    .Y(_2328_));
 sg13g2_nand3b_1 _3921_ (.B(net2078),
    .C(net2141),
    .Y(_2339_),
    .A_N(_2251_));
 sg13g2_nor2_2 _3922_ (.A(net2456),
    .B(net2360),
    .Y(_2350_));
 sg13g2_nand2_1 _3923_ (.Y(_2361_),
    .A(net2458),
    .B(net2369));
 sg13g2_nor2_2 _3924_ (.A(net2278),
    .B(net2228),
    .Y(_2372_));
 sg13g2_nand2_2 _3925_ (.Y(_2383_),
    .A(net2250),
    .B(net2226));
 sg13g2_nor2_2 _3926_ (.A(net2140),
    .B(_2383_),
    .Y(_2394_));
 sg13g2_nand2_1 _3927_ (.Y(_2405_),
    .A(net2103),
    .B(net2077));
 sg13g2_nor2_2 _3928_ (.A(net2289),
    .B(net2245),
    .Y(_2416_));
 sg13g2_nand2_2 _3929_ (.Y(_2427_),
    .A(net2252),
    .B(_1855_));
 sg13g2_nor2_2 _3930_ (.A(net2174),
    .B(_2427_),
    .Y(_2438_));
 sg13g2_o21ai_1 _3931_ (.B1(net2092),
    .Y(_2449_),
    .A1(net2349),
    .A2(net2077));
 sg13g2_a21oi_2 _3932_ (.B1(net2133),
    .Y(_2460_),
    .A2(_2383_),
    .A1(net2345));
 sg13g2_o21ai_1 _3933_ (.B1(net2344),
    .Y(_2471_),
    .A1(_2328_),
    .A2(_2460_));
 sg13g2_nand2_1 _3934_ (.Y(_2482_),
    .A(net2050),
    .B(_2449_));
 sg13g2_nand2_1 _3935_ (.Y(_2493_),
    .A(net2538),
    .B(_2482_));
 sg13g2_o21ai_1 _3936_ (.B1(net2470),
    .Y(_2504_),
    .A1(_1888_),
    .A2(_2086_));
 sg13g2_nand4_1 _3937_ (.B(_2471_),
    .C(_2493_),
    .A(net2483),
    .Y(_2515_),
    .D(_2504_));
 sg13g2_nor2_1 _3938_ (.A(net2487),
    .B(net2544),
    .Y(_2526_));
 sg13g2_nand2_2 _3939_ (.Y(_2537_),
    .A(net2501),
    .B(net2521));
 sg13g2_nand2_2 _3940_ (.Y(_2548_),
    .A(net2285),
    .B(net2239));
 sg13g2_nor2_2 _3941_ (.A(net2459),
    .B(net2277),
    .Y(_2559_));
 sg13g2_nand2_2 _3942_ (.Y(_2570_),
    .A(net2455),
    .B(net2251));
 sg13g2_o21ai_1 _3943_ (.B1(_1833_),
    .Y(_2581_),
    .A1(net2459),
    .A2(net2364));
 sg13g2_a21oi_2 _3944_ (.B1(net2358),
    .Y(_2592_),
    .A2(net2366),
    .A1(net2455));
 sg13g2_nor2_1 _3945_ (.A(net2275),
    .B(_2592_),
    .Y(_2603_));
 sg13g2_nand2_2 _3946_ (.Y(_2614_),
    .A(net2258),
    .B(_2581_));
 sg13g2_nor2_2 _3947_ (.A(net2100),
    .B(_2603_),
    .Y(_2625_));
 sg13g2_nand3_1 _3948_ (.B(_2548_),
    .C(_2614_),
    .A(net2143),
    .Y(_2636_));
 sg13g2_nor2_2 _3949_ (.A(net2142),
    .B(net2254),
    .Y(_2647_));
 sg13g2_nor2_1 _3950_ (.A(net2457),
    .B(net2372),
    .Y(_2658_));
 sg13g2_nand2_2 _3951_ (.Y(_2669_),
    .A(net2458),
    .B(net2361));
 sg13g2_nor2_2 _3952_ (.A(net2375),
    .B(net2224),
    .Y(_2680_));
 sg13g2_nor2_2 _3953_ (.A(net2270),
    .B(net2225),
    .Y(_2691_));
 sg13g2_nand2_2 _3954_ (.Y(_2702_),
    .A(net2275),
    .B(_2669_));
 sg13g2_nor2_2 _3955_ (.A(net2140),
    .B(_2702_),
    .Y(_2713_));
 sg13g2_nand2_2 _3956_ (.Y(_2724_),
    .A(net2122),
    .B(_2691_));
 sg13g2_nand3_1 _3957_ (.B(net2275),
    .C(_2680_),
    .A(net2096),
    .Y(_2734_));
 sg13g2_nand4_1 _3958_ (.B(net2046),
    .C(net2044),
    .A(net2502),
    .Y(_2744_),
    .D(_2734_));
 sg13g2_o21ai_1 _3959_ (.B1(net2133),
    .Y(_2750_),
    .A1(_2031_),
    .A2(_2592_));
 sg13g2_nor2_1 _3960_ (.A(net2361),
    .B(net2355),
    .Y(_2757_));
 sg13g2_nand2_2 _3961_ (.Y(_2767_),
    .A(net2367),
    .B(net2356));
 sg13g2_nand2_2 _3962_ (.Y(_2778_),
    .A(net2253),
    .B(net2222));
 sg13g2_nor2_2 _3963_ (.A(net2274),
    .B(net2223),
    .Y(_2787_));
 sg13g2_nor2_2 _3964_ (.A(net2145),
    .B(_2778_),
    .Y(_2797_));
 sg13g2_nand2_2 _3965_ (.Y(_2806_),
    .A(net2089),
    .B(_2787_));
 sg13g2_nor2_2 _3966_ (.A(net2261),
    .B(net2359),
    .Y(_2816_));
 sg13g2_nand2_2 _3967_ (.Y(_2826_),
    .A(net2277),
    .B(net2357));
 sg13g2_nor2_2 _3968_ (.A(net2371),
    .B(net2355),
    .Y(_2836_));
 sg13g2_nand2_1 _3969_ (.Y(_2844_),
    .A(net2364),
    .B(_1943_));
 sg13g2_nor3_2 _3970_ (.A(net2264),
    .B(net2358),
    .C(_2836_),
    .Y(_2853_));
 sg13g2_o21ai_1 _3971_ (.B1(net2089),
    .Y(_2863_),
    .A1(_2787_),
    .A2(_2853_));
 sg13g2_and2_1 _3972_ (.A(net2580),
    .B(_2863_),
    .X(_2872_));
 sg13g2_nand2_1 _3973_ (.Y(_2882_),
    .A(_2750_),
    .B(_2872_));
 sg13g2_and2_1 _3974_ (.A(net2559),
    .B(net2044),
    .X(_2892_));
 sg13g2_nor2_2 _3975_ (.A(net2455),
    .B(net2279),
    .Y(_2901_));
 sg13g2_nand2_2 _3976_ (.Y(_2912_),
    .A(net2458),
    .B(net2256));
 sg13g2_nor2_2 _3977_ (.A(net2277),
    .B(net2222),
    .Y(_2922_));
 sg13g2_nand2_1 _3978_ (.Y(_2931_),
    .A(net2269),
    .B(_2757_));
 sg13g2_nor2_2 _3979_ (.A(net2174),
    .B(_2922_),
    .Y(_2936_));
 sg13g2_nand2_2 _3980_ (.Y(_2941_),
    .A(net2121),
    .B(_2931_));
 sg13g2_nor2_2 _3981_ (.A(net2453),
    .B(net2361),
    .Y(_2948_));
 sg13g2_nand2_1 _3982_ (.Y(_2954_),
    .A(net2451),
    .B(net2366));
 sg13g2_xnor2_1 _3983_ (.Y(_2963_),
    .A(net2453),
    .B(net2366));
 sg13g2_xnor2_1 _3984_ (.Y(_2972_),
    .A(net2451),
    .B(net2366));
 sg13g2_nor2_2 _3985_ (.A(net2375),
    .B(net2362),
    .Y(_2982_));
 sg13g2_nand2_2 _3986_ (.Y(_2991_),
    .A(net2364),
    .B(_1954_));
 sg13g2_nor2_2 _3987_ (.A(net2371),
    .B(_1943_),
    .Y(_2999_));
 sg13g2_nor2_2 _3988_ (.A(_1668_),
    .B(net2217),
    .Y(_3007_));
 sg13g2_nand2_2 _3989_ (.Y(_3011_),
    .A(net2460),
    .B(_2972_));
 sg13g2_o21ai_1 _3990_ (.B1(_2936_),
    .Y(_3012_),
    .A1(net2261),
    .A2(_3011_));
 sg13g2_a21oi_1 _3991_ (.A1(_2892_),
    .A2(_3012_),
    .Y(_3013_),
    .B1(net2538));
 sg13g2_a22oi_1 _3992_ (.Y(_3014_),
    .B1(_2882_),
    .B2(_3013_),
    .A2(_2744_),
    .A1(net2336));
 sg13g2_nor2_2 _3993_ (.A(net2487),
    .B(net2527),
    .Y(_3015_));
 sg13g2_nand2_2 _3994_ (.Y(_3016_),
    .A(net2501),
    .B(net2538));
 sg13g2_nor2_2 _3995_ (.A(net2364),
    .B(_1833_),
    .Y(_3017_));
 sg13g2_nand2_2 _3996_ (.Y(_3018_),
    .A(net2370),
    .B(net2359));
 sg13g2_nor2_2 _3997_ (.A(net2290),
    .B(_3017_),
    .Y(_3019_));
 sg13g2_o21ai_1 _3998_ (.B1(_1954_),
    .Y(_3020_),
    .A1(net2457),
    .A2(net2370));
 sg13g2_nand2_2 _3999_ (.Y(_3021_),
    .A(net2251),
    .B(_2240_));
 sg13g2_nor3_2 _4000_ (.A(net2275),
    .B(_2229_),
    .C(net2224),
    .Y(_3022_));
 sg13g2_nand3_1 _4001_ (.B(_2240_),
    .C(_2669_),
    .A(net2251),
    .Y(_3023_));
 sg13g2_nor2_2 _4002_ (.A(net2559),
    .B(net2089),
    .Y(_3024_));
 sg13g2_nand2_2 _4003_ (.Y(_3025_),
    .A(net2579),
    .B(net2138));
 sg13g2_nor2_2 _4004_ (.A(net2130),
    .B(_3022_),
    .Y(_3026_));
 sg13g2_nor2_2 _4005_ (.A(net2587),
    .B(net2109),
    .Y(_3027_));
 sg13g2_nand2_2 _4006_ (.Y(_3028_),
    .A(net2559),
    .B(net2140));
 sg13g2_nand2_2 _4007_ (.Y(_3029_),
    .A(net2256),
    .B(net2349));
 sg13g2_and2_2 _4008_ (.A(net2135),
    .B(net2074),
    .X(_3030_));
 sg13g2_nand2_2 _4009_ (.Y(_3031_),
    .A(net2139),
    .B(net2074));
 sg13g2_nand2_1 _4010_ (.Y(_3032_),
    .A(net2560),
    .B(_3030_));
 sg13g2_nor2_2 _4011_ (.A(net2136),
    .B(net2081),
    .Y(_3033_));
 sg13g2_nand2_2 _4012_ (.Y(_3034_),
    .A(net2089),
    .B(net2080));
 sg13g2_o21ai_1 _4013_ (.B1(net2093),
    .Y(_3035_),
    .A1(net2249),
    .A2(_2020_));
 sg13g2_a21oi_1 _4014_ (.A1(net2247),
    .A2(net2081),
    .Y(_3036_),
    .B1(net2139));
 sg13g2_a21oi_1 _4015_ (.A1(net2579),
    .A2(_3026_),
    .Y(_3037_),
    .B1(_3036_));
 sg13g2_a21oi_1 _4016_ (.A1(_3032_),
    .A2(_3037_),
    .Y(_3038_),
    .B1(net2330));
 sg13g2_nor2_2 _4017_ (.A(net2508),
    .B(net2526),
    .Y(_3039_));
 sg13g2_nand2_2 _4018_ (.Y(_3040_),
    .A(net2487),
    .B(net2547));
 sg13g2_a21oi_1 _4019_ (.A1(net2081),
    .A2(net2217),
    .Y(_3041_),
    .B1(net2149));
 sg13g2_o21ai_1 _4020_ (.B1(net2102),
    .Y(_3042_),
    .A1(net2080),
    .A2(net2216));
 sg13g2_o21ai_1 _4021_ (.B1(net2585),
    .Y(_3043_),
    .A1(net2045),
    .A2(_3041_));
 sg13g2_nor2_2 _4022_ (.A(net2094),
    .B(_2559_),
    .Y(_3044_));
 sg13g2_nand2_2 _4023_ (.Y(_3045_),
    .A(net2138),
    .B(_2570_));
 sg13g2_nor2_1 _4024_ (.A(_3041_),
    .B(_3044_),
    .Y(_3046_));
 sg13g2_a21oi_1 _4025_ (.A1(_3043_),
    .A2(_3046_),
    .Y(_3047_),
    .B1(net2325));
 sg13g2_nand2_1 _4026_ (.Y(_3048_),
    .A(net2498),
    .B(net2599));
 sg13g2_nor2_1 _4027_ (.A(net2517),
    .B(net2555),
    .Y(_3049_));
 sg13g2_nand2_1 _4028_ (.Y(_3050_),
    .A(net2499),
    .B(net2535));
 sg13g2_nor2_1 _4029_ (.A(net2508),
    .B(net2462),
    .Y(_3051_));
 sg13g2_nand2_2 _4030_ (.Y(_3052_),
    .A(net2483),
    .B(net2470));
 sg13g2_o21ai_1 _4031_ (.B1(net2102),
    .Y(_3053_),
    .A1(net2080),
    .A2(_2948_));
 sg13g2_a21oi_2 _4032_ (.B1(net2148),
    .Y(_3054_),
    .A2(net2220),
    .A1(net2082));
 sg13g2_nand3_1 _4033_ (.B(net2346),
    .C(net2226),
    .A(net2256),
    .Y(_3055_));
 sg13g2_and2_1 _4034_ (.A(net2149),
    .B(_3055_),
    .X(_3056_));
 sg13g2_nand2_2 _4035_ (.Y(_3057_),
    .A(net2149),
    .B(_3055_));
 sg13g2_a21oi_1 _4036_ (.A1(_3053_),
    .A2(_3057_),
    .Y(_3058_),
    .B1(net2462));
 sg13g2_a21oi_1 _4037_ (.A1(_3053_),
    .A2(_3057_),
    .Y(_3059_),
    .B1(_3052_));
 sg13g2_nor2_2 _4038_ (.A(_3036_),
    .B(_3044_),
    .Y(_3060_));
 sg13g2_nor2_2 _4039_ (.A(net2507),
    .B(net2402),
    .Y(_3061_));
 sg13g2_nand2_2 _4040_ (.Y(_3062_),
    .A(net2488),
    .B(net2409));
 sg13g2_o21ai_1 _4041_ (.B1(_3061_),
    .Y(_3063_),
    .A1(net2045),
    .A2(_3041_));
 sg13g2_nor2_1 _4042_ (.A(net2295),
    .B(_3014_),
    .Y(_3064_));
 sg13g2_o21ai_1 _4043_ (.B1(_3063_),
    .Y(_3065_),
    .A1(net2336),
    .A2(_3060_));
 sg13g2_nor4_2 _4044_ (.A(_3038_),
    .B(_3047_),
    .C(_3059_),
    .Y(_3066_),
    .D(_3065_));
 sg13g2_o21ai_1 _4045_ (.B1(net2376),
    .Y(_3067_),
    .A1(net2301),
    .A2(_3066_));
 sg13g2_a21oi_1 _4046_ (.A1(_2515_),
    .A2(_3064_),
    .Y(_3068_),
    .B1(_3067_));
 sg13g2_xor2_1 _4047_ (.B(net2606),
    .A(\logo_top[5] ),
    .X(_3069_));
 sg13g2_a21oi_2 _4048_ (.B1(_1239_),
    .Y(_3070_),
    .A2(net2607),
    .A1(_0713_));
 sg13g2_nor2_1 _4049_ (.A(_3069_),
    .B(_3070_),
    .Y(_3071_));
 sg13g2_xor2_1 _4050_ (.B(_3070_),
    .A(_3069_),
    .X(_3072_));
 sg13g2_xnor2_1 _4051_ (.Y(_3073_),
    .A(_3069_),
    .B(_3070_));
 sg13g2_nor2_2 _4052_ (.A(net2091),
    .B(net2075),
    .Y(_3074_));
 sg13g2_nand2_2 _4053_ (.Y(_3075_),
    .A(net2137),
    .B(_2912_));
 sg13g2_nor2_2 _4054_ (.A(net2363),
    .B(net2353),
    .Y(_3076_));
 sg13g2_nand2_2 _4055_ (.Y(_3077_),
    .A(net2370),
    .B(net2351));
 sg13g2_nor2_2 _4056_ (.A(net2363),
    .B(net2350),
    .Y(_3078_));
 sg13g2_nand2_2 _4057_ (.Y(_3079_),
    .A(net2367),
    .B(net2346));
 sg13g2_a21oi_1 _4058_ (.A1(net2273),
    .A2(_3079_),
    .Y(_3080_),
    .B1(net2135));
 sg13g2_nand2_2 _4059_ (.Y(_3081_),
    .A(net2460),
    .B(net2218));
 sg13g2_o21ai_1 _4060_ (.B1(net2247),
    .Y(_3082_),
    .A1(net2362),
    .A2(net2345));
 sg13g2_a21o_2 _4061_ (.A2(_3082_),
    .A1(net2273),
    .B1(net2136),
    .X(_3083_));
 sg13g2_a21oi_1 _4062_ (.A1(net2273),
    .A2(_3082_),
    .Y(_3084_),
    .B1(net2136));
 sg13g2_nor2_2 _4063_ (.A(net2118),
    .B(net2285),
    .Y(_3085_));
 sg13g2_nand2_1 _4064_ (.Y(_3086_),
    .A(net2136),
    .B(net2075));
 sg13g2_a21oi_1 _4065_ (.A1(_3075_),
    .A2(_3083_),
    .Y(_3087_),
    .B1(net2429));
 sg13g2_o21ai_1 _4066_ (.B1(net2153),
    .Y(_3088_),
    .A1(net2245),
    .A2(net2074));
 sg13g2_nor2_2 _4067_ (.A(net2416),
    .B(_3088_),
    .Y(_3089_));
 sg13g2_nor2_2 _4068_ (.A(net2571),
    .B(net2166),
    .Y(_3090_));
 sg13g2_nand2_2 _4069_ (.Y(_3091_),
    .A(net2586),
    .B(net2102));
 sg13g2_nor3_2 _4070_ (.A(net2250),
    .B(net2358),
    .C(net2223),
    .Y(_3092_));
 sg13g2_nor2_2 _4071_ (.A(net2134),
    .B(_3092_),
    .Y(_3093_));
 sg13g2_nor3_1 _4072_ (.A(net2134),
    .B(net2416),
    .C(_3092_),
    .Y(_3094_));
 sg13g2_nor2_2 _4073_ (.A(net2093),
    .B(net2074),
    .Y(_3095_));
 sg13g2_o21ai_1 _4074_ (.B1(net2319),
    .Y(_3096_),
    .A1(_3030_),
    .A2(_3093_));
 sg13g2_nor2_2 _4075_ (.A(net2136),
    .B(_2262_),
    .Y(_3097_));
 sg13g2_nand2_2 _4076_ (.Y(_3098_),
    .A(net2104),
    .B(_2273_));
 sg13g2_nor2_2 _4077_ (.A(net2279),
    .B(net2235),
    .Y(_3099_));
 sg13g2_nand2_2 _4078_ (.Y(_3100_),
    .A(net2250),
    .B(net2234));
 sg13g2_nor2_2 _4079_ (.A(net2285),
    .B(net2354),
    .Y(_3101_));
 sg13g2_nand2_2 _4080_ (.Y(_3102_),
    .A(net2268),
    .B(net2352));
 sg13g2_nand3_1 _4081_ (.B(net2352),
    .C(net2234),
    .A(net2252),
    .Y(_3103_));
 sg13g2_and2_2 _4082_ (.A(net2133),
    .B(_3103_),
    .X(_3104_));
 sg13g2_o21ai_1 _4083_ (.B1(net2578),
    .Y(_3105_),
    .A1(_3097_),
    .A2(_3104_));
 sg13g2_o21ai_1 _4084_ (.B1(net2421),
    .Y(_3106_),
    .A1(_3097_),
    .A2(_3104_));
 sg13g2_a21oi_1 _4085_ (.A1(_3075_),
    .A2(_3098_),
    .Y(_3107_),
    .B1(net2539));
 sg13g2_o21ai_1 _4086_ (.B1(net2521),
    .Y(_3108_),
    .A1(net2034),
    .A2(_3097_));
 sg13g2_a22oi_1 _4087_ (.Y(_3109_),
    .B1(_3085_),
    .B2(net2347),
    .A2(_2713_),
    .A1(net2373));
 sg13g2_nand2_1 _4088_ (.Y(_3110_),
    .A(net2439),
    .B(_3109_));
 sg13g2_and4_1 _4089_ (.A(net2501),
    .B(_3106_),
    .C(_3108_),
    .D(_3110_),
    .X(_3111_));
 sg13g2_nor4_1 _4090_ (.A(net2501),
    .B(_3087_),
    .C(_3089_),
    .D(_3094_),
    .Y(_3112_));
 sg13g2_o21ai_1 _4091_ (.B1(_3096_),
    .Y(_3113_),
    .A1(_3111_),
    .A2(_3112_));
 sg13g2_nand3_1 _4092_ (.B(net2237),
    .C(_2767_),
    .A(net2291),
    .Y(_3114_));
 sg13g2_nand2b_2 _4093_ (.Y(_3115_),
    .B(net2124),
    .A_N(_3114_));
 sg13g2_nor2_2 _4094_ (.A(net2276),
    .B(_2948_),
    .Y(_3116_));
 sg13g2_nand2_2 _4095_ (.Y(_3117_),
    .A(net2269),
    .B(net2219));
 sg13g2_nand2_2 _4096_ (.Y(_3118_),
    .A(net2174),
    .B(_2372_));
 sg13g2_nor2_1 _4097_ (.A(net2286),
    .B(_3076_),
    .Y(_3119_));
 sg13g2_nand2_1 _4098_ (.Y(_3120_),
    .A(net2160),
    .B(net2067));
 sg13g2_nor2_2 _4099_ (.A(net2373),
    .B(net2368),
    .Y(_3121_));
 sg13g2_nand2_2 _4100_ (.Y(_3122_),
    .A(net2375),
    .B(net2362));
 sg13g2_nor2_1 _4101_ (.A(net2268),
    .B(_3121_),
    .Y(_3123_));
 sg13g2_nand2_2 _4102_ (.Y(_3124_),
    .A(net2285),
    .B(_3122_));
 sg13g2_nor2_2 _4103_ (.A(net2113),
    .B(net2066),
    .Y(_3125_));
 sg13g2_nor2_1 _4104_ (.A(net2364),
    .B(net2352),
    .Y(_3126_));
 sg13g2_nand2_1 _4105_ (.Y(_3127_),
    .A(net2372),
    .B(net2354));
 sg13g2_nor2_1 _4106_ (.A(net2285),
    .B(net2213),
    .Y(_3128_));
 sg13g2_nand2_2 _4107_ (.Y(_3129_),
    .A(net2268),
    .B(net2211));
 sg13g2_nor2_2 _4108_ (.A(net2166),
    .B(net2064),
    .Y(_3130_));
 sg13g2_nor2_2 _4109_ (.A(net2127),
    .B(_2273_),
    .Y(_3131_));
 sg13g2_nand2_2 _4110_ (.Y(_3132_),
    .A(net2174),
    .B(_2262_));
 sg13g2_nor2_2 _4111_ (.A(net2123),
    .B(_1932_),
    .Y(_3133_));
 sg13g2_nand2_1 _4112_ (.Y(_3134_),
    .A(net2170),
    .B(net2085));
 sg13g2_nor2_2 _4113_ (.A(net2111),
    .B(_3124_),
    .Y(_3135_));
 sg13g2_nand2_2 _4114_ (.Y(_3136_),
    .A(net2160),
    .B(net2066));
 sg13g2_nor2_2 _4115_ (.A(net2143),
    .B(_3129_),
    .Y(_3137_));
 sg13g2_nand2_1 _4116_ (.Y(_3138_),
    .A(net2113),
    .B(net2063));
 sg13g2_nand4_1 _4117_ (.B(_3120_),
    .C(_3136_),
    .A(_3115_),
    .Y(_3139_),
    .D(_3138_));
 sg13g2_a21oi_1 _4118_ (.A1(net2443),
    .A2(_3139_),
    .Y(_3140_),
    .B1(net2493));
 sg13g2_nor2_1 _4119_ (.A(_1943_),
    .B(net2068),
    .Y(_3141_));
 sg13g2_nand3_1 _4120_ (.B(net2355),
    .C(net2069),
    .A(net2146),
    .Y(_3142_));
 sg13g2_nor2_1 _4121_ (.A(net2373),
    .B(net2362),
    .Y(_3143_));
 sg13g2_nand2_2 _4122_ (.Y(_3144_),
    .A(_1712_),
    .B(net2370));
 sg13g2_nor2_2 _4123_ (.A(net2277),
    .B(net2210),
    .Y(_3145_));
 sg13g2_nand2_2 _4124_ (.Y(_3146_),
    .A(net2261),
    .B(_3144_));
 sg13g2_nor3_2 _4125_ (.A(net2286),
    .B(net2213),
    .C(net2209),
    .Y(_3147_));
 sg13g2_nand3_1 _4126_ (.B(net2211),
    .C(_3144_),
    .A(net2262),
    .Y(_3148_));
 sg13g2_nor2_2 _4127_ (.A(net2144),
    .B(net2062),
    .Y(_3149_));
 sg13g2_nand2_2 _4128_ (.Y(_3150_),
    .A(net2095),
    .B(_3147_));
 sg13g2_nor2_2 _4129_ (.A(net2370),
    .B(net2351),
    .Y(_3151_));
 sg13g2_nand2_2 _4130_ (.Y(_3152_),
    .A(net2362),
    .B(net2353));
 sg13g2_nand2_2 _4131_ (.Y(_3153_),
    .A(net2275),
    .B(net2208));
 sg13g2_nor2_2 _4132_ (.A(net2269),
    .B(_3151_),
    .Y(_3154_));
 sg13g2_nand3_1 _4133_ (.B(_3079_),
    .C(_3152_),
    .A(net2284),
    .Y(_3155_));
 sg13g2_nand2b_1 _4134_ (.Y(_3156_),
    .B(net2120),
    .A_N(_3155_));
 sg13g2_a21o_1 _4135_ (.A2(_3155_),
    .A1(net2062),
    .B1(net2158),
    .X(_3157_));
 sg13g2_a21oi_1 _4136_ (.A1(net2062),
    .A2(_3155_),
    .Y(_3158_),
    .B1(net2142));
 sg13g2_nand3_1 _4137_ (.B(_3142_),
    .C(_3157_),
    .A(_3136_),
    .Y(_3159_));
 sg13g2_nand2_2 _4138_ (.Y(_3160_),
    .A(net2274),
    .B(net2345));
 sg13g2_nand2_2 _4139_ (.Y(_3161_),
    .A(net2360),
    .B(net2357));
 sg13g2_nor2_1 _4140_ (.A(net2370),
    .B(net2359),
    .Y(_3162_));
 sg13g2_nor2_2 _4141_ (.A(net2371),
    .B(net2347),
    .Y(_3163_));
 sg13g2_nand2_2 _4142_ (.Y(_3164_),
    .A(net2363),
    .B(net2350));
 sg13g2_nand2_1 _4143_ (.Y(_3165_),
    .A(net2283),
    .B(_3164_));
 sg13g2_nor2_2 _4144_ (.A(net2263),
    .B(_3163_),
    .Y(_3166_));
 sg13g2_nand2_2 _4145_ (.Y(_3167_),
    .A(net2118),
    .B(_3166_));
 sg13g2_o21ai_1 _4146_ (.B1(net2110),
    .Y(_3168_),
    .A1(_3147_),
    .A2(_3166_));
 sg13g2_nor2_2 _4147_ (.A(net2254),
    .B(net2353),
    .Y(_3169_));
 sg13g2_a221oi_1 _4148_ (.B2(net2061),
    .C1(net2159),
    .B1(net2062),
    .A1(net2282),
    .Y(_3170_),
    .A2(net2215));
 sg13g2_nand2_2 _4149_ (.Y(_3171_),
    .A(net2273),
    .B(net2349));
 sg13g2_nor2_2 _4150_ (.A(net2253),
    .B(_3164_),
    .Y(_3172_));
 sg13g2_nand2_2 _4151_ (.Y(_3173_),
    .A(net2363),
    .B(net2347));
 sg13g2_nor2_2 _4152_ (.A(net2366),
    .B(net2349),
    .Y(_3174_));
 sg13g2_nor2_2 _4153_ (.A(net2282),
    .B(_3173_),
    .Y(_3175_));
 sg13g2_nor2_2 _4154_ (.A(net2096),
    .B(_3175_),
    .Y(_3176_));
 sg13g2_nor2_1 _4155_ (.A(net2290),
    .B(net2220),
    .Y(_3177_));
 sg13g2_nand2_1 _4156_ (.Y(_3178_),
    .A(net2268),
    .B(_2948_));
 sg13g2_nor4_1 _4157_ (.A(net2095),
    .B(_3172_),
    .C(_3175_),
    .D(net2060),
    .Y(_3179_));
 sg13g2_or2_1 _4158_ (.X(_3180_),
    .B(_3179_),
    .A(_3170_));
 sg13g2_a221oi_1 _4159_ (.B2(net2261),
    .C1(net2112),
    .B1(_3174_),
    .A1(_3148_),
    .Y(_3181_),
    .A2(_3165_));
 sg13g2_xnor2_1 _4160_ (.Y(_3182_),
    .A(net2374),
    .B(net2372));
 sg13g2_nand2_2 _4161_ (.Y(_3183_),
    .A(net2105),
    .B(_3169_));
 sg13g2_or2_2 _4162_ (.X(_3184_),
    .B(_3182_),
    .A(net2354));
 sg13g2_nor3_1 _4163_ (.A(net2144),
    .B(net2254),
    .C(_3184_),
    .Y(_3185_));
 sg13g2_nor2_1 _4164_ (.A(_3149_),
    .B(_3185_),
    .Y(_3186_));
 sg13g2_nor3_1 _4165_ (.A(_3149_),
    .B(net2028),
    .C(_3185_),
    .Y(_3187_));
 sg13g2_nor2_1 _4166_ (.A(net2464),
    .B(_3187_),
    .Y(_3188_));
 sg13g2_a221oi_1 _4167_ (.B2(net2408),
    .C1(_3188_),
    .B1(_3180_),
    .A1(net2423),
    .Y(_3189_),
    .A2(_3159_));
 sg13g2_nand2_1 _4168_ (.Y(_3190_),
    .A(_3140_),
    .B(_3189_));
 sg13g2_nor2_1 _4169_ (.A(net2228),
    .B(_3034_),
    .Y(_3191_));
 sg13g2_nand3_1 _4170_ (.B(net2080),
    .C(net2226),
    .A(net2090),
    .Y(_3192_));
 sg13g2_nand3_1 _4171_ (.B(net2044),
    .C(_3192_),
    .A(net2485),
    .Y(_3193_));
 sg13g2_nor2_2 _4172_ (.A(net2143),
    .B(_3146_),
    .Y(_3194_));
 sg13g2_nand2_2 _4173_ (.Y(_3195_),
    .A(net2092),
    .B(_3145_));
 sg13g2_nor3_2 _4174_ (.A(net2143),
    .B(net2245),
    .C(net2061),
    .Y(_3196_));
 sg13g2_nor2_1 _4175_ (.A(_3194_),
    .B(_3196_),
    .Y(_3197_));
 sg13g2_a21oi_1 _4176_ (.A1(net2581),
    .A2(net2358),
    .Y(_3198_),
    .B1(net2028));
 sg13g2_a21oi_1 _4177_ (.A1(_3197_),
    .A2(_3198_),
    .Y(_3199_),
    .B1(net2524));
 sg13g2_nand2_2 _4178_ (.Y(_3200_),
    .A(net2062),
    .B(_3153_));
 sg13g2_nand2_1 _4179_ (.Y(_3201_),
    .A(net2163),
    .B(_3147_));
 sg13g2_nand2_1 _4180_ (.Y(_3202_),
    .A(net2154),
    .B(_3154_));
 sg13g2_nand2_1 _4181_ (.Y(_3203_),
    .A(net2143),
    .B(_3200_));
 sg13g2_nand3_1 _4182_ (.B(net2355),
    .C(_2691_),
    .A(net2122),
    .Y(_3204_));
 sg13g2_nand3_1 _4183_ (.B(_3203_),
    .C(net2025),
    .A(net2046),
    .Y(_3205_));
 sg13g2_a221oi_1 _4184_ (.B2(net2408),
    .C1(_3199_),
    .B1(_3205_),
    .A1(_1371_),
    .Y(_3206_),
    .A2(_3193_));
 sg13g2_nor2_1 _4185_ (.A(net2295),
    .B(_3206_),
    .Y(_3207_));
 sg13g2_a221oi_1 _4186_ (.B2(_3207_),
    .C1(net2376),
    .B1(_3190_),
    .A1(net2295),
    .Y(_3208_),
    .A2(_3113_));
 sg13g2_or3_2 _4187_ (.A(_3068_),
    .B(net2035),
    .C(_3208_),
    .X(_3209_));
 sg13g2_xor2_1 _4188_ (.B(net2604),
    .A(\logo_top[6] ),
    .X(_3210_));
 sg13g2_a21oi_2 _4189_ (.B1(_3071_),
    .Y(_3211_),
    .A2(net2606),
    .A1(_0702_));
 sg13g2_nor2_1 _4190_ (.A(_3210_),
    .B(_3211_),
    .Y(_3212_));
 sg13g2_xor2_1 _4191_ (.B(_3211_),
    .A(_3210_),
    .X(_3213_));
 sg13g2_xnor2_1 _4192_ (.Y(_3214_),
    .A(_3210_),
    .B(_3211_));
 sg13g2_nor2_2 _4193_ (.A(net2385),
    .B(net2499),
    .Y(_3215_));
 sg13g2_nand2_1 _4194_ (.Y(_3216_),
    .A(net2391),
    .B(net2508));
 sg13g2_nor2_2 _4195_ (.A(net2239),
    .B(_2350_),
    .Y(_3217_));
 sg13g2_nand2_1 _4196_ (.Y(_3218_),
    .A(net2237),
    .B(net2227));
 sg13g2_nand2_1 _4197_ (.Y(_3219_),
    .A(net2234),
    .B(_2844_));
 sg13g2_nor3_2 _4198_ (.A(net2286),
    .B(net2229),
    .C(_2999_),
    .Y(_3220_));
 sg13g2_nand2_2 _4199_ (.Y(_3221_),
    .A(net2367),
    .B(net2357));
 sg13g2_nor2_2 _4200_ (.A(net2364),
    .B(net2359),
    .Y(_3222_));
 sg13g2_mux2_2 _4201_ (.A0(net2358),
    .A1(net2356),
    .S(net2361),
    .X(_3223_));
 sg13g2_nand2_2 _4202_ (.Y(_3224_),
    .A(_2991_),
    .B(_3221_));
 sg13g2_nand2_1 _4203_ (.Y(_3225_),
    .A(net2256),
    .B(_3223_));
 sg13g2_nor2_2 _4204_ (.A(net2280),
    .B(_2669_),
    .Y(_3226_));
 sg13g2_nand2_2 _4205_ (.Y(_3227_),
    .A(net2256),
    .B(net2224));
 sg13g2_a22oi_1 _4206_ (.Y(_3228_),
    .B1(_3227_),
    .B2(net2041),
    .A2(_3225_),
    .A1(_3027_));
 sg13g2_nor2_1 _4207_ (.A(net2544),
    .B(_3228_),
    .Y(_3229_));
 sg13g2_nand2_1 _4208_ (.Y(_3230_),
    .A(net2278),
    .B(net2356));
 sg13g2_nor2_2 _4209_ (.A(net2266),
    .B(net2221),
    .Y(_3231_));
 sg13g2_nand2_1 _4210_ (.Y(_3232_),
    .A(net2291),
    .B(_2836_));
 sg13g2_nor2_1 _4211_ (.A(net2151),
    .B(_3231_),
    .Y(_3233_));
 sg13g2_nand2_1 _4212_ (.Y(_3234_),
    .A(net2526),
    .B(_3233_));
 sg13g2_nor2_2 _4213_ (.A(net2257),
    .B(_2669_),
    .Y(_3235_));
 sg13g2_nand2_2 _4214_ (.Y(_3236_),
    .A(net2279),
    .B(net2224));
 sg13g2_nor2_1 _4215_ (.A(net2150),
    .B(_3235_),
    .Y(_3237_));
 sg13g2_and2_2 _4216_ (.A(net2150),
    .B(_3225_),
    .X(_3238_));
 sg13g2_nand2_1 _4217_ (.Y(_3239_),
    .A(net2149),
    .B(_3225_));
 sg13g2_o21ai_1 _4218_ (.B1(net2424),
    .Y(_3240_),
    .A1(_3237_),
    .A2(_3238_));
 sg13g2_nor2_2 _4219_ (.A(net2523),
    .B(net2097),
    .Y(_3241_));
 sg13g2_o21ai_1 _4220_ (.B1(net2544),
    .Y(_3242_),
    .A1(_3056_),
    .A2(_3237_));
 sg13g2_nand3_1 _4221_ (.B(_3240_),
    .C(_3242_),
    .A(_3234_),
    .Y(_3243_));
 sg13g2_o21ai_1 _4222_ (.B1(net2203),
    .Y(_3244_),
    .A1(_3229_),
    .A2(_3243_));
 sg13g2_nand2_2 _4223_ (.Y(_3245_),
    .A(net2268),
    .B(_3163_));
 sg13g2_and2_1 _4224_ (.A(net2151),
    .B(_3245_),
    .X(_3246_));
 sg13g2_nand2_2 _4225_ (.Y(_3247_),
    .A(net2155),
    .B(_3245_));
 sg13g2_nor2_1 _4226_ (.A(net2601),
    .B(net2024),
    .Y(_3248_));
 sg13g2_nand3_1 _4227_ (.B(net2151),
    .C(_3245_),
    .A(net2564),
    .Y(_3249_));
 sg13g2_nor2_2 _4228_ (.A(net2257),
    .B(net2226),
    .Y(_3250_));
 sg13g2_nand2_1 _4229_ (.Y(_3251_),
    .A(net2278),
    .B(net2228));
 sg13g2_nor2_1 _4230_ (.A(net2578),
    .B(net2133),
    .Y(_3252_));
 sg13g2_nand2_2 _4231_ (.Y(_3253_),
    .A(net2565),
    .B(net2107));
 sg13g2_nand2_1 _4232_ (.Y(_3254_),
    .A(net2268),
    .B(_2999_));
 sg13g2_nand2_2 _4233_ (.Y(_3255_),
    .A(net2177),
    .B(_3254_));
 sg13g2_and2_2 _4234_ (.A(net2177),
    .B(_3254_),
    .X(_3256_));
 sg13g2_o21ai_1 _4235_ (.B1(_3255_),
    .Y(_3257_),
    .A1(net2154),
    .A2(_3250_));
 sg13g2_a221oi_1 _4236_ (.B2(net2103),
    .C1(_3256_),
    .B1(_3251_),
    .A1(net2564),
    .Y(_3258_),
    .A2(_3246_));
 sg13g2_nand2_1 _4237_ (.Y(_3259_),
    .A(net2093),
    .B(net2081));
 sg13g2_nor2_2 _4238_ (.A(net2270),
    .B(net2222),
    .Y(_3260_));
 sg13g2_nand2_2 _4239_ (.Y(_3261_),
    .A(net2289),
    .B(net2223));
 sg13g2_nor2_2 _4240_ (.A(net2173),
    .B(_3261_),
    .Y(_3262_));
 sg13g2_nand2_1 _4241_ (.Y(_3263_),
    .A(net2107),
    .B(_3260_));
 sg13g2_nor2_1 _4242_ (.A(net2546),
    .B(_3262_),
    .Y(_3264_));
 sg13g2_nand2_1 _4243_ (.Y(_3265_),
    .A(net2527),
    .B(net2021));
 sg13g2_nor2_2 _4244_ (.A(net2279),
    .B(net2236),
    .Y(_3266_));
 sg13g2_nand2_2 _4245_ (.Y(_3267_),
    .A(net2258),
    .B(net2238));
 sg13g2_o21ai_1 _4246_ (.B1(_3264_),
    .Y(_3268_),
    .A1(net2107),
    .A2(_3267_));
 sg13g2_nor2_2 _4247_ (.A(net2108),
    .B(_3266_),
    .Y(_3269_));
 sg13g2_nor2_1 _4248_ (.A(net2151),
    .B(_3251_),
    .Y(_3270_));
 sg13g2_nand2_2 _4249_ (.Y(_3271_),
    .A(net2107),
    .B(_3250_));
 sg13g2_mux2_2 _4250_ (.A0(_3250_),
    .A1(_3266_),
    .S(net2154),
    .X(_3272_));
 sg13g2_nand3_1 _4251_ (.B(_3268_),
    .C(_3272_),
    .A(net2488),
    .Y(_3273_));
 sg13g2_nor3_2 _4252_ (.A(net2256),
    .B(net2360),
    .C(net2345),
    .Y(_3274_));
 sg13g2_nand3_1 _4253_ (.B(net2369),
    .C(net2350),
    .A(net2278),
    .Y(_3275_));
 sg13g2_nor2_2 _4254_ (.A(net2156),
    .B(_3274_),
    .Y(_3276_));
 sg13g2_nand2_2 _4255_ (.Y(_3277_),
    .A(net2103),
    .B(_3275_));
 sg13g2_mux2_2 _4256_ (.A0(_3245_),
    .A1(_3275_),
    .S(net2103),
    .X(_3278_));
 sg13g2_o21ai_1 _4257_ (.B1(net2378),
    .Y(_3279_),
    .A1(net2330),
    .A2(_3278_));
 sg13g2_a21oi_1 _4258_ (.A1(net2339),
    .A2(_3258_),
    .Y(_3280_),
    .B1(_3279_));
 sg13g2_nor2_1 _4259_ (.A(net2378),
    .B(net2509),
    .Y(_3281_));
 sg13g2_nand2_1 _4260_ (.Y(_3282_),
    .A(net2392),
    .B(net2487));
 sg13g2_o21ai_1 _4261_ (.B1(net2151),
    .Y(_3283_),
    .A1(net2278),
    .A2(_3161_));
 sg13g2_nand2_1 _4262_ (.Y(_3284_),
    .A(_3277_),
    .B(_3283_));
 sg13g2_nor2_1 _4263_ (.A(net2107),
    .B(_3226_),
    .Y(_3285_));
 sg13g2_nand2_2 _4264_ (.Y(_3286_),
    .A(net2156),
    .B(_3227_));
 sg13g2_a21oi_1 _4265_ (.A1(_3277_),
    .A2(_3286_),
    .Y(_3287_),
    .B1(net2587));
 sg13g2_or2_1 _4266_ (.X(_3288_),
    .B(_3287_),
    .A(_3284_));
 sg13g2_nor2_2 _4267_ (.A(net2378),
    .B(net2326),
    .Y(_3289_));
 sg13g2_nand2_2 _4268_ (.Y(_3290_),
    .A(net2388),
    .B(net2328));
 sg13g2_o21ai_1 _4269_ (.B1(net2301),
    .Y(_3291_),
    .A1(net2224),
    .A2(_3290_));
 sg13g2_a221oi_1 _4270_ (.B2(_3288_),
    .C1(_3291_),
    .B1(net2195),
    .A1(_3273_),
    .Y(_3292_),
    .A2(_3280_));
 sg13g2_nor2_2 _4271_ (.A(net2092),
    .B(_2570_),
    .Y(_3293_));
 sg13g2_nor3_2 _4272_ (.A(net2103),
    .B(net2280),
    .C(net2231),
    .Y(_3294_));
 sg13g2_nand3_1 _4273_ (.B(net2257),
    .C(net2232),
    .A(net2154),
    .Y(_3295_));
 sg13g2_a21oi_2 _4274_ (.B1(net2201),
    .Y(_3296_),
    .A2(_3295_),
    .A1(net2021));
 sg13g2_nor2_2 _4275_ (.A(net2550),
    .B(net2169),
    .Y(_3297_));
 sg13g2_nand3_1 _4276_ (.B(net2253),
    .C(net2232),
    .A(net2562),
    .Y(_3298_));
 sg13g2_nand2_2 _4277_ (.Y(_3299_),
    .A(net2523),
    .B(_3298_));
 sg13g2_nor2_2 _4278_ (.A(net2299),
    .B(net2038),
    .Y(_3300_));
 sg13g2_nand2_2 _4279_ (.Y(_3301_),
    .A(net2300),
    .B(net2035));
 sg13g2_a21o_1 _4280_ (.A2(_3299_),
    .A1(_3296_),
    .B1(net2037),
    .X(_3302_));
 sg13g2_a22oi_1 _4281_ (.Y(_3303_),
    .B1(net1985),
    .B2(_3302_),
    .A2(_3292_),
    .A1(_3244_));
 sg13g2_nor2_1 _4282_ (.A(net1978),
    .B(_3303_),
    .Y(_3304_));
 sg13g2_a21oi_2 _4283_ (.B1(_3212_),
    .Y(_3305_),
    .A2(net2604),
    .A1(_0691_));
 sg13g2_xnor2_1 _4284_ (.Y(_3306_),
    .A(\logo_top[7] ),
    .B(\pix_y[7] ));
 sg13g2_nor2b_1 _4285_ (.A(_3305_),
    .B_N(_3306_),
    .Y(_3307_));
 sg13g2_xnor2_1 _4286_ (.Y(_3308_),
    .A(_3305_),
    .B(_3306_));
 sg13g2_xor2_1 _4287_ (.B(_3306_),
    .A(_3305_),
    .X(_3309_));
 sg13g2_nor2_1 _4288_ (.A(net2300),
    .B(net2037),
    .Y(_3310_));
 sg13g2_nand2_2 _4289_ (.Y(_3311_),
    .A(net2294),
    .B(net2035));
 sg13g2_nor2_2 _4290_ (.A(net2254),
    .B(_3173_),
    .Y(_3312_));
 sg13g2_nand2_2 _4291_ (.Y(_3313_),
    .A(net2283),
    .B(_3174_));
 sg13g2_nand2_2 _4292_ (.Y(_3314_),
    .A(net2128),
    .B(net2075));
 sg13g2_a21oi_1 _4293_ (.A1(net2245),
    .A2(_2912_),
    .Y(_3315_),
    .B1(net2161));
 sg13g2_and2_2 _4294_ (.A(_3313_),
    .B(_3315_),
    .X(_3316_));
 sg13g2_nand3_1 _4295_ (.B(_1855_),
    .C(_3313_),
    .A(net2115),
    .Y(_3317_));
 sg13g2_nand2_1 _4296_ (.Y(_3318_),
    .A(net2246),
    .B(net2347));
 sg13g2_nand3_1 _4297_ (.B(net2261),
    .C(_3318_),
    .A(net2159),
    .Y(_3319_));
 sg13g2_nor2_2 _4298_ (.A(net2261),
    .B(_3174_),
    .Y(_3320_));
 sg13g2_nand2_2 _4299_ (.Y(_3321_),
    .A(net2283),
    .B(_3173_));
 sg13g2_nand2_2 _4300_ (.Y(_3322_),
    .A(net2169),
    .B(_3320_));
 sg13g2_nand4_1 _4301_ (.B(_3317_),
    .C(_3319_),
    .A(net2513),
    .Y(_3323_),
    .D(_3322_));
 sg13g2_a21oi_1 _4302_ (.A1(net2592),
    .A2(_3316_),
    .Y(_3324_),
    .B1(_3323_));
 sg13g2_nor2_1 _4303_ (.A(net2335),
    .B(_3324_),
    .Y(_3325_));
 sg13g2_nand2_2 _4304_ (.Y(_3326_),
    .A(_2592_),
    .B(net2221));
 sg13g2_a221oi_1 _4305_ (.B2(net2283),
    .C1(net2116),
    .B1(_3174_),
    .A1(_2372_),
    .Y(_3327_),
    .A2(_3164_));
 sg13g2_nand2_1 _4306_ (.Y(_3328_),
    .A(net2444),
    .B(_3327_));
 sg13g2_o21ai_1 _4307_ (.B1(net2347),
    .Y(_3329_),
    .A1(net2267),
    .A2(net2363));
 sg13g2_nand3_1 _4308_ (.B(net2273),
    .C(_2592_),
    .A(net2092),
    .Y(_3330_));
 sg13g2_a221oi_1 _4309_ (.B2(_3329_),
    .C1(_2438_),
    .B1(net2040),
    .A1(_2592_),
    .Y(_3331_),
    .A2(_2647_));
 sg13g2_o21ai_1 _4310_ (.B1(_3328_),
    .Y(_3332_),
    .A1(net2531),
    .A2(_3331_));
 sg13g2_o21ai_1 _4311_ (.B1(net2110),
    .Y(_3333_),
    .A1(_3101_),
    .A2(_3163_));
 sg13g2_nand3_1 _4312_ (.B(_3322_),
    .C(_3333_),
    .A(_3319_),
    .Y(_3334_));
 sg13g2_nor3_2 _4313_ (.A(net2182),
    .B(net2270),
    .C(_3218_),
    .Y(_3335_));
 sg13g2_nor3_1 _4314_ (.A(_3135_),
    .B(_3137_),
    .C(_3335_),
    .Y(_3336_));
 sg13g2_nand2_1 _4315_ (.Y(_3337_),
    .A(_3120_),
    .B(_3336_));
 sg13g2_nor2_1 _4316_ (.A(_2691_),
    .B(_3119_),
    .Y(_3338_));
 sg13g2_mux2_1 _4317_ (.A0(_3130_),
    .A1(net2169),
    .S(_3338_),
    .X(_3339_));
 sg13g2_a21oi_2 _4318_ (.B1(net2214),
    .Y(_3340_),
    .A2(net2211),
    .A1(net2262));
 sg13g2_nor2_1 _4319_ (.A(net2167),
    .B(_3340_),
    .Y(_3341_));
 sg13g2_nor2_1 _4320_ (.A(net2284),
    .B(_3078_),
    .Y(_3342_));
 sg13g2_nand2_2 _4321_ (.Y(_3343_),
    .A(net2263),
    .B(_3079_));
 sg13g2_a21oi_1 _4322_ (.A1(_2702_),
    .A2(_3343_),
    .Y(_3344_),
    .B1(net2529));
 sg13g2_a221oi_1 _4323_ (.B2(net2040),
    .C1(net2512),
    .B1(_3344_),
    .A1(net2426),
    .Y(_3345_),
    .A2(_3341_));
 sg13g2_o21ai_1 _4324_ (.B1(_3345_),
    .Y(_3346_),
    .A1(net2405),
    .A2(_3339_));
 sg13g2_a221oi_1 _4325_ (.B2(net2477),
    .C1(_3346_),
    .B1(_3337_),
    .A1(net2444),
    .Y(_3347_),
    .A2(_3334_));
 sg13g2_o21ai_1 _4326_ (.B1(net2382),
    .Y(_3348_),
    .A1(_3325_),
    .A2(_3332_));
 sg13g2_nand2_1 _4327_ (.Y(_3349_),
    .A(net2130),
    .B(net2065));
 sg13g2_nor3_2 _4328_ (.A(net2263),
    .B(net2249),
    .C(net2239),
    .Y(_3350_));
 sg13g2_nand2_2 _4329_ (.Y(_3351_),
    .A(_1800_),
    .B(net2237));
 sg13g2_nor2_2 _4330_ (.A(net2098),
    .B(net2073),
    .Y(_3352_));
 sg13g2_a21oi_2 _4331_ (.B1(net2121),
    .Y(_3353_),
    .A2(net2072),
    .A1(net2221));
 sg13g2_nor2_2 _4332_ (.A(net2173),
    .B(_2416_),
    .Y(_3354_));
 sg13g2_nand2_1 _4333_ (.Y(_3355_),
    .A(_3018_),
    .B(net2066));
 sg13g2_a22oi_1 _4334_ (.Y(_3356_),
    .B1(_3354_),
    .B2(_3355_),
    .A2(_3353_),
    .A1(_3351_));
 sg13g2_nand2_1 _4335_ (.Y(_3357_),
    .A(net2425),
    .B(_3356_));
 sg13g2_nor2_2 _4336_ (.A(net2089),
    .B(net2429),
    .Y(_3358_));
 sg13g2_o21ai_1 _4337_ (.B1(_3358_),
    .Y(_3359_),
    .A1(net2073),
    .A2(_3350_));
 sg13g2_a21o_2 _4338_ (.A2(_3018_),
    .A1(_2647_),
    .B1(_2438_),
    .X(_3360_));
 sg13g2_o21ai_1 _4339_ (.B1(net2531),
    .Y(_3361_),
    .A1(_2438_),
    .A2(_3327_));
 sg13g2_a21oi_1 _4340_ (.A1(net2593),
    .A2(_2196_),
    .Y(_3362_),
    .B1(_3124_));
 sg13g2_a22oi_1 _4341_ (.Y(_3363_),
    .B1(_3362_),
    .B2(_3297_),
    .A2(_3360_),
    .A1(net2447));
 sg13g2_nand4_1 _4342_ (.B(_3359_),
    .C(_3361_),
    .A(_3357_),
    .Y(_3364_),
    .D(_3363_));
 sg13g2_a21oi_2 _4343_ (.B1(net2145),
    .Y(_3365_),
    .A2(net2076),
    .A1(_1811_));
 sg13g2_nor2_2 _4344_ (.A(net2128),
    .B(_1811_),
    .Y(_3366_));
 sg13g2_nand2_2 _4345_ (.Y(_3367_),
    .A(net2181),
    .B(_1800_));
 sg13g2_a21oi_2 _4346_ (.B1(net2116),
    .Y(_3368_),
    .A2(net2062),
    .A1(_1811_));
 sg13g2_nor2_2 _4347_ (.A(net2144),
    .B(net2403),
    .Y(_3369_));
 sg13g2_nand2_1 _4348_ (.Y(_3370_),
    .A(net2076),
    .B(_3153_));
 sg13g2_a22oi_1 _4349_ (.Y(_3371_),
    .B1(_3369_),
    .B2(_3370_),
    .A2(_3365_),
    .A1(net2541));
 sg13g2_a21oi_1 _4350_ (.A1(net2477),
    .A2(_3360_),
    .Y(_3372_),
    .B1(_3368_));
 sg13g2_nand2_1 _4351_ (.Y(_3373_),
    .A(_3371_),
    .B(_3372_));
 sg13g2_nor2_2 _4352_ (.A(net2299),
    .B(net2035),
    .Y(_3374_));
 sg13g2_nand2_2 _4353_ (.Y(_3375_),
    .A(net2300),
    .B(net2037));
 sg13g2_nand2_2 _4354_ (.Y(_3376_),
    .A(net2119),
    .B(net2067));
 sg13g2_nor2_2 _4355_ (.A(net2233),
    .B(net2210),
    .Y(_3377_));
 sg13g2_nand3_1 _4356_ (.B(net2291),
    .C(_3377_),
    .A(net2131),
    .Y(_3378_));
 sg13g2_nand2_2 _4357_ (.Y(_3379_),
    .A(net2151),
    .B(_2948_));
 sg13g2_nor2_2 _4358_ (.A(net2266),
    .B(net2247),
    .Y(_3380_));
 sg13g2_nand2_2 _4359_ (.Y(_3381_),
    .A(net2289),
    .B(net2248));
 sg13g2_nand3_1 _4360_ (.B(net2251),
    .C(net2247),
    .A(net2459),
    .Y(_3382_));
 sg13g2_nand2_1 _4361_ (.Y(_3383_),
    .A(net2137),
    .B(_3382_));
 sg13g2_nand3_1 _4362_ (.B(_3381_),
    .C(_3382_),
    .A(net2175),
    .Y(_3384_));
 sg13g2_nand2_2 _4363_ (.Y(_3385_),
    .A(_3379_),
    .B(_3384_));
 sg13g2_nand4_1 _4364_ (.B(_3378_),
    .C(_3379_),
    .A(_3376_),
    .Y(_3386_),
    .D(_3384_));
 sg13g2_nor2_1 _4365_ (.A(net2480),
    .B(_3386_),
    .Y(_3387_));
 sg13g2_nand2_2 _4366_ (.Y(_3388_),
    .A(net2116),
    .B(_3019_));
 sg13g2_and2_1 _4367_ (.A(_3378_),
    .B(_3388_),
    .X(_3389_));
 sg13g2_nand4_1 _4368_ (.B(_3379_),
    .C(_3384_),
    .A(_3378_),
    .Y(_3390_),
    .D(_3388_));
 sg13g2_o21ai_1 _4369_ (.B1(net2205),
    .Y(_3391_),
    .A1(net2467),
    .A2(_3390_));
 sg13g2_nor2_2 _4370_ (.A(net2172),
    .B(net2071),
    .Y(_3392_));
 sg13g2_nand2_2 _4371_ (.Y(_3393_),
    .A(net2119),
    .B(net2072));
 sg13g2_nor2_2 _4372_ (.A(_2948_),
    .B(_3393_),
    .Y(_3394_));
 sg13g2_nand3_1 _4373_ (.B(net2219),
    .C(net2072),
    .A(net2129),
    .Y(_3395_));
 sg13g2_o21ai_1 _4374_ (.B1(net2553),
    .Y(_3396_),
    .A1(_3335_),
    .A2(_3394_));
 sg13g2_nor2_2 _4375_ (.A(net2264),
    .B(net2233),
    .Y(_3397_));
 sg13g2_nand2_2 _4376_ (.Y(_3398_),
    .A(net2286),
    .B(net2230));
 sg13g2_nor2_1 _4377_ (.A(net2174),
    .B(_3398_),
    .Y(_3399_));
 sg13g2_nor3_2 _4378_ (.A(net2180),
    .B(net2229),
    .C(_3398_),
    .Y(_3400_));
 sg13g2_o21ai_1 _4379_ (.B1(net2533),
    .Y(_3401_),
    .A1(_3394_),
    .A2(_3400_));
 sg13g2_nor3_2 _4380_ (.A(net2292),
    .B(net2223),
    .C(_2999_),
    .Y(_3402_));
 sg13g2_nand2_1 _4381_ (.Y(_3403_),
    .A(net2184),
    .B(_3402_));
 sg13g2_o21ai_1 _4382_ (.B1(net2185),
    .Y(_3404_),
    .A1(_3154_),
    .A2(_3402_));
 sg13g2_a21oi_2 _4383_ (.B1(_3169_),
    .Y(_3405_),
    .A2(net2222),
    .A1(net2237));
 sg13g2_nor2_1 _4384_ (.A(net2128),
    .B(_3405_),
    .Y(_3406_));
 sg13g2_o21ai_1 _4385_ (.B1(net2497),
    .Y(_3407_),
    .A1(net2128),
    .A2(_3405_));
 sg13g2_nand2_1 _4386_ (.Y(_3408_),
    .A(_1371_),
    .B(_3407_));
 sg13g2_nand4_1 _4387_ (.B(_3401_),
    .C(_3404_),
    .A(_3396_),
    .Y(_3409_),
    .D(_3408_));
 sg13g2_nor2_2 _4388_ (.A(net2488),
    .B(net2463),
    .Y(_3410_));
 sg13g2_nand2_2 _4389_ (.Y(_3411_),
    .A(net2508),
    .B(net2475));
 sg13g2_o21ai_1 _4390_ (.B1(net2174),
    .Y(_3412_),
    .A1(net2088),
    .A2(_3219_));
 sg13g2_nor3_1 _4391_ (.A(_3335_),
    .B(_3394_),
    .C(_3411_),
    .Y(_3413_));
 sg13g2_o21ai_1 _4392_ (.B1(net2292),
    .Y(_3414_),
    .A1(net2233),
    .A2(net2209));
 sg13g2_nand2_2 _4393_ (.Y(_3415_),
    .A(net2131),
    .B(_3414_));
 sg13g2_nand3_1 _4394_ (.B(net2291),
    .C(net2221),
    .A(net2169),
    .Y(_3416_));
 sg13g2_and2_1 _4395_ (.A(_3415_),
    .B(_3416_),
    .X(_3417_));
 sg13g2_nand3_1 _4396_ (.B(_2372_),
    .C(_3164_),
    .A(net2163),
    .Y(_3418_));
 sg13g2_nor2_2 _4397_ (.A(net2487),
    .B(net2473),
    .Y(_3419_));
 sg13g2_nand2_2 _4398_ (.Y(_3420_),
    .A(net2508),
    .B(net2462));
 sg13g2_mux2_2 _4399_ (.A0(net2355),
    .A1(net2347),
    .S(net2364),
    .X(_3421_));
 sg13g2_nor2_2 _4400_ (.A(net2274),
    .B(net2429),
    .Y(_3422_));
 sg13g2_a221oi_1 _4401_ (.B2(_3422_),
    .C1(_3420_),
    .B1(_3421_),
    .A1(_3085_),
    .Y(_3423_),
    .A2(_3326_));
 sg13g2_a221oi_1 _4402_ (.B2(_3423_),
    .C1(net2397),
    .B1(_3417_),
    .A1(_3412_),
    .Y(_3424_),
    .A2(_3413_));
 sg13g2_a21oi_2 _4403_ (.B1(net2291),
    .Y(_3425_),
    .A2(net2218),
    .A1(net2460));
 sg13g2_o21ai_1 _4404_ (.B1(net2269),
    .Y(_3426_),
    .A1(net2457),
    .A2(net2216));
 sg13g2_nand2_2 _4405_ (.Y(_3427_),
    .A(net2179),
    .B(_3425_));
 sg13g2_nand2_1 _4406_ (.Y(_3428_),
    .A(_3417_),
    .B(_3427_));
 sg13g2_a22oi_1 _4407_ (.Y(_3429_),
    .B1(_3428_),
    .B2(net2198),
    .A2(_3424_),
    .A1(_3409_));
 sg13g2_o21ai_1 _4408_ (.B1(_3429_),
    .Y(_3430_),
    .A1(_3387_),
    .A2(_3391_));
 sg13g2_nor2_2 _4409_ (.A(net2300),
    .B(net2035),
    .Y(_3431_));
 sg13g2_nand2_2 _4410_ (.Y(_3432_),
    .A(net2294),
    .B(net2037));
 sg13g2_nor2_1 _4411_ (.A(net2183),
    .B(_3117_),
    .Y(_3433_));
 sg13g2_nand2_1 _4412_ (.Y(_3434_),
    .A(net2121),
    .B(_3116_));
 sg13g2_nor2_2 _4413_ (.A(_3400_),
    .B(_3433_),
    .Y(_3435_));
 sg13g2_nand2b_2 _4414_ (.Y(_3436_),
    .B(net2016),
    .A_N(_3400_));
 sg13g2_a21oi_1 _4415_ (.A1(_3404_),
    .A2(_3435_),
    .Y(_3437_),
    .B1(net2467));
 sg13g2_nor2_1 _4416_ (.A(net2437),
    .B(_3406_),
    .Y(_3438_));
 sg13g2_a21oi_1 _4417_ (.A1(net2437),
    .A2(_3404_),
    .Y(_3439_),
    .B1(_3438_));
 sg13g2_or4_1 _4418_ (.A(_3394_),
    .B(_3400_),
    .C(_3437_),
    .D(_3439_),
    .X(_3440_));
 sg13g2_nand3_1 _4419_ (.B(net2291),
    .C(_3161_),
    .A(net2184),
    .Y(_3441_));
 sg13g2_nand2_1 _4420_ (.Y(_3442_),
    .A(net2166),
    .B(_3166_));
 sg13g2_a21oi_2 _4421_ (.B1(net2129),
    .Y(_3443_),
    .A2(_3426_),
    .A1(net2061));
 sg13g2_nor2_1 _4422_ (.A(_2922_),
    .B(_3415_),
    .Y(_3444_));
 sg13g2_nor2_1 _4423_ (.A(net2311),
    .B(_3389_),
    .Y(_3445_));
 sg13g2_a21oi_1 _4424_ (.A1(_3427_),
    .A2(_3441_),
    .Y(_3446_),
    .B1(_3420_));
 sg13g2_a221oi_1 _4425_ (.B2(net2311),
    .C1(_3446_),
    .B1(_3444_),
    .A1(_3420_),
    .Y(_3447_),
    .A2(_3443_));
 sg13g2_nor2b_1 _4426_ (.A(_3445_),
    .B_N(_3447_),
    .Y(_3448_));
 sg13g2_nor2_1 _4427_ (.A(net2508),
    .B(net2431),
    .Y(_3449_));
 sg13g2_nand2_2 _4428_ (.Y(_3450_),
    .A(net2489),
    .B(net2442));
 sg13g2_nor2_2 _4429_ (.A(net2380),
    .B(net2308),
    .Y(_3451_));
 sg13g2_nand3_1 _4430_ (.B(_3404_),
    .C(_3435_),
    .A(_3314_),
    .Y(_3452_));
 sg13g2_nor2_2 _4431_ (.A(net2508),
    .B(net2416),
    .Y(_3453_));
 sg13g2_nand2_2 _4432_ (.Y(_3454_),
    .A(net2483),
    .B(net2421));
 sg13g2_nand2_1 _4433_ (.Y(_3455_),
    .A(net2397),
    .B(net2307));
 sg13g2_nand3_1 _4434_ (.B(net2271),
    .C(_3421_),
    .A(net2184),
    .Y(_3456_));
 sg13g2_and2_1 _4435_ (.A(net2027),
    .B(net2010),
    .X(_3457_));
 sg13g2_a21oi_1 _4436_ (.A1(_3389_),
    .A2(_3457_),
    .Y(_3458_),
    .B1(_3455_));
 sg13g2_nor2_2 _4437_ (.A(net2384),
    .B(net2315),
    .Y(_3459_));
 sg13g2_nand2_2 _4438_ (.Y(_3460_),
    .A(net2392),
    .B(net2318));
 sg13g2_nor2_2 _4439_ (.A(net2487),
    .B(net2431),
    .Y(_3461_));
 sg13g2_a21o_1 _4440_ (.A2(net2305),
    .A1(net2383),
    .B1(_3459_),
    .X(_3462_));
 sg13g2_a221oi_1 _4441_ (.B2(_3390_),
    .C1(_3458_),
    .B1(_3462_),
    .A1(_3451_),
    .Y(_3463_),
    .A2(_3452_));
 sg13g2_o21ai_1 _4442_ (.B1(_3463_),
    .Y(_3464_),
    .A1(net2398),
    .A2(_3448_));
 sg13g2_a21o_1 _4443_ (.A2(_3440_),
    .A1(net2205),
    .B1(_3464_),
    .X(_3465_));
 sg13g2_nor2_1 _4444_ (.A(net2553),
    .B(_2438_),
    .Y(_3466_));
 sg13g2_o21ai_1 _4445_ (.B1(net2532),
    .Y(_3467_),
    .A1(net2174),
    .A2(_2427_));
 sg13g2_a21oi_2 _4446_ (.B1(net2116),
    .Y(_3468_),
    .A2(net2068),
    .A1(_1811_));
 sg13g2_nor3_2 _4447_ (.A(net2145),
    .B(net2253),
    .C(_2836_),
    .Y(_3469_));
 sg13g2_o21ai_1 _4448_ (.B1(net2574),
    .Y(_3470_),
    .A1(_3293_),
    .A2(_3468_));
 sg13g2_or2_1 _4449_ (.X(_3471_),
    .B(_3469_),
    .A(_3368_));
 sg13g2_a221oi_1 _4450_ (.B2(net2592),
    .C1(_3467_),
    .B1(_3471_),
    .A1(net2023),
    .Y(_3472_),
    .A2(_3320_));
 sg13g2_nor3_2 _4451_ (.A(net2130),
    .B(net2291),
    .C(_3218_),
    .Y(_3473_));
 sg13g2_and2_1 _4452_ (.A(net2374),
    .B(_3335_),
    .X(_3474_));
 sg13g2_nor3_2 _4453_ (.A(_3366_),
    .B(_3473_),
    .C(_3474_),
    .Y(_3475_));
 sg13g2_o21ai_1 _4454_ (.B1(net2553),
    .Y(_3476_),
    .A1(net2174),
    .A2(_2427_));
 sg13g2_xnor2_1 _4455_ (.Y(_3477_),
    .A(net2136),
    .B(net2273));
 sg13g2_mux2_2 _4456_ (.A0(_3227_),
    .A1(_3236_),
    .S(net2102),
    .X(_3478_));
 sg13g2_nor2_2 _4457_ (.A(net2563),
    .B(_3478_),
    .Y(_3479_));
 sg13g2_nor2_1 _4458_ (.A(_3476_),
    .B(_3479_),
    .Y(_3480_));
 sg13g2_a22oi_1 _4459_ (.Y(_3481_),
    .B1(_3475_),
    .B2(_3480_),
    .A2(_3472_),
    .A1(_3470_));
 sg13g2_o21ai_1 _4460_ (.B1(net2511),
    .Y(_3482_),
    .A1(net2403),
    .A2(_3257_));
 sg13g2_a21oi_1 _4461_ (.A1(_3217_),
    .A2(net2023),
    .Y(_3483_),
    .B1(_3476_));
 sg13g2_o21ai_1 _4462_ (.B1(net2181),
    .Y(_3484_),
    .A1(net2088),
    .A2(_3402_));
 sg13g2_nand2_2 _4463_ (.Y(_3485_),
    .A(_3367_),
    .B(_3403_));
 sg13g2_nand3b_1 _4464_ (.B(_3483_),
    .C(_3484_),
    .Y(_3486_),
    .A_N(_3474_));
 sg13g2_a21oi_1 _4465_ (.A1(_3466_),
    .A2(_3475_),
    .Y(_3487_),
    .B1(_3482_));
 sg13g2_a221oi_1 _4466_ (.B2(_3487_),
    .C1(net2398),
    .B1(_3486_),
    .A1(net2497),
    .Y(_3488_),
    .A2(_3481_));
 sg13g2_o21ai_1 _4467_ (.B1(net2127),
    .Y(_3489_),
    .A1(_2416_),
    .A2(net2055));
 sg13g2_nor3_1 _4468_ (.A(net2419),
    .B(_2797_),
    .C(_3400_),
    .Y(_3490_));
 sg13g2_a21oi_1 _4469_ (.A1(net2419),
    .A2(_3489_),
    .Y(_3491_),
    .B1(_3490_));
 sg13g2_nor3_1 _4470_ (.A(net2192),
    .B(_3485_),
    .C(_3491_),
    .Y(_3492_));
 sg13g2_nor3_2 _4471_ (.A(net2264),
    .B(net2225),
    .C(_2982_),
    .Y(_3493_));
 sg13g2_nor2_1 _4472_ (.A(_2941_),
    .B(_3493_),
    .Y(_3494_));
 sg13g2_a21oi_1 _4473_ (.A1(net2575),
    .A2(_2559_),
    .Y(_3495_),
    .B1(_3494_));
 sg13g2_nand4_1 _4474_ (.B(_3441_),
    .C(net2010),
    .A(net2534),
    .Y(_3496_),
    .D(_3495_));
 sg13g2_or3_1 _4475_ (.A(net2534),
    .B(_3443_),
    .C(_3444_),
    .X(_3497_));
 sg13g2_a21oi_1 _4476_ (.A1(_3496_),
    .A2(_3497_),
    .Y(_3498_),
    .B1(net2201));
 sg13g2_nor4_2 _4477_ (.A(net2039),
    .B(_3488_),
    .C(_3492_),
    .Y(_3499_),
    .D(_3498_));
 sg13g2_a221oi_1 _4478_ (.B2(net2207),
    .C1(net2302),
    .B1(_3373_),
    .A1(net2197),
    .Y(_3500_),
    .A2(_3364_));
 sg13g2_o21ai_1 _4479_ (.B1(_3500_),
    .Y(_3501_),
    .A1(_3347_),
    .A2(_3348_));
 sg13g2_o21ai_1 _4480_ (.B1(_3501_),
    .Y(_3502_),
    .A1(_3310_),
    .A2(_3499_));
 sg13g2_a221oi_1 _4481_ (.B2(_3465_),
    .C1(_3214_),
    .B1(_3431_),
    .A1(_3374_),
    .Y(_3503_),
    .A2(_3430_));
 sg13g2_a221oi_1 _4482_ (.B2(_3503_),
    .C1(_3308_),
    .B1(_3502_),
    .A1(_3209_),
    .Y(_3504_),
    .A2(_3304_));
 sg13g2_xnor2_1 _4483_ (.Y(_3505_),
    .A(\logo_left[0] ),
    .B(\pix_x[0] ));
 sg13g2_xor2_1 _4484_ (.B(\pix_x[0] ),
    .A(\logo_left[0] ),
    .X(_3506_));
 sg13g2_a22oi_1 _4485_ (.Y(_3507_),
    .B1(_3360_),
    .B2(_3236_),
    .A2(_3313_),
    .A1(net2045));
 sg13g2_nor2_1 _4486_ (.A(net2466),
    .B(_3507_),
    .Y(_3508_));
 sg13g2_nand2_2 _4487_ (.Y(_3509_),
    .A(net2175),
    .B(net2243));
 sg13g2_o21ai_1 _4488_ (.B1(net2351),
    .Y(_3510_),
    .A1(net2374),
    .A2(net2363));
 sg13g2_a21oi_2 _4489_ (.B1(net2354),
    .Y(_3511_),
    .A2(net2372),
    .A1(net2375));
 sg13g2_nor2_2 _4490_ (.A(net2290),
    .B(_3511_),
    .Y(_3512_));
 sg13g2_nand2_2 _4491_ (.Y(_3513_),
    .A(net2261),
    .B(_3510_));
 sg13g2_nor2_2 _4492_ (.A(net2097),
    .B(_3513_),
    .Y(_3514_));
 sg13g2_a21oi_1 _4493_ (.A1(_3321_),
    .A2(_3513_),
    .Y(_3515_),
    .B1(net2111));
 sg13g2_nand2_1 _4494_ (.Y(_3516_),
    .A(net2447),
    .B(_3515_));
 sg13g2_nor3_2 _4495_ (.A(net2258),
    .B(_2581_),
    .C(_2836_),
    .Y(_3517_));
 sg13g2_nand3_1 _4496_ (.B(_2592_),
    .C(net2221),
    .A(net2283),
    .Y(_3518_));
 sg13g2_a21oi_1 _4497_ (.A1(net2076),
    .A2(_3518_),
    .Y(_3519_),
    .B1(net2161));
 sg13g2_a22oi_1 _4498_ (.Y(_3520_),
    .B1(_3519_),
    .B2(net2343),
    .A2(_3327_),
    .A1(net2411));
 sg13g2_nor2_1 _4499_ (.A(net2435),
    .B(_3317_),
    .Y(_3521_));
 sg13g2_nor2_1 _4500_ (.A(net2513),
    .B(_3521_),
    .Y(_3522_));
 sg13g2_nand3_1 _4501_ (.B(_3152_),
    .C(_3321_),
    .A(_3144_),
    .Y(_3523_));
 sg13g2_nand3_1 _4502_ (.B(net2427),
    .C(_3523_),
    .A(net2159),
    .Y(_3524_));
 sg13g2_nand4_1 _4503_ (.B(_3520_),
    .C(_3522_),
    .A(_3516_),
    .Y(_3525_),
    .D(_3524_));
 sg13g2_nor2_2 _4504_ (.A(net2093),
    .B(_3021_),
    .Y(_3526_));
 sg13g2_nand2_1 _4505_ (.Y(_3527_),
    .A(net2592),
    .B(_3526_));
 sg13g2_nand2_2 _4506_ (.Y(_3528_),
    .A(net2257),
    .B(net2217));
 sg13g2_nand3_1 _4507_ (.B(net2077),
    .C(net2217),
    .A(net2137),
    .Y(_3529_));
 sg13g2_nor2_1 _4508_ (.A(net2592),
    .B(_3529_),
    .Y(_3530_));
 sg13g2_a221oi_1 _4509_ (.B2(net2245),
    .C1(net2161),
    .B1(_2912_),
    .A1(net2288),
    .Y(_3531_),
    .A2(net2238));
 sg13g2_o21ai_1 _4510_ (.B1(net2335),
    .Y(_3532_),
    .A1(net2111),
    .A2(_2702_));
 sg13g2_nor3_1 _4511_ (.A(_3530_),
    .B(_3531_),
    .C(_3532_),
    .Y(_3533_));
 sg13g2_nor3_1 _4512_ (.A(_2537_),
    .B(_3316_),
    .C(_3514_),
    .Y(_3534_));
 sg13g2_a221oi_1 _4513_ (.B2(_3322_),
    .C1(net2395),
    .B1(_3534_),
    .A1(_3527_),
    .Y(_3535_),
    .A2(_3533_));
 sg13g2_o21ai_1 _4514_ (.B1(_3535_),
    .Y(_3536_),
    .A1(_3508_),
    .A2(_3525_));
 sg13g2_nor2_2 _4515_ (.A(_3170_),
    .B(net2028),
    .Y(_3537_));
 sg13g2_o21ai_1 _4516_ (.B1(net2476),
    .Y(_3538_),
    .A1(_3170_),
    .A2(net2028));
 sg13g2_a21oi_1 _4517_ (.A1(net2283),
    .A2(net2246),
    .Y(_3539_),
    .B1(net2347));
 sg13g2_and2_1 _4518_ (.A(_3267_),
    .B(_3539_),
    .X(_3540_));
 sg13g2_a21oi_2 _4519_ (.B1(net2110),
    .Y(_3541_),
    .A2(_3539_),
    .A1(_3267_));
 sg13g2_nand3_1 _4520_ (.B(net2243),
    .C(net2355),
    .A(net2279),
    .Y(_3542_));
 sg13g2_nor2_1 _4521_ (.A(net2153),
    .B(_3542_),
    .Y(_3543_));
 sg13g2_a21oi_2 _4522_ (.B1(net2140),
    .Y(_3544_),
    .A2(_3542_),
    .A1(_2383_));
 sg13g2_o21ai_1 _4523_ (.B1(net2443),
    .Y(_3545_),
    .A1(_3541_),
    .A2(_3544_));
 sg13g2_nand2_2 _4524_ (.Y(_3546_),
    .A(net2120),
    .B(net2085));
 sg13g2_a21oi_1 _4525_ (.A1(net2083),
    .A2(_2383_),
    .Y(_3547_),
    .B1(net2158));
 sg13g2_nor2_1 _4526_ (.A(net2358),
    .B(net2238),
    .Y(_3548_));
 sg13g2_nor3_2 _4527_ (.A(net2375),
    .B(net2224),
    .C(net2212),
    .Y(_3549_));
 sg13g2_nand3_1 _4528_ (.B(_3079_),
    .C(_3166_),
    .A(net2110),
    .Y(_3550_));
 sg13g2_nand3_1 _4529_ (.B(net2242),
    .C(_3147_),
    .A(net2158),
    .Y(_3551_));
 sg13g2_nand4_1 _4530_ (.B(net2011),
    .C(_3550_),
    .A(net2048),
    .Y(_3552_),
    .D(_3551_));
 sg13g2_nand3_1 _4531_ (.B(net2086),
    .C(net2237),
    .A(net2130),
    .Y(_3553_));
 sg13g2_nand4_1 _4532_ (.B(_1921_),
    .C(net2237),
    .A(net2111),
    .Y(_3554_),
    .D(_3318_));
 sg13g2_nand4_1 _4533_ (.B(net2011),
    .C(_3551_),
    .A(net2048),
    .Y(_3555_),
    .D(_3554_));
 sg13g2_a22oi_1 _4534_ (.Y(_3556_),
    .B1(_3555_),
    .B2(net2425),
    .A2(_3552_),
    .A1(net2410));
 sg13g2_nand3_1 _4535_ (.B(_3545_),
    .C(_3556_),
    .A(_3538_),
    .Y(_3557_));
 sg13g2_nand2_1 _4536_ (.Y(_3558_),
    .A(net2207),
    .B(_3557_));
 sg13g2_nand2_1 _4537_ (.Y(_3559_),
    .A(net2588),
    .B(net2361));
 sg13g2_nand2_2 _4538_ (.Y(_3560_),
    .A(net2593),
    .B(_2836_));
 sg13g2_nand3_1 _4539_ (.B(_3529_),
    .C(_3560_),
    .A(_3136_),
    .Y(_3561_));
 sg13g2_o21ai_1 _4540_ (.B1(_3459_),
    .Y(_3562_),
    .A1(_3531_),
    .A2(_3561_));
 sg13g2_nand2_1 _4541_ (.Y(_3563_),
    .A(_3200_),
    .B(_3315_));
 sg13g2_nor3_2 _4542_ (.A(net2273),
    .B(net2356),
    .C(net2228),
    .Y(_3564_));
 sg13g2_nand3_1 _4543_ (.B(net2355),
    .C(net2226),
    .A(net2252),
    .Y(_3565_));
 sg13g2_o21ai_1 _4544_ (.B1(net2158),
    .Y(_3566_),
    .A1(net2065),
    .A2(_3564_));
 sg13g2_a21oi_1 _4545_ (.A1(_3124_),
    .A2(_3565_),
    .Y(_3567_),
    .B1(net2122));
 sg13g2_nand3_1 _4546_ (.B(_3563_),
    .C(_3566_),
    .A(net2593),
    .Y(_3568_));
 sg13g2_nand2_1 _4547_ (.Y(_3569_),
    .A(_3085_),
    .B(_3184_));
 sg13g2_and3_1 _4548_ (.X(_3570_),
    .A(net2570),
    .B(net2012),
    .C(_3569_));
 sg13g2_a21oi_1 _4549_ (.A1(_3186_),
    .A2(_3570_),
    .Y(_3571_),
    .B1(_3290_));
 sg13g2_a21oi_1 _4550_ (.A1(_3568_),
    .A2(_3571_),
    .Y(_3572_),
    .B1(net2302));
 sg13g2_nand4_1 _4551_ (.B(_3558_),
    .C(_3562_),
    .A(_3536_),
    .Y(_3573_),
    .D(_3572_));
 sg13g2_nor2_2 _4552_ (.A(net2135),
    .B(_3171_),
    .Y(_3574_));
 sg13g2_nand2b_2 _4553_ (.Y(_3575_),
    .B(net2093),
    .A_N(_3171_));
 sg13g2_nor2_1 _4554_ (.A(net2249),
    .B(_2826_),
    .Y(_3576_));
 sg13g2_nand3_1 _4555_ (.B(net2246),
    .C(_2816_),
    .A(net2112),
    .Y(_3577_));
 sg13g2_nor3_2 _4556_ (.A(net2135),
    .B(net2249),
    .C(_3171_),
    .Y(_3578_));
 sg13g2_nor3_2 _4557_ (.A(net2520),
    .B(_3095_),
    .C(net2009),
    .Y(_3579_));
 sg13g2_nor2_2 _4558_ (.A(net2484),
    .B(_3579_),
    .Y(_3580_));
 sg13g2_nand2_1 _4559_ (.Y(_3581_),
    .A(net2042),
    .B(_3330_));
 sg13g2_nand3_1 _4560_ (.B(_3330_),
    .C(_3383_),
    .A(net2042),
    .Y(_3582_));
 sg13g2_nor2_1 _4561_ (.A(net2346),
    .B(net2079),
    .Y(_3583_));
 sg13g2_o21ai_1 _4562_ (.B1(_3383_),
    .Y(_3584_),
    .A1(_2941_),
    .A2(_3583_));
 sg13g2_a221oi_1 _4563_ (.B2(net2407),
    .C1(_3089_),
    .B1(_3584_),
    .A1(net2471),
    .Y(_3585_),
    .A2(_3582_));
 sg13g2_nand2_2 _4564_ (.Y(_3586_),
    .A(net2127),
    .B(_2559_));
 sg13g2_a21oi_2 _4565_ (.B1(net2137),
    .Y(_3587_),
    .A2(_2570_),
    .A1(_1866_));
 sg13g2_or3_1 _4566_ (.A(net2503),
    .B(_2086_),
    .C(_3587_),
    .X(_3588_));
 sg13g2_a22oi_1 _4567_ (.Y(_3589_),
    .B1(_3588_),
    .B2(net2325),
    .A2(_3382_),
    .A1(_3358_));
 sg13g2_nand3_1 _4568_ (.B(net2240),
    .C(net2226),
    .A(net2133),
    .Y(_3590_));
 sg13g2_o21ai_1 _4569_ (.B1(_3590_),
    .Y(_3591_),
    .A1(net2089),
    .A2(net2250));
 sg13g2_a22oi_1 _4570_ (.Y(_3592_),
    .B1(_3591_),
    .B2(net2422),
    .A2(_3581_),
    .A1(net2539));
 sg13g2_a221oi_1 _4571_ (.B2(_3592_),
    .C1(net2376),
    .B1(_3589_),
    .A1(_3580_),
    .Y(_3593_),
    .A2(_3585_));
 sg13g2_nor2_2 _4572_ (.A(net2095),
    .B(net2079),
    .Y(_3594_));
 sg13g2_nand2_2 _4573_ (.Y(_3595_),
    .A(net2146),
    .B(_2075_));
 sg13g2_nand3_1 _4574_ (.B(net2242),
    .C(net2063),
    .A(net2158),
    .Y(_3596_));
 sg13g2_and3_1 _4575_ (.X(_3597_),
    .A(net2583),
    .B(_3595_),
    .C(_3596_));
 sg13g2_nor2_1 _4576_ (.A(net2314),
    .B(_3544_),
    .Y(_3598_));
 sg13g2_o21ai_1 _4577_ (.B1(_3598_),
    .Y(_3599_),
    .A1(_2892_),
    .A2(_3597_));
 sg13g2_nand4_1 _4578_ (.B(net2141),
    .C(net2231),
    .A(net2578),
    .Y(_3600_),
    .D(_2570_));
 sg13g2_and2_1 _4579_ (.A(net2090),
    .B(_3160_),
    .X(_3601_));
 sg13g2_nor3_1 _4580_ (.A(_2328_),
    .B(net2330),
    .C(_3601_),
    .Y(_3602_));
 sg13g2_a21oi_1 _4581_ (.A1(net2338),
    .A2(_3600_),
    .Y(_3603_),
    .B1(_3602_));
 sg13g2_nor3_2 _4582_ (.A(net2251),
    .B(net2349),
    .C(net2228),
    .Y(_3604_));
 sg13g2_nor2_1 _4583_ (.A(net2140),
    .B(_3604_),
    .Y(_3605_));
 sg13g2_nor2_2 _4584_ (.A(net2461),
    .B(net2134),
    .Y(_3606_));
 sg13g2_nand2_2 _4585_ (.Y(_3607_),
    .A(net2470),
    .B(net2089));
 sg13g2_o21ai_1 _4586_ (.B1(net2407),
    .Y(_3608_),
    .A1(_2086_),
    .A2(_3601_));
 sg13g2_o21ai_1 _4587_ (.B1(_3608_),
    .Y(_3609_),
    .A1(_3604_),
    .A2(_3607_));
 sg13g2_nor3_2 _4588_ (.A(net2096),
    .B(net2238),
    .C(_2559_),
    .Y(_3610_));
 sg13g2_a21oi_1 _4589_ (.A1(net2561),
    .A2(net2075),
    .Y(_3611_),
    .B1(_3610_));
 sg13g2_nand2_2 _4590_ (.Y(_3612_),
    .A(net2240),
    .B(_2713_));
 sg13g2_nand4_1 _4591_ (.B(net2329),
    .C(_3611_),
    .A(net2046),
    .Y(_3613_),
    .D(_3612_));
 sg13g2_o21ai_1 _4592_ (.B1(_3613_),
    .Y(_3614_),
    .A1(_3603_),
    .A2(_3609_));
 sg13g2_nand3b_1 _4593_ (.B(_3599_),
    .C(net2376),
    .Y(_3615_),
    .A_N(_3614_));
 sg13g2_nand3b_1 _4594_ (.B(_3615_),
    .C(net2301),
    .Y(_3616_),
    .A_N(_3593_));
 sg13g2_nand3_1 _4595_ (.B(_3573_),
    .C(_3616_),
    .A(net2038),
    .Y(_3617_));
 sg13g2_nor2_2 _4596_ (.A(net2223),
    .B(_3153_),
    .Y(_3618_));
 sg13g2_nand2_1 _4597_ (.Y(_3619_),
    .A(net2222),
    .B(_3154_));
 sg13g2_nand2_1 _4598_ (.Y(_3620_),
    .A(net2099),
    .B(_3618_));
 sg13g2_a21oi_2 _4599_ (.B1(net2180),
    .Y(_3621_),
    .A2(_3619_),
    .A1(net2076));
 sg13g2_nor3_1 _4600_ (.A(_3293_),
    .B(_3468_),
    .C(_3621_),
    .Y(_3622_));
 sg13g2_nor2_1 _4601_ (.A(net2532),
    .B(_3622_),
    .Y(_3623_));
 sg13g2_a22oi_1 _4602_ (.Y(_3624_),
    .B1(_3269_),
    .B2(_3381_),
    .A2(net2222),
    .A1(net2126));
 sg13g2_o21ai_1 _4603_ (.B1(net2480),
    .Y(_3625_),
    .A1(net2088),
    .A2(_2787_));
 sg13g2_o21ai_1 _4604_ (.B1(_3625_),
    .Y(_3626_),
    .A1(net2553),
    .A2(_3624_));
 sg13g2_nor3_1 _4605_ (.A(net2518),
    .B(_3623_),
    .C(_3626_),
    .Y(_3627_));
 sg13g2_o21ai_1 _4606_ (.B1(net2436),
    .Y(_3628_),
    .A1(_3366_),
    .A2(_3621_));
 sg13g2_o21ai_1 _4607_ (.B1(net2117),
    .Y(_3629_),
    .A1(_2416_),
    .A2(_3166_));
 sg13g2_a21oi_1 _4608_ (.A1(net2076),
    .A2(net2061),
    .Y(_3630_),
    .B1(net2180));
 sg13g2_nand2_2 _4609_ (.Y(_3631_),
    .A(net2180),
    .B(_2931_));
 sg13g2_nor2_1 _4610_ (.A(_3380_),
    .B(_3631_),
    .Y(_3632_));
 sg13g2_o21ai_1 _4611_ (.B1(net2448),
    .Y(_0086_),
    .A1(_3630_),
    .A2(_3632_));
 sg13g2_nand3_1 _4612_ (.B(net2169),
    .C(_3147_),
    .A(net2530),
    .Y(_0087_));
 sg13g2_nand3_1 _4613_ (.B(net2230),
    .C(net2064),
    .A(net2171),
    .Y(_0088_));
 sg13g2_or2_1 _4614_ (.X(_0089_),
    .B(_0088_),
    .A(net2420));
 sg13g2_nand4_1 _4615_ (.B(_0086_),
    .C(_0087_),
    .A(_3628_),
    .Y(_0090_),
    .D(_0089_));
 sg13g2_o21ai_1 _4616_ (.B1(net2385),
    .Y(_0091_),
    .A1(net2498),
    .A2(_0090_));
 sg13g2_a21oi_1 _4617_ (.A1(_3236_),
    .A2(_3360_),
    .Y(_0092_),
    .B1(net2531));
 sg13g2_nand3_1 _4618_ (.B(net2268),
    .C(_3224_),
    .A(net2173),
    .Y(_0093_));
 sg13g2_nand2_2 _4619_ (.Y(_0094_),
    .A(net2171),
    .B(_3350_));
 sg13g2_a21oi_1 _4620_ (.A1(_0093_),
    .A2(_0094_),
    .Y(_0095_),
    .B1(net2574));
 sg13g2_nand3_1 _4621_ (.B(_2625_),
    .C(_3313_),
    .A(net2574),
    .Y(_0096_));
 sg13g2_nand3b_1 _4622_ (.B(_0096_),
    .C(_0092_),
    .Y(_0097_),
    .A_N(_0095_));
 sg13g2_nand3_1 _4623_ (.B(net2263),
    .C(_3011_),
    .A(net2167),
    .Y(_0098_));
 sg13g2_nand2_1 _4624_ (.Y(_0099_),
    .A(_0094_),
    .B(_0098_));
 sg13g2_o21ai_1 _4625_ (.B1(net2351),
    .Y(_0100_),
    .A1(net2460),
    .A2(net2370));
 sg13g2_nor2_2 _4626_ (.A(net2353),
    .B(net2239),
    .Y(_0101_));
 sg13g2_nand2_2 _4627_ (.Y(_0102_),
    .A(net2265),
    .B(_0100_));
 sg13g2_a21oi_1 _4628_ (.A1(net2248),
    .A2(_2570_),
    .Y(_0103_),
    .B1(net2060));
 sg13g2_a221oi_1 _4629_ (.B2(net2040),
    .C1(_3467_),
    .B1(_0103_),
    .A1(net2570),
    .Y(_0104_),
    .A2(_0099_));
 sg13g2_a21oi_1 _4630_ (.A1(_2724_),
    .A2(_0104_),
    .Y(_0105_),
    .B1(net2201));
 sg13g2_nor4_1 _4631_ (.A(net2435),
    .B(_2438_),
    .C(_2713_),
    .D(_3468_),
    .Y(_0106_));
 sg13g2_o21ai_1 _4632_ (.B1(net2163),
    .Y(_0107_),
    .A1(net2088),
    .A2(net2067));
 sg13g2_nand3_1 _4633_ (.B(_3629_),
    .C(_0107_),
    .A(net2435),
    .Y(_0108_));
 sg13g2_nor2_1 _4634_ (.A(net2192),
    .B(_0106_),
    .Y(_0109_));
 sg13g2_nand2_2 _4635_ (.Y(_0110_),
    .A(net2472),
    .B(net2196));
 sg13g2_o21ai_1 _4636_ (.B1(net2302),
    .Y(_0111_),
    .A1(net2357),
    .A2(_0110_));
 sg13g2_a221oi_1 _4637_ (.B2(_0109_),
    .C1(_0111_),
    .B1(_0108_),
    .A1(_0097_),
    .Y(_0112_),
    .A2(_0105_));
 sg13g2_o21ai_1 _4638_ (.B1(_0112_),
    .Y(_0113_),
    .A1(_3627_),
    .A2(_0091_));
 sg13g2_nor2_2 _4639_ (.A(_3266_),
    .B(_3384_),
    .Y(_0114_));
 sg13g2_nand4_1 _4640_ (.B(_3267_),
    .C(_3381_),
    .A(net2175),
    .Y(_0115_),
    .D(_3382_));
 sg13g2_nor4_1 _4641_ (.A(net2404),
    .B(_2797_),
    .C(_3400_),
    .D(_0114_),
    .Y(_0116_));
 sg13g2_nor3_1 _4642_ (.A(net2467),
    .B(_2394_),
    .C(_3399_),
    .Y(_0117_));
 sg13g2_a221oi_1 _4643_ (.B2(_2936_),
    .C1(net2532),
    .B1(_2317_),
    .A1(net2574),
    .Y(_0118_),
    .A2(net2452));
 sg13g2_o21ai_1 _4644_ (.B1(_3118_),
    .Y(_0119_),
    .A1(_0117_),
    .A2(_0118_));
 sg13g2_o21ai_1 _4645_ (.B1(net2205),
    .Y(_0120_),
    .A1(_3366_),
    .A2(_0119_));
 sg13g2_or2_1 _4646_ (.X(_0121_),
    .B(_0120_),
    .A(_0116_));
 sg13g2_a21o_1 _4647_ (.A2(net2305),
    .A1(net2383),
    .B1(net2198),
    .X(_0122_));
 sg13g2_nand4_1 _4648_ (.B(_3378_),
    .C(_3379_),
    .A(net2049),
    .Y(_0123_),
    .D(_3384_));
 sg13g2_nor2_2 _4649_ (.A(net2392),
    .B(net2488),
    .Y(_0124_));
 sg13g2_nand3_1 _4650_ (.B(_3390_),
    .C(_0124_),
    .A(net2414),
    .Y(_0125_));
 sg13g2_nand2_1 _4651_ (.Y(_0126_),
    .A(net2296),
    .B(_0125_));
 sg13g2_a221oi_1 _4652_ (.B2(_0123_),
    .C1(_0126_),
    .B1(_0122_),
    .A1(net2383),
    .Y(_0127_),
    .A2(_3386_));
 sg13g2_a21oi_1 _4653_ (.A1(_0121_),
    .A2(_0127_),
    .Y(_0128_),
    .B1(_3072_));
 sg13g2_a21oi_1 _4654_ (.A1(_0113_),
    .A2(_0128_),
    .Y(_0129_),
    .B1(net1980));
 sg13g2_nor3_2 _4655_ (.A(net2161),
    .B(_1811_),
    .C(net2209),
    .Y(_0130_));
 sg13g2_nor3_1 _4656_ (.A(_2394_),
    .B(_3135_),
    .C(_0130_),
    .Y(_0131_));
 sg13g2_nand3_1 _4657_ (.B(net2266),
    .C(net2221),
    .A(net2169),
    .Y(_0132_));
 sg13g2_nand3_1 _4658_ (.B(net2221),
    .C(net2063),
    .A(net2162),
    .Y(_0133_));
 sg13g2_and2_1 _4659_ (.A(_0131_),
    .B(_0133_),
    .X(_0134_));
 sg13g2_o21ai_1 _4660_ (.B1(net2562),
    .Y(_0135_),
    .A1(_2797_),
    .A2(_0130_));
 sg13g2_nand3_1 _4661_ (.B(_0134_),
    .C(_0135_),
    .A(net2523),
    .Y(_0136_));
 sg13g2_nor2_1 _4662_ (.A(_3007_),
    .B(_3183_),
    .Y(_0137_));
 sg13g2_mux2_2 _4663_ (.A0(_1899_),
    .A1(net2213),
    .S(net2266),
    .X(_0138_));
 sg13g2_nor3_2 _4664_ (.A(net2457),
    .B(net2286),
    .C(net2246),
    .Y(_0139_));
 sg13g2_nor2_2 _4665_ (.A(net2123),
    .B(_0139_),
    .Y(_0140_));
 sg13g2_or3_2 _4666_ (.A(net2124),
    .B(_0138_),
    .C(_0139_),
    .X(_0141_));
 sg13g2_a21oi_1 _4667_ (.A1(net2569),
    .A2(net2359),
    .Y(_0142_),
    .B1(_0137_));
 sg13g2_nand4_1 _4668_ (.B(net2043),
    .C(_0141_),
    .A(net2548),
    .Y(_0143_),
    .D(_0142_));
 sg13g2_a21oi_1 _4669_ (.A1(_0136_),
    .A2(_0143_),
    .Y(_0144_),
    .B1(net2504));
 sg13g2_a21oi_1 _4670_ (.A1(net2275),
    .A2(_3076_),
    .Y(_0145_),
    .B1(_3091_));
 sg13g2_nor2_1 _4671_ (.A(net2065),
    .B(net2063),
    .Y(_0146_));
 sg13g2_a22oi_1 _4672_ (.Y(_0147_),
    .B1(_0146_),
    .B2(net2041),
    .A2(_0145_),
    .A1(_2778_));
 sg13g2_o21ai_1 _4673_ (.B1(net2390),
    .Y(_0148_),
    .A1(net2336),
    .A2(_0147_));
 sg13g2_nand2_2 _4674_ (.Y(_0149_),
    .A(net2552),
    .B(net2116));
 sg13g2_nor4_2 _4675_ (.A(net2523),
    .B(net2145),
    .C(net2252),
    .Y(_0150_),
    .D(net2235));
 sg13g2_nand2_1 _4676_ (.Y(_0151_),
    .A(net2241),
    .B(_0150_));
 sg13g2_a21oi_2 _4677_ (.B1(net2589),
    .Y(_0152_),
    .A2(_3250_),
    .A1(net2107));
 sg13g2_nor2_2 _4678_ (.A(net2546),
    .B(_0152_),
    .Y(_0153_));
 sg13g2_nand2_2 _4679_ (.Y(_0154_),
    .A(net2236),
    .B(net2218));
 sg13g2_nand3_1 _4680_ (.B(net2236),
    .C(net2217),
    .A(net2252),
    .Y(_0155_));
 sg13g2_inv_1 _4681_ (.Y(_0156_),
    .A(_0155_));
 sg13g2_nor2_2 _4682_ (.A(net2265),
    .B(net2208),
    .Y(_0157_));
 sg13g2_nand2_1 _4683_ (.Y(_0158_),
    .A(net2291),
    .B(_3151_));
 sg13g2_nor2_2 _4684_ (.A(net2099),
    .B(_0157_),
    .Y(_0159_));
 sg13g2_a221oi_1 _4685_ (.B2(_0159_),
    .C1(net2486),
    .B1(_0155_),
    .A1(net2441),
    .Y(_0160_),
    .A2(net2232));
 sg13g2_nand3_1 _4686_ (.B(_0151_),
    .C(_0160_),
    .A(net2049),
    .Y(_0161_));
 sg13g2_nor2_1 _4687_ (.A(_0153_),
    .B(_0161_),
    .Y(_0162_));
 sg13g2_nor3_1 _4688_ (.A(_0144_),
    .B(_0148_),
    .C(_0162_),
    .Y(_0163_));
 sg13g2_nor3_1 _4689_ (.A(net2095),
    .B(_2603_),
    .C(_3172_),
    .Y(_0164_));
 sg13g2_nor2_2 _4690_ (.A(net2263),
    .B(_3122_),
    .Y(_0165_));
 sg13g2_nand2_2 _4691_ (.Y(_0166_),
    .A(net2279),
    .B(net2214));
 sg13g2_nor2_2 _4692_ (.A(net2252),
    .B(net2234),
    .Y(_0167_));
 sg13g2_nor2_2 _4693_ (.A(net2271),
    .B(net2211),
    .Y(_0168_));
 sg13g2_nand2_2 _4694_ (.Y(_0169_),
    .A(net2280),
    .B(net2212));
 sg13g2_o21ai_1 _4695_ (.B1(net2279),
    .Y(_0170_),
    .A1(net2214),
    .A2(net2213));
 sg13g2_or2_1 _4696_ (.X(_0171_),
    .B(_0170_),
    .A(net2143));
 sg13g2_nor2_1 _4697_ (.A(_2394_),
    .B(_0164_),
    .Y(_0172_));
 sg13g2_a21oi_1 _4698_ (.A1(_0171_),
    .A2(_0172_),
    .Y(_0173_),
    .B1(net2417));
 sg13g2_nand2_1 _4699_ (.Y(_0174_),
    .A(net2282),
    .B(_3182_));
 sg13g2_nor2_1 _4700_ (.A(net2143),
    .B(_2787_),
    .Y(_0175_));
 sg13g2_a221oi_1 _4701_ (.B2(_0175_),
    .C1(net2430),
    .B1(_0174_),
    .A1(net2070),
    .Y(_0176_),
    .A2(_3125_));
 sg13g2_nor3_2 _4702_ (.A(net2142),
    .B(net2254),
    .C(_3549_),
    .Y(_0177_));
 sg13g2_a21oi_1 _4703_ (.A1(_3528_),
    .A2(_0159_),
    .Y(_0178_),
    .B1(_0177_));
 sg13g2_a21oi_1 _4704_ (.A1(net2048),
    .A2(_0178_),
    .Y(_0179_),
    .B1(net2541));
 sg13g2_nor4_2 _4705_ (.A(net2504),
    .B(_0173_),
    .C(_0176_),
    .Y(_0180_),
    .D(_0179_));
 sg13g2_nand3_1 _4706_ (.B(net2221),
    .C(net2072),
    .A(net2163),
    .Y(_0181_));
 sg13g2_a21oi_1 _4707_ (.A1(_0131_),
    .A2(_0181_),
    .Y(_0182_),
    .B1(net2419));
 sg13g2_nand2_2 _4708_ (.Y(_0183_),
    .A(net2504),
    .B(net2042));
 sg13g2_nor3_1 _4709_ (.A(_3135_),
    .B(_0130_),
    .C(_0183_),
    .Y(_0184_));
 sg13g2_a21oi_1 _4710_ (.A1(_0181_),
    .A2(_0184_),
    .Y(_0185_),
    .B1(net2334));
 sg13g2_nor2_1 _4711_ (.A(net2429),
    .B(_0134_),
    .Y(_0186_));
 sg13g2_nor3_1 _4712_ (.A(_0182_),
    .B(_0185_),
    .C(_0186_),
    .Y(_0187_));
 sg13g2_nor3_1 _4713_ (.A(net2390),
    .B(_0180_),
    .C(_0187_),
    .Y(_0188_));
 sg13g2_o21ai_1 _4714_ (.B1(net2038),
    .Y(_0189_),
    .A1(_0163_),
    .A2(_0188_));
 sg13g2_and2_1 _4715_ (.A(net2587),
    .B(_3278_),
    .X(_0190_));
 sg13g2_a221oi_1 _4716_ (.B2(net2587),
    .C1(_3246_),
    .B1(_3276_),
    .A1(_3251_),
    .Y(_0191_),
    .A2(net2022));
 sg13g2_nor2_1 _4717_ (.A(net2326),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_a22oi_1 _4718_ (.Y(_0193_),
    .B1(_3269_),
    .B2(_3419_),
    .A2(_3257_),
    .A1(net2510));
 sg13g2_and3_1 _4719_ (.X(_0194_),
    .A(_3249_),
    .B(_3277_),
    .C(_3283_));
 sg13g2_o21ai_1 _4720_ (.B1(_0193_),
    .Y(_0195_),
    .A1(net2313),
    .A2(_0194_));
 sg13g2_o21ai_1 _4721_ (.B1(net2379),
    .Y(_0196_),
    .A1(_0192_),
    .A2(_0195_));
 sg13g2_nor3_1 _4722_ (.A(net2528),
    .B(_3154_),
    .C(_3425_),
    .Y(_0197_));
 sg13g2_a21oi_2 _4723_ (.B1(net2199),
    .Y(_0198_),
    .A2(_0197_),
    .A1(_3027_));
 sg13g2_a21oi_1 _4724_ (.A1(net2462),
    .A2(net2021),
    .Y(_0199_),
    .B1(net2442));
 sg13g2_o21ai_1 _4725_ (.B1(_3268_),
    .Y(_0200_),
    .A1(_3294_),
    .A2(_0199_));
 sg13g2_a21oi_1 _4726_ (.A1(net2195),
    .A2(_0200_),
    .Y(_0201_),
    .B1(_0198_));
 sg13g2_a21oi_1 _4727_ (.A1(_0196_),
    .A2(_0201_),
    .Y(_0202_),
    .B1(net2294));
 sg13g2_nand2_2 _4728_ (.Y(_0203_),
    .A(net1979),
    .B(_3375_));
 sg13g2_or3_1 _4729_ (.A(net2560),
    .B(_3095_),
    .C(net2009),
    .X(_0204_));
 sg13g2_a21o_1 _4730_ (.A2(_0204_),
    .A1(_3032_),
    .B1(net2314),
    .X(_0205_));
 sg13g2_nand2_2 _4731_ (.Y(_0206_),
    .A(net2136),
    .B(_3021_));
 sg13g2_nand2_1 _4732_ (.Y(_0207_),
    .A(_3034_),
    .B(_0206_));
 sg13g2_o21ai_1 _4733_ (.B1(net2102),
    .Y(_0208_),
    .A1(net2349),
    .A2(net2079));
 sg13g2_a21oi_2 _4734_ (.B1(net2138),
    .Y(_0209_),
    .A2(_2075_),
    .A1(net2345));
 sg13g2_nand2_2 _4735_ (.Y(_0210_),
    .A(net2374),
    .B(net2067));
 sg13g2_nor2_1 _4736_ (.A(net2128),
    .B(_3420_),
    .Y(_0211_));
 sg13g2_a22oi_1 _4737_ (.Y(_0212_),
    .B1(_0210_),
    .B2(_0211_),
    .A2(_3461_),
    .A1(_3151_));
 sg13g2_o21ai_1 _4738_ (.B1(_0212_),
    .Y(_0213_),
    .A1(_3035_),
    .A2(_3062_));
 sg13g2_a221oi_1 _4739_ (.B2(net2332),
    .C1(_0213_),
    .B1(_0209_),
    .A1(net2306),
    .Y(_0214_),
    .A2(_0207_));
 sg13g2_nor2_1 _4740_ (.A(net2585),
    .B(_3053_),
    .Y(_0215_));
 sg13g2_nor2_2 _4741_ (.A(net2091),
    .B(_3564_),
    .Y(_0216_));
 sg13g2_nand2_1 _4742_ (.Y(_0217_),
    .A(net2135),
    .B(_3565_));
 sg13g2_mux2_2 _4743_ (.A0(net2081),
    .A1(_3564_),
    .S(net2135),
    .X(_0218_));
 sg13g2_nor2_1 _4744_ (.A(net2563),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_o21ai_1 _4745_ (.B1(net2339),
    .Y(_0220_),
    .A1(_0215_),
    .A2(_0219_));
 sg13g2_nor2_1 _4746_ (.A(net2501),
    .B(net2578),
    .Y(_0221_));
 sg13g2_or2_1 _4747_ (.X(_0222_),
    .B(_0218_),
    .A(net2308));
 sg13g2_and4_1 _4748_ (.A(net2379),
    .B(_0214_),
    .C(_0220_),
    .D(_0222_),
    .X(_0223_));
 sg13g2_nand2_2 _4749_ (.Y(_0224_),
    .A(net2571),
    .B(net2353));
 sg13g2_o21ai_1 _4750_ (.B1(net2318),
    .Y(_0225_),
    .A1(_3176_),
    .A2(_0209_));
 sg13g2_a21oi_1 _4751_ (.A1(net2278),
    .A2(_3223_),
    .Y(_0226_),
    .B1(net2149));
 sg13g2_o21ai_1 _4752_ (.B1(net2103),
    .Y(_0227_),
    .A1(net2257),
    .A2(_3224_));
 sg13g2_o21ai_1 _4753_ (.B1(net2306),
    .Y(_0228_),
    .A1(_0140_),
    .A2(_0226_));
 sg13g2_nor2_2 _4754_ (.A(net2138),
    .B(_0167_),
    .Y(_0229_));
 sg13g2_or2_2 _4755_ (.X(_0230_),
    .B(_0167_),
    .A(net2148));
 sg13g2_o21ai_1 _4756_ (.B1(net2309),
    .Y(_0231_),
    .A1(_0140_),
    .A2(_0229_));
 sg13g2_nand4_1 _4757_ (.B(_0225_),
    .C(_0228_),
    .A(net2391),
    .Y(_0232_),
    .D(_0231_));
 sg13g2_a21oi_1 _4758_ (.A1(_3286_),
    .A2(_0230_),
    .Y(_0233_),
    .B1(net2567));
 sg13g2_o21ai_1 _4759_ (.B1(net2332),
    .Y(_0234_),
    .A1(_3287_),
    .A2(_0233_));
 sg13g2_a21oi_2 _4760_ (.B1(net2487),
    .Y(_0235_),
    .A2(_0230_),
    .A1(_3286_));
 sg13g2_nand2_1 _4761_ (.Y(_0236_),
    .A(net2527),
    .B(_0235_));
 sg13g2_a221oi_1 _4762_ (.B2(net2526),
    .C1(_0232_),
    .B1(_0235_),
    .A1(net2223),
    .Y(_0237_),
    .A2(_3061_));
 sg13g2_a221oi_1 _4763_ (.B2(_0237_),
    .C1(net1983),
    .B1(_0234_),
    .A1(_0205_),
    .Y(_0238_),
    .A2(_0223_));
 sg13g2_nor3_2 _4764_ (.A(_0202_),
    .B(_0203_),
    .C(_0238_),
    .Y(_0239_));
 sg13g2_a221oi_1 _4765_ (.B2(_0239_),
    .C1(net1976),
    .B1(_0189_),
    .A1(_3617_),
    .Y(_0240_),
    .A2(_0129_));
 sg13g2_nor3_1 _4766_ (.A(_3504_),
    .B(_3506_),
    .C(_0240_),
    .Y(_0241_));
 sg13g2_nand3_1 _4767_ (.B(_2691_),
    .C(_3018_),
    .A(net2121),
    .Y(_0242_));
 sg13g2_nor2_1 _4768_ (.A(net2569),
    .B(_2797_),
    .Y(_0243_));
 sg13g2_a21oi_1 _4769_ (.A1(net2116),
    .A2(net2066),
    .Y(_0244_),
    .B1(net2592));
 sg13g2_a22oi_1 _4770_ (.Y(_0245_),
    .B1(_0244_),
    .B2(net2043),
    .A2(_0243_),
    .A1(_0242_));
 sg13g2_o21ai_1 _4771_ (.B1(net2531),
    .Y(_0246_),
    .A1(_3327_),
    .A2(_0245_));
 sg13g2_nand3_1 _4772_ (.B(_3018_),
    .C(net2065),
    .A(net2117),
    .Y(_0247_));
 sg13g2_nand4_1 _4773_ (.B(_3322_),
    .C(_0181_),
    .A(net2043),
    .Y(_0248_),
    .D(_0247_));
 sg13g2_nor2_1 _4774_ (.A(_2941_),
    .B(_3017_),
    .Y(_0249_));
 sg13g2_o21ai_1 _4775_ (.B1(net2163),
    .Y(_0250_),
    .A1(net2072),
    .A2(_3320_));
 sg13g2_o21ai_1 _4776_ (.B1(_0250_),
    .Y(_0251_),
    .A1(_2941_),
    .A2(_3017_));
 sg13g2_a221oi_1 _4777_ (.B2(net2444),
    .C1(net2513),
    .B1(_0251_),
    .A1(net2425),
    .Y(_0252_),
    .A2(_0248_));
 sg13g2_nand2_1 _4778_ (.Y(_0253_),
    .A(net2120),
    .B(_3342_));
 sg13g2_a21oi_1 _4779_ (.A1(_1811_),
    .A2(_3343_),
    .Y(_0254_),
    .B1(net2164));
 sg13g2_nand2_1 _4780_ (.Y(_0255_),
    .A(net2121),
    .B(_3350_));
 sg13g2_nand2_1 _4781_ (.Y(_0256_),
    .A(_3388_),
    .B(_0255_));
 sg13g2_nand3_1 _4782_ (.B(net2246),
    .C(_3018_),
    .A(net2288),
    .Y(_0257_));
 sg13g2_nor3_2 _4783_ (.A(net2265),
    .B(_3017_),
    .C(_3151_),
    .Y(_0258_));
 sg13g2_nor3_1 _4784_ (.A(net2169),
    .B(net2054),
    .C(_0258_),
    .Y(_0259_));
 sg13g2_nand3_1 _4785_ (.B(net2071),
    .C(_3321_),
    .A(net2168),
    .Y(_0260_));
 sg13g2_nor2b_1 _4786_ (.A(_0259_),
    .B_N(_0260_),
    .Y(_0261_));
 sg13g2_a21oi_1 _4787_ (.A1(_3201_),
    .A2(_3416_),
    .Y(_0262_),
    .B1(net2404));
 sg13g2_a221oi_1 _4788_ (.B2(net2444),
    .C1(_0262_),
    .B1(_0256_),
    .A1(net2548),
    .Y(_0263_),
    .A2(_3368_));
 sg13g2_a221oi_1 _4789_ (.B2(net2477),
    .C1(net2495),
    .B1(_0261_),
    .A1(net2343),
    .Y(_0264_),
    .A2(_0254_));
 sg13g2_a221oi_1 _4790_ (.B2(_0264_),
    .C1(net2382),
    .B1(_0263_),
    .A1(_0246_),
    .Y(_0265_),
    .A2(_0252_));
 sg13g2_nand2_2 _4791_ (.Y(_0266_),
    .A(net2501),
    .B(net2421));
 sg13g2_o21ai_1 _4792_ (.B1(net2161),
    .Y(_0267_),
    .A1(net2248),
    .A2(_3329_));
 sg13g2_nor2b_1 _4793_ (.A(_3519_),
    .B_N(_0267_),
    .Y(_0268_));
 sg13g2_nor2_1 _4794_ (.A(_0266_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_nand2_1 _4795_ (.Y(_0270_),
    .A(net2101),
    .B(_2826_));
 sg13g2_o21ai_1 _4796_ (.B1(net2129),
    .Y(_0271_),
    .A1(_2826_),
    .A2(net2055));
 sg13g2_nor2_1 _4797_ (.A(_2787_),
    .B(_0271_),
    .Y(_0272_));
 sg13g2_o21ai_1 _4798_ (.B1(net2226),
    .Y(_0273_),
    .A1(net2258),
    .A2(net2361));
 sg13g2_nor3_2 _4799_ (.A(net2105),
    .B(net2350),
    .C(_0273_),
    .Y(_0274_));
 sg13g2_nor4_2 _4800_ (.A(net2497),
    .B(net2437),
    .C(_0272_),
    .Y(_0275_),
    .D(_0274_));
 sg13g2_o21ai_1 _4801_ (.B1(net2593),
    .Y(_0276_),
    .A1(net2029),
    .A2(_3335_));
 sg13g2_nand2_2 _4802_ (.Y(_0277_),
    .A(_3129_),
    .B(_0170_));
 sg13g2_nand3_1 _4803_ (.B(net2351),
    .C(_2702_),
    .A(net2246),
    .Y(_0278_));
 sg13g2_a22oi_1 _4804_ (.Y(_0279_),
    .B1(_0278_),
    .B2(net2159),
    .A2(_0277_),
    .A1(net2023));
 sg13g2_a21oi_1 _4805_ (.A1(_0276_),
    .A2(_0279_),
    .Y(_0280_),
    .B1(net2316));
 sg13g2_nor3_1 _4806_ (.A(_0269_),
    .B(_0275_),
    .C(_0280_),
    .Y(_0281_));
 sg13g2_o21ai_1 _4807_ (.B1(net2133),
    .Y(_0282_),
    .A1(net2087),
    .A2(_3082_));
 sg13g2_a21oi_1 _4808_ (.A1(_3317_),
    .A2(_0282_),
    .Y(_0283_),
    .B1(net2570));
 sg13g2_a21oi_1 _4809_ (.A1(_3317_),
    .A2(_0267_),
    .Y(_0284_),
    .B1(net2592));
 sg13g2_or2_1 _4810_ (.X(_0285_),
    .B(_0284_),
    .A(_0283_));
 sg13g2_nand2_1 _4811_ (.Y(_0286_),
    .A(_3090_),
    .B(_0277_));
 sg13g2_nand2_1 _4812_ (.Y(_0287_),
    .A(_3132_),
    .B(_0282_));
 sg13g2_nand2_2 _4813_ (.Y(_0288_),
    .A(net2260),
    .B(net2212));
 sg13g2_nand3_1 _4814_ (.B(net2022),
    .C(_0288_),
    .A(_3160_),
    .Y(_0289_));
 sg13g2_nand4_1 _4815_ (.B(_0282_),
    .C(_0286_),
    .A(_3132_),
    .Y(_0290_),
    .D(_0289_));
 sg13g2_a22oi_1 _4816_ (.Y(_0291_),
    .B1(_0290_),
    .B2(net2329),
    .A2(_0285_),
    .A1(net2340));
 sg13g2_a21oi_1 _4817_ (.A1(_0281_),
    .A2(_0291_),
    .Y(_0292_),
    .B1(net2395));
 sg13g2_or3_2 _4818_ (.A(net2302),
    .B(_0265_),
    .C(_0292_),
    .X(_0293_));
 sg13g2_a21oi_1 _4819_ (.A1(net2013),
    .A2(_3475_),
    .Y(_0294_),
    .B1(_3411_));
 sg13g2_nand3_1 _4820_ (.B(_3169_),
    .C(net2055),
    .A(net2127),
    .Y(_0295_));
 sg13g2_nand2_2 _4821_ (.Y(_0296_),
    .A(net2015),
    .B(net2004));
 sg13g2_nand2_1 _4822_ (.Y(_0297_),
    .A(net2556),
    .B(_0296_));
 sg13g2_nor2_1 _4823_ (.A(net2185),
    .B(net2059),
    .Y(_0298_));
 sg13g2_nand2_1 _4824_ (.Y(_0299_),
    .A(net2131),
    .B(net2057));
 sg13g2_nor2_2 _4825_ (.A(net2258),
    .B(_3223_),
    .Y(_0300_));
 sg13g2_nor2_1 _4826_ (.A(net2001),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_or3_1 _4827_ (.A(net2184),
    .B(net2058),
    .C(_0300_),
    .X(_0302_));
 sg13g2_a22oi_1 _4828_ (.Y(_0303_),
    .B1(_0301_),
    .B2(net2414),
    .A2(_0296_),
    .A1(net2556));
 sg13g2_a22oi_1 _4829_ (.Y(_0304_),
    .B1(_0114_),
    .B2(net2342),
    .A2(_3485_),
    .A1(net2449));
 sg13g2_a21oi_1 _4830_ (.A1(_0303_),
    .A2(_0304_),
    .Y(_0305_),
    .B1(net2499));
 sg13g2_nor3_1 _4831_ (.A(net2292),
    .B(net2239),
    .C(net2209),
    .Y(_0306_));
 sg13g2_nand2_1 _4832_ (.Y(_0307_),
    .A(net2181),
    .B(_0306_));
 sg13g2_nand2_2 _4833_ (.Y(_0308_),
    .A(net2601),
    .B(net2214));
 sg13g2_nand3_1 _4834_ (.B(_0307_),
    .C(_0308_),
    .A(_3388_),
    .Y(_0309_));
 sg13g2_nor3_1 _4835_ (.A(_3366_),
    .B(_3474_),
    .C(_0309_),
    .Y(_0310_));
 sg13g2_mux2_2 _4836_ (.A0(net2242),
    .A1(net2219),
    .S(net2269),
    .X(_0311_));
 sg13g2_nand2b_2 _4837_ (.Y(_0312_),
    .B(net2457),
    .A_N(_0311_));
 sg13g2_a21o_1 _4838_ (.A2(_0312_),
    .A1(net2023),
    .B1(_3368_),
    .X(_0313_));
 sg13g2_a221oi_1 _4839_ (.B2(net2324),
    .C1(net2395),
    .B1(_0313_),
    .A1(net2312),
    .Y(_0314_),
    .A2(_0256_));
 sg13g2_o21ai_1 _4840_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_3040_),
    .A2(_0310_));
 sg13g2_nor3_1 _4841_ (.A(_0294_),
    .B(_0305_),
    .C(_0315_),
    .Y(_0316_));
 sg13g2_nor3_2 _4842_ (.A(net2262),
    .B(net2215),
    .C(_3162_),
    .Y(_0317_));
 sg13g2_nor2_2 _4843_ (.A(net2177),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_or2_2 _4844_ (.X(_0319_),
    .B(_0317_),
    .A(net2178));
 sg13g2_nor2_1 _4845_ (.A(net2060),
    .B(_0319_),
    .Y(_0320_));
 sg13g2_or3_2 _4846_ (.A(net2178),
    .B(net2060),
    .C(_0317_),
    .X(_0321_));
 sg13g2_nand2b_1 _4847_ (.Y(_0322_),
    .B(_0321_),
    .A_N(_3443_));
 sg13g2_nand3_1 _4848_ (.B(_3221_),
    .C(_3397_),
    .A(net2126),
    .Y(_0323_));
 sg13g2_nand2_2 _4849_ (.Y(_0324_),
    .A(net2014),
    .B(net1999));
 sg13g2_a21oi_2 _4850_ (.B1(net2577),
    .Y(_0325_),
    .A2(net1999),
    .A1(net2013));
 sg13g2_and4_1 _4851_ (.A(_3403_),
    .B(net2013),
    .C(_3441_),
    .D(net2004),
    .X(_0326_));
 sg13g2_nand2b_1 _4852_ (.Y(_0327_),
    .B(_0326_),
    .A_N(_0325_));
 sg13g2_nor3_2 _4853_ (.A(net2265),
    .B(net2225),
    .C(net2215),
    .Y(_0328_));
 sg13g2_nor2_2 _4854_ (.A(net2002),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_or3_1 _4855_ (.A(net2184),
    .B(net2058),
    .C(_0328_),
    .X(_0330_));
 sg13g2_nand3_1 _4856_ (.B(_3456_),
    .C(_0330_),
    .A(_3441_),
    .Y(_0331_));
 sg13g2_a21oi_1 _4857_ (.A1(net2340),
    .A2(_0331_),
    .Y(_0332_),
    .B1(net2384));
 sg13g2_a21oi_1 _4858_ (.A1(net2014),
    .A2(net1998),
    .Y(_0333_),
    .B1(net2601));
 sg13g2_nor3_1 _4859_ (.A(_3485_),
    .B(_0296_),
    .C(_0333_),
    .Y(_0334_));
 sg13g2_o21ai_1 _4860_ (.B1(_0332_),
    .Y(_0335_),
    .A1(net2316),
    .A2(_0334_));
 sg13g2_a221oi_1 _4861_ (.B2(_3039_),
    .C1(_0335_),
    .B1(_0327_),
    .A1(net2335),
    .Y(_0336_),
    .A2(_0322_));
 sg13g2_o21ai_1 _4862_ (.B1(net2303),
    .Y(_0337_),
    .A1(_0316_),
    .A2(_0336_));
 sg13g2_nand3_1 _4863_ (.B(_0293_),
    .C(_0337_),
    .A(net2036),
    .Y(_0338_));
 sg13g2_nand4_1 _4864_ (.B(net2292),
    .C(net2211),
    .A(net2131),
    .Y(_0339_),
    .D(_3377_));
 sg13g2_nand2_1 _4865_ (.Y(_0340_),
    .A(_3376_),
    .B(_0339_));
 sg13g2_nand3_1 _4866_ (.B(_3384_),
    .C(_0339_),
    .A(net2019),
    .Y(_0341_));
 sg13g2_nor2_2 _4867_ (.A(_3385_),
    .B(_0340_),
    .Y(_0342_));
 sg13g2_nand3_1 _4868_ (.B(_3384_),
    .C(_0321_),
    .A(_3379_),
    .Y(_0343_));
 sg13g2_a21oi_1 _4869_ (.A1(_3388_),
    .A2(_0339_),
    .Y(_0344_),
    .B1(net2467));
 sg13g2_a21oi_1 _4870_ (.A1(net2534),
    .A2(_0343_),
    .Y(_0345_),
    .B1(_0344_));
 sg13g2_o21ai_1 _4871_ (.B1(_0345_),
    .Y(_0346_),
    .A1(net2534),
    .A2(_0342_));
 sg13g2_nand3_1 _4872_ (.B(net2010),
    .C(_0319_),
    .A(_3416_),
    .Y(_0347_));
 sg13g2_nand3_1 _4873_ (.B(_3418_),
    .C(_0319_),
    .A(_3416_),
    .Y(_0348_));
 sg13g2_a22oi_1 _4874_ (.Y(_0349_),
    .B1(_0348_),
    .B2(net2342),
    .A2(_0347_),
    .A1(net2449));
 sg13g2_nand3_1 _4875_ (.B(_3412_),
    .C(net2003),
    .A(net2017),
    .Y(_0350_));
 sg13g2_a21oi_1 _4876_ (.A1(net2480),
    .A2(_0350_),
    .Y(_0351_),
    .B1(net2497));
 sg13g2_nand2_1 _4877_ (.Y(_0352_),
    .A(_0349_),
    .B(_0351_));
 sg13g2_and3_1 _4878_ (.X(_0353_),
    .A(_3395_),
    .B(_3404_),
    .C(net2003));
 sg13g2_nand2_2 _4879_ (.Y(_0354_),
    .A(net2017),
    .B(net1999));
 sg13g2_a22oi_1 _4880_ (.Y(_0355_),
    .B1(_0354_),
    .B2(net2533),
    .A2(_3407_),
    .A1(_1371_));
 sg13g2_a21oi_1 _4881_ (.A1(_0353_),
    .A2(_0355_),
    .Y(_0356_),
    .B1(net2398));
 sg13g2_a21o_1 _4882_ (.A2(_0347_),
    .A1(net2198),
    .B1(net2296),
    .X(_0357_));
 sg13g2_a221oi_1 _4883_ (.B2(_0356_),
    .C1(_0357_),
    .B1(_0352_),
    .A1(net2206),
    .Y(_0358_),
    .A2(_0346_));
 sg13g2_nand4_1 _4884_ (.B(net2017),
    .C(_3404_),
    .A(net2534),
    .Y(_0359_),
    .D(net1998));
 sg13g2_nor3_1 _4885_ (.A(net2532),
    .B(_3406_),
    .C(_0354_),
    .Y(_0360_));
 sg13g2_o21ai_1 _4886_ (.B1(net2206),
    .Y(_0361_),
    .A1(_0325_),
    .A2(_0359_));
 sg13g2_o21ai_1 _4887_ (.B1(net2296),
    .Y(_0362_),
    .A1(_0360_),
    .A2(_0361_));
 sg13g2_nand3_1 _4888_ (.B(net2014),
    .C(net1998),
    .A(_3404_),
    .Y(_0363_));
 sg13g2_nand3_1 _4889_ (.B(net2010),
    .C(net2000),
    .A(net2027),
    .Y(_0364_));
 sg13g2_a22oi_1 _4890_ (.Y(_0365_),
    .B1(_0364_),
    .B2(net2428),
    .A2(_0363_),
    .A1(net2448));
 sg13g2_nand2_1 _4891_ (.Y(_0366_),
    .A(_3367_),
    .B(net2010));
 sg13g2_nand3_1 _4892_ (.B(net2010),
    .C(net2000),
    .A(_3367_),
    .Y(_0367_));
 sg13g2_a22oi_1 _4893_ (.Y(_0368_),
    .B1(_0367_),
    .B2(net2534),
    .A2(_3385_),
    .A1(net2482));
 sg13g2_nand2_1 _4894_ (.Y(_0369_),
    .A(_0365_),
    .B(_0368_));
 sg13g2_nand3_1 _4895_ (.B(_3441_),
    .C(net2000),
    .A(_3427_),
    .Y(_0370_));
 sg13g2_mux2_1 _4896_ (.A0(_0322_),
    .A1(_0370_),
    .S(net2517),
    .X(_0371_));
 sg13g2_a221oi_1 _4897_ (.B2(net2384),
    .C1(_0362_),
    .B1(_0371_),
    .A1(net2197),
    .Y(_0372_),
    .A2(_0369_));
 sg13g2_nor3_2 _4898_ (.A(net2036),
    .B(_0358_),
    .C(_0372_),
    .Y(_0373_));
 sg13g2_nor2_1 _4899_ (.A(_3214_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_a21oi_1 _4900_ (.A1(_2734_),
    .A2(net2042),
    .Y(_0375_),
    .B1(net2578));
 sg13g2_nor3_2 _4901_ (.A(net2116),
    .B(net2460),
    .C(_0311_),
    .Y(_0376_));
 sg13g2_xnor2_1 _4902_ (.Y(_0377_),
    .A(net2090),
    .B(_0312_));
 sg13g2_a21oi_1 _4903_ (.A1(_2872_),
    .A2(_0377_),
    .Y(_0378_),
    .B1(_2892_));
 sg13g2_o21ai_1 _4904_ (.B1(net2521),
    .Y(_0379_),
    .A1(_0375_),
    .A2(_0378_));
 sg13g2_a22oi_1 _4905_ (.Y(_0380_),
    .B1(_3422_),
    .B2(net2232),
    .A2(_2744_),
    .A1(net2336));
 sg13g2_a21oi_1 _4906_ (.A1(_2339_),
    .A2(_2863_),
    .Y(_0381_),
    .B1(net2521));
 sg13g2_a21oi_1 _4907_ (.A1(_3160_),
    .A2(_3606_),
    .Y(_0382_),
    .B1(net2501));
 sg13g2_a21oi_1 _4908_ (.A1(net2521),
    .A2(_2482_),
    .Y(_0383_),
    .B1(_0381_));
 sg13g2_a221oi_1 _4909_ (.B2(_0383_),
    .C1(net2388),
    .B1(_0382_),
    .A1(_0379_),
    .Y(_0384_),
    .A2(_0380_));
 sg13g2_nand3_1 _4910_ (.B(net2230),
    .C(net2077),
    .A(net2161),
    .Y(_0385_));
 sg13g2_nand3_1 _4911_ (.B(_3157_),
    .C(_0385_),
    .A(_3136_),
    .Y(_0386_));
 sg13g2_nand3_1 _4912_ (.B(net2357),
    .C(net2077),
    .A(net2162),
    .Y(_0387_));
 sg13g2_nand4_1 _4913_ (.B(_3136_),
    .C(_3138_),
    .A(_3115_),
    .Y(_0388_),
    .D(_0387_));
 sg13g2_a22oi_1 _4914_ (.Y(_0389_),
    .B1(_0388_),
    .B2(net2441),
    .A2(_0386_),
    .A1(net2423));
 sg13g2_o21ai_1 _4915_ (.B1(_0389_),
    .Y(_0390_),
    .A1(net2403),
    .A2(_3537_));
 sg13g2_o21ai_1 _4916_ (.B1(net2204),
    .Y(_0391_),
    .A1(_3188_),
    .A2(_0390_));
 sg13g2_nand3_1 _4917_ (.B(_3176_),
    .C(_3200_),
    .A(net2582),
    .Y(_0392_));
 sg13g2_nor3_1 _4918_ (.A(_3149_),
    .B(net2028),
    .C(_3196_),
    .Y(_0393_));
 sg13g2_a21oi_1 _4919_ (.A1(_0392_),
    .A2(_0393_),
    .Y(_0394_),
    .B1(_3290_));
 sg13g2_o21ai_1 _4920_ (.B1(net2581),
    .Y(_0395_),
    .A1(_3194_),
    .A2(_3196_));
 sg13g2_a21oi_2 _4921_ (.B1(_3194_),
    .Y(_0396_),
    .A2(_0154_),
    .A1(_2647_));
 sg13g2_a221oi_1 _4922_ (.B2(_0396_),
    .C1(_3460_),
    .B1(_3203_),
    .A1(_1129_),
    .Y(_0397_),
    .A2(_1294_));
 sg13g2_nand2_2 _4923_ (.Y(_0398_),
    .A(net2079),
    .B(net2070));
 sg13g2_o21ai_1 _4924_ (.B1(net2137),
    .Y(_0399_),
    .A1(_2075_),
    .A2(net2073));
 sg13g2_nor2_1 _4925_ (.A(_2394_),
    .B(_2713_),
    .Y(_0400_));
 sg13g2_a21oi_1 _4926_ (.A1(_0399_),
    .A2(_0400_),
    .Y(_0401_),
    .B1(_0110_));
 sg13g2_nor3_1 _4927_ (.A(net2295),
    .B(_0397_),
    .C(_0401_),
    .Y(_0402_));
 sg13g2_nand3_1 _4928_ (.B(_0393_),
    .C(_0395_),
    .A(_0392_),
    .Y(_0403_));
 sg13g2_nand2_1 _4929_ (.Y(_0404_),
    .A(_3289_),
    .B(_0403_));
 sg13g2_nand3_1 _4930_ (.B(_0402_),
    .C(_0404_),
    .A(_0391_),
    .Y(_0405_));
 sg13g2_a21oi_1 _4931_ (.A1(_3043_),
    .A2(_3060_),
    .Y(_0406_),
    .B1(net2526));
 sg13g2_a21oi_1 _4932_ (.A1(_3042_),
    .A2(_3057_),
    .Y(_0407_),
    .B1(net2402));
 sg13g2_nor4_1 _4933_ (.A(net2506),
    .B(_3058_),
    .C(_0406_),
    .D(_0407_),
    .Y(_0408_));
 sg13g2_a21oi_1 _4934_ (.A1(_0206_),
    .A2(_0270_),
    .Y(_0409_),
    .B1(net2431));
 sg13g2_nor2_1 _4935_ (.A(net2442),
    .B(_3060_),
    .Y(_0410_));
 sg13g2_o21ai_1 _4936_ (.B1(net2506),
    .Y(_0411_),
    .A1(net2416),
    .A2(_3379_));
 sg13g2_nor3_1 _4937_ (.A(_0409_),
    .B(_0410_),
    .C(_0411_),
    .Y(_0412_));
 sg13g2_or3_1 _4938_ (.A(net2391),
    .B(_0408_),
    .C(_0412_),
    .X(_0413_));
 sg13g2_nor3_1 _4939_ (.A(net2440),
    .B(_3030_),
    .C(_3093_),
    .Y(_0414_));
 sg13g2_nor2_1 _4940_ (.A(net2194),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_o21ai_1 _4941_ (.B1(net2137),
    .Y(_0416_),
    .A1(net2070),
    .A2(_3174_));
 sg13g2_nand3_1 _4942_ (.B(_3083_),
    .C(_0416_),
    .A(net2440),
    .Y(_0417_));
 sg13g2_nand2_2 _4943_ (.Y(_0418_),
    .A(net2176),
    .B(_3101_));
 sg13g2_o21ai_1 _4944_ (.B1(_2734_),
    .Y(_0419_),
    .A1(net2235),
    .A2(_0418_));
 sg13g2_nand3_1 _4945_ (.B(_3108_),
    .C(_0419_),
    .A(_3105_),
    .Y(_0420_));
 sg13g2_a221oi_1 _4946_ (.B2(net2202),
    .C1(net2301),
    .B1(_0420_),
    .A1(_0415_),
    .Y(_0421_),
    .A2(_0417_));
 sg13g2_a21oi_1 _4947_ (.A1(_0413_),
    .A2(_0421_),
    .Y(_0422_),
    .B1(net2035));
 sg13g2_o21ai_1 _4948_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_0384_),
    .A2(_0405_));
 sg13g2_nand2_1 _4949_ (.Y(_0424_),
    .A(net2463),
    .B(_3296_));
 sg13g2_nand3_1 _4950_ (.B(net2021),
    .C(_3295_),
    .A(net2312),
    .Y(_0425_));
 sg13g2_nor2_2 _4951_ (.A(net2487),
    .B(net2402),
    .Y(_0426_));
 sg13g2_nor2_2 _4952_ (.A(net2260),
    .B(_3221_),
    .Y(_0427_));
 sg13g2_nor2_2 _4953_ (.A(net2154),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_or2_2 _4954_ (.X(_0429_),
    .B(_0427_),
    .A(net2154));
 sg13g2_o21ai_1 _4955_ (.B1(_0426_),
    .Y(_0430_),
    .A1(_3246_),
    .A2(_0428_));
 sg13g2_nand2_1 _4956_ (.Y(_0431_),
    .A(net2332),
    .B(_3278_));
 sg13g2_nand2b_1 _4957_ (.Y(_0432_),
    .B(_3420_),
    .A_N(_3272_));
 sg13g2_nand4_1 _4958_ (.B(_0430_),
    .C(_0431_),
    .A(_0425_),
    .Y(_0433_),
    .D(_0432_));
 sg13g2_nor2_2 _4959_ (.A(net2177),
    .B(_0168_),
    .Y(_0434_));
 sg13g2_nor3_1 _4960_ (.A(net2473),
    .B(net2020),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_o21ai_1 _4961_ (.B1(net2195),
    .Y(_0436_),
    .A1(net2462),
    .A2(_3278_));
 sg13g2_o21ai_1 _4962_ (.B1(net2475),
    .Y(_0437_),
    .A1(_3233_),
    .A2(net2020));
 sg13g2_o21ai_1 _4963_ (.B1(net2344),
    .Y(_0438_),
    .A1(_3237_),
    .A2(_3238_));
 sg13g2_nand3_1 _4964_ (.B(_0437_),
    .C(_0438_),
    .A(_3242_),
    .Y(_0439_));
 sg13g2_a22oi_1 _4965_ (.Y(_0440_),
    .B1(_0439_),
    .B2(net2203),
    .A2(_0433_),
    .A1(net2378));
 sg13g2_o21ai_1 _4966_ (.B1(_0440_),
    .Y(_0441_),
    .A1(_0435_),
    .A2(_0436_));
 sg13g2_a221oi_1 _4967_ (.B2(_3300_),
    .C1(net1979),
    .B1(_0441_),
    .A1(net1984),
    .Y(_0442_),
    .A2(_0424_));
 sg13g2_a221oi_1 _4968_ (.B2(_0442_),
    .C1(_3308_),
    .B1(_0423_),
    .A1(_0338_),
    .Y(_0443_),
    .A2(_0374_));
 sg13g2_o21ai_1 _4969_ (.B1(net2563),
    .Y(_0444_),
    .A1(_2922_),
    .A2(_3274_));
 sg13g2_nor3_2 _4970_ (.A(net2139),
    .B(_2922_),
    .C(_0167_),
    .Y(_0445_));
 sg13g2_o21ai_1 _4971_ (.B1(_0444_),
    .Y(_0446_),
    .A1(net2022),
    .A2(_0445_));
 sg13g2_a21oi_1 _4972_ (.A1(_3383_),
    .A2(_0446_),
    .Y(_0447_),
    .B1(net2539));
 sg13g2_o21ai_1 _4973_ (.B1(net2202),
    .Y(_0448_),
    .A1(_3579_),
    .A2(_0447_));
 sg13g2_and3_1 _4974_ (.X(_0449_),
    .A(net2542),
    .B(_3195_),
    .C(_3611_));
 sg13g2_a21oi_2 _4975_ (.B1(net2096),
    .Y(_0450_),
    .A2(_3103_),
    .A1(net2079));
 sg13g2_nor2_2 _4976_ (.A(net2279),
    .B(net2352),
    .Y(_0451_));
 sg13g2_nor2_2 _4977_ (.A(net2282),
    .B(net2208),
    .Y(_0452_));
 sg13g2_nor3_1 _4978_ (.A(net2561),
    .B(net2275),
    .C(net2208),
    .Y(_0453_));
 sg13g2_nor4_1 _4979_ (.A(net2542),
    .B(_2394_),
    .C(_0450_),
    .D(_0453_),
    .Y(_0454_));
 sg13g2_a21oi_1 _4980_ (.A1(net2240),
    .A2(_2713_),
    .Y(_0455_),
    .B1(net2504));
 sg13g2_o21ai_1 _4981_ (.B1(_0455_),
    .Y(_0456_),
    .A1(_0449_),
    .A2(_0454_));
 sg13g2_or2_1 _4982_ (.X(_0457_),
    .B(_3605_),
    .A(_2328_));
 sg13g2_o21ai_1 _4983_ (.B1(net2439),
    .Y(_0458_),
    .A1(_2086_),
    .A2(_3601_));
 sg13g2_o21ai_1 _4984_ (.B1(net2141),
    .Y(_0459_),
    .A1(net2087),
    .A2(_3548_));
 sg13g2_o21ai_1 _4985_ (.B1(_0459_),
    .Y(_0460_),
    .A1(net2140),
    .A2(_3312_));
 sg13g2_a221oi_1 _4986_ (.B2(net2472),
    .C1(net2485),
    .B1(_0460_),
    .A1(net2344),
    .Y(_0461_),
    .A2(_0457_));
 sg13g2_a21oi_1 _4987_ (.A1(_0458_),
    .A2(_0461_),
    .Y(_0462_),
    .B1(net2388));
 sg13g2_o21ai_1 _4988_ (.B1(net2439),
    .Y(_0463_),
    .A1(net2034),
    .A2(_3581_));
 sg13g2_a21oi_2 _4989_ (.B1(net2099),
    .Y(_0464_),
    .A2(_3164_),
    .A1(_3099_));
 sg13g2_o21ai_1 _4990_ (.B1(net2408),
    .Y(_0465_),
    .A1(_3587_),
    .A2(_0464_));
 sg13g2_o21ai_1 _4991_ (.B1(net2470),
    .Y(_0466_),
    .A1(_2086_),
    .A2(_3601_));
 sg13g2_o21ai_1 _4992_ (.B1(net2421),
    .Y(_0467_),
    .A1(_3104_),
    .A2(_3587_));
 sg13g2_nand4_1 _4993_ (.B(_0465_),
    .C(_0466_),
    .A(_0463_),
    .Y(_0468_),
    .D(_0467_));
 sg13g2_a221oi_1 _4994_ (.B2(net2196),
    .C1(net2295),
    .B1(_0468_),
    .A1(_0456_),
    .Y(_0469_),
    .A2(_0462_));
 sg13g2_nand4_1 _4995_ (.B(net2026),
    .C(_3550_),
    .A(net2048),
    .Y(_0470_),
    .D(_3551_));
 sg13g2_nor2_2 _4996_ (.A(net2289),
    .B(_3222_),
    .Y(_0471_));
 sg13g2_nand2_2 _4997_ (.Y(_0472_),
    .A(net2261),
    .B(_3221_));
 sg13g2_nor2_2 _4998_ (.A(net2159),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_nand2_2 _4999_ (.Y(_0474_),
    .A(net2105),
    .B(_0471_));
 sg13g2_nand4_1 _5000_ (.B(_3550_),
    .C(_3551_),
    .A(net2011),
    .Y(_0475_),
    .D(net1997));
 sg13g2_nand2_1 _5001_ (.Y(_0476_),
    .A(net2410),
    .B(_0475_));
 sg13g2_a21o_1 _5002_ (.A2(_3547_),
    .A1(net2222),
    .B1(_3541_),
    .X(_0477_));
 sg13g2_a22oi_1 _5003_ (.Y(_0478_),
    .B1(_0477_),
    .B2(net2443),
    .A2(_0470_),
    .A1(net2425));
 sg13g2_nand3_1 _5004_ (.B(_0476_),
    .C(_0478_),
    .A(_3538_),
    .Y(_0479_));
 sg13g2_nor3_2 _5005_ (.A(net2284),
    .B(net2225),
    .C(net2213),
    .Y(_0480_));
 sg13g2_nor2_1 _5006_ (.A(net2112),
    .B(_0165_),
    .Y(_0481_));
 sg13g2_nand2_1 _5007_ (.Y(_0482_),
    .A(net2162),
    .B(_0166_));
 sg13g2_nor2_1 _5008_ (.A(_0480_),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_nor3_1 _5009_ (.A(net2584),
    .B(net2363),
    .C(net2357),
    .Y(_0484_));
 sg13g2_nor2_1 _5010_ (.A(net2543),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_a21oi_2 _5011_ (.B1(net2163),
    .Y(_0486_),
    .A2(_3340_),
    .A1(net2220));
 sg13g2_nor4_1 _5012_ (.A(net2541),
    .B(_0483_),
    .C(_0484_),
    .D(_0486_),
    .Y(_0487_));
 sg13g2_nor2_1 _5013_ (.A(net2194),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_a221oi_1 _5014_ (.B2(_0464_),
    .C1(net2417),
    .B1(_0166_),
    .A1(net2099),
    .Y(_0489_),
    .A2(_3147_));
 sg13g2_a22oi_1 _5015_ (.Y(_0490_),
    .B1(_3620_),
    .B2(_0489_),
    .A2(_3537_),
    .A1(net2441));
 sg13g2_o21ai_1 _5016_ (.B1(net2552),
    .Y(_0491_),
    .A1(net2115),
    .A2(_3398_));
 sg13g2_nand2_1 _5017_ (.Y(_0492_),
    .A(net2076),
    .B(_3171_));
 sg13g2_a221oi_1 _5018_ (.B2(net2033),
    .C1(_0491_),
    .B1(_0492_),
    .A1(net2161),
    .Y(_0493_),
    .A2(_3512_));
 sg13g2_nand2_2 _5019_ (.Y(_0494_),
    .A(net2122),
    .B(_0328_));
 sg13g2_nand2_1 _5020_ (.Y(_0495_),
    .A(net2043),
    .B(_0494_));
 sg13g2_o21ai_1 _5021_ (.B1(net2531),
    .Y(_0496_),
    .A1(net2592),
    .A2(net2374));
 sg13g2_nor3_1 _5022_ (.A(_3327_),
    .B(_0495_),
    .C(_0496_),
    .Y(_0497_));
 sg13g2_o21ai_1 _5023_ (.B1(_3522_),
    .Y(_0498_),
    .A1(_0493_),
    .A2(_0497_));
 sg13g2_a21oi_1 _5024_ (.A1(_3122_),
    .A2(net2063),
    .Y(_0499_),
    .B1(_0482_));
 sg13g2_o21ai_1 _5025_ (.B1(net2569),
    .Y(_0500_),
    .A1(_0486_),
    .A2(_0499_));
 sg13g2_nand2_1 _5026_ (.Y(_0501_),
    .A(_3029_),
    .B(_3124_));
 sg13g2_a21oi_1 _5027_ (.A1(net2074),
    .A2(_3124_),
    .Y(_0502_),
    .B1(net2569));
 sg13g2_a221oi_1 _5028_ (.B2(_3269_),
    .C1(net2331),
    .B1(_0502_),
    .A1(net2592),
    .Y(_0503_),
    .A2(_3316_));
 sg13g2_a22oi_1 _5029_ (.Y(_0504_),
    .B1(_0501_),
    .B2(_3027_),
    .A2(_3316_),
    .A1(net2569));
 sg13g2_nor2_1 _5030_ (.A(_2537_),
    .B(_0283_),
    .Y(_0505_));
 sg13g2_a22oi_1 _5031_ (.Y(_0506_),
    .B1(_0504_),
    .B2(_0505_),
    .A2(_0503_),
    .A1(_0500_));
 sg13g2_nand3_1 _5032_ (.B(_0498_),
    .C(_0506_),
    .A(net2382),
    .Y(_0507_));
 sg13g2_a221oi_1 _5033_ (.B2(_0490_),
    .C1(net2301),
    .B1(_0488_),
    .A1(net2204),
    .Y(_0508_),
    .A2(_0479_));
 sg13g2_a221oi_1 _5034_ (.B2(_0508_),
    .C1(net2035),
    .B1(_0507_),
    .A1(_0448_),
    .Y(_0509_),
    .A2(_0469_));
 sg13g2_nor2_1 _5035_ (.A(net2316),
    .B(_0342_),
    .Y(_0510_));
 sg13g2_o21ai_1 _5036_ (.B1(net2499),
    .Y(_0511_),
    .A1(net2420),
    .A2(_3379_));
 sg13g2_a21oi_1 _5037_ (.A1(net2556),
    .A2(_0341_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_nor2_1 _5038_ (.A(_2306_),
    .B(net2001),
    .Y(_0513_));
 sg13g2_nand3_1 _5039_ (.B(net2078),
    .C(net2056),
    .A(net2127),
    .Y(_0514_));
 sg13g2_o21ai_1 _5040_ (.B1(net2448),
    .Y(_0515_),
    .A1(_3632_),
    .A2(_0513_));
 sg13g2_nand3_1 _5041_ (.B(_3367_),
    .C(_0514_),
    .A(_3118_),
    .Y(_0516_));
 sg13g2_nand4_1 _5042_ (.B(net2013),
    .C(_0115_),
    .A(net2515),
    .Y(_0517_),
    .D(net1998));
 sg13g2_a21oi_1 _5043_ (.A1(net2597),
    .A2(_0516_),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_a21oi_1 _5044_ (.A1(_0515_),
    .A2(_0518_),
    .Y(_0519_),
    .B1(_0512_));
 sg13g2_o21ai_1 _5045_ (.B1(net2297),
    .Y(_0520_),
    .A1(_0510_),
    .A2(_0519_));
 sg13g2_nand2_1 _5046_ (.Y(_0521_),
    .A(net2572),
    .B(net2209));
 sg13g2_a21oi_1 _5047_ (.A1(net2560),
    .A2(net2210),
    .Y(_0522_),
    .B1(net2539));
 sg13g2_nand4_1 _5048_ (.B(_0098_),
    .C(net2007),
    .A(_2724_),
    .Y(_0523_),
    .D(_0521_));
 sg13g2_nand2_1 _5049_ (.Y(_0524_),
    .A(net2530),
    .B(_0523_));
 sg13g2_nand4_1 _5050_ (.B(net2042),
    .C(_0088_),
    .A(net2572),
    .Y(_0525_),
    .D(_0494_));
 sg13g2_nand4_1 _5051_ (.B(net2042),
    .C(_0132_),
    .A(net2594),
    .Y(_0526_),
    .D(_0242_));
 sg13g2_nand3_1 _5052_ (.B(_0525_),
    .C(_0526_),
    .A(net2550),
    .Y(_0527_));
 sg13g2_nand4_1 _5053_ (.B(_3322_),
    .C(_0524_),
    .A(net2514),
    .Y(_0528_),
    .D(_0527_));
 sg13g2_o21ai_1 _5054_ (.B1(net2121),
    .Y(_0529_),
    .A1(net2069),
    .A2(_3166_));
 sg13g2_inv_1 _5055_ (.Y(_0530_),
    .A(_0529_));
 sg13g2_o21ai_1 _5056_ (.B1(net2117),
    .Y(_0531_),
    .A1(_3019_),
    .A2(_3166_));
 sg13g2_nand2_1 _5057_ (.Y(_0532_),
    .A(_3167_),
    .B(_3388_));
 sg13g2_a21oi_1 _5058_ (.A1(_0107_),
    .A2(_0531_),
    .Y(_0533_),
    .B1(net2548));
 sg13g2_nand2b_1 _5059_ (.Y(_0534_),
    .B(_0531_),
    .A_N(_3468_));
 sg13g2_nand3_1 _5060_ (.B(net2056),
    .C(_3232_),
    .A(net2180),
    .Y(_0535_));
 sg13g2_nand3_1 _5061_ (.B(net2008),
    .C(_0535_),
    .A(_3167_),
    .Y(_0536_));
 sg13g2_a22oi_1 _5062_ (.Y(_0537_),
    .B1(_0536_),
    .B2(net2449),
    .A2(_0534_),
    .A1(net2428));
 sg13g2_nor2_1 _5063_ (.A(net2513),
    .B(_0533_),
    .Y(_0538_));
 sg13g2_a21oi_1 _5064_ (.A1(_0537_),
    .A2(_0538_),
    .Y(_0539_),
    .B1(net2298));
 sg13g2_a21oi_2 _5065_ (.B1(net2382),
    .Y(_0540_),
    .A2(_0539_),
    .A1(_0528_));
 sg13g2_o21ai_1 _5066_ (.B1(net2448),
    .Y(_0541_),
    .A1(_3632_),
    .A2(_0532_));
 sg13g2_nand2_1 _5067_ (.Y(_0542_),
    .A(net2068),
    .B(_3619_));
 sg13g2_nand3_1 _5068_ (.B(_3018_),
    .C(_3161_),
    .A(net2269),
    .Y(_0543_));
 sg13g2_nor3_1 _5069_ (.A(net2575),
    .B(net2129),
    .C(_3380_),
    .Y(_0544_));
 sg13g2_a221oi_1 _5070_ (.B2(_0544_),
    .C1(net2331),
    .B1(_0543_),
    .A1(_3090_),
    .Y(_0545_),
    .A2(_0542_));
 sg13g2_and3_1 _5071_ (.X(_0546_),
    .A(net2123),
    .B(_2548_),
    .C(net2056));
 sg13g2_nand3_1 _5072_ (.B(_2548_),
    .C(net2056),
    .A(net2123),
    .Y(_0547_));
 sg13g2_nand2_1 _5073_ (.Y(_0548_),
    .A(net2253),
    .B(_3222_));
 sg13g2_o21ai_1 _5074_ (.B1(net2173),
    .Y(_0549_),
    .A1(net2088),
    .A2(_0471_));
 sg13g2_a21oi_1 _5075_ (.A1(net2575),
    .A2(_1899_),
    .Y(_0550_),
    .B1(net2337));
 sg13g2_and3_1 _5076_ (.X(_0551_),
    .A(_0547_),
    .B(_0549_),
    .C(_0550_));
 sg13g2_o21ai_1 _5077_ (.B1(_0541_),
    .Y(_0552_),
    .A1(_0545_),
    .A2(_0551_));
 sg13g2_nand3_1 _5078_ (.B(_0547_),
    .C(_0549_),
    .A(_3039_),
    .Y(_0553_));
 sg13g2_nor3_2 _5079_ (.A(net2263),
    .B(net2233),
    .C(net2223),
    .Y(_0554_));
 sg13g2_o21ai_1 _5080_ (.B1(net2122),
    .Y(_0555_),
    .A1(net2069),
    .A2(_0554_));
 sg13g2_nand4_1 _5081_ (.B(_3367_),
    .C(_0385_),
    .A(net2322),
    .Y(_0556_),
    .D(_0555_));
 sg13g2_a22oi_1 _5082_ (.Y(_0557_),
    .B1(_0553_),
    .B2(_0556_),
    .A2(_0516_),
    .A1(net2597));
 sg13g2_nor2_1 _5083_ (.A(_3301_),
    .B(_0557_),
    .Y(_0558_));
 sg13g2_nor2_1 _5084_ (.A(net2385),
    .B(net2039),
    .Y(_0559_));
 sg13g2_nand2_2 _5085_ (.Y(_0560_),
    .A(net2490),
    .B(net2432));
 sg13g2_nor2_2 _5086_ (.A(net2517),
    .B(net2449),
    .Y(_0561_));
 sg13g2_nand2_1 _5087_ (.Y(_0562_),
    .A(net2008),
    .B(_0339_));
 sg13g2_or3_1 _5088_ (.A(_3385_),
    .B(_0561_),
    .C(_0562_),
    .X(_0563_));
 sg13g2_a21oi_1 _5089_ (.A1(_0342_),
    .A2(_0561_),
    .Y(_0564_),
    .B1(_3311_));
 sg13g2_a221oi_1 _5090_ (.B2(_0564_),
    .C1(_0559_),
    .B1(_0563_),
    .A1(_0552_),
    .Y(_0565_),
    .A2(_0558_));
 sg13g2_a21oi_2 _5091_ (.B1(_0565_),
    .Y(_0566_),
    .A2(_0540_),
    .A1(_0520_));
 sg13g2_nor3_1 _5092_ (.A(net1978),
    .B(_0509_),
    .C(_0566_),
    .Y(_0567_));
 sg13g2_a21oi_1 _5093_ (.A1(_3035_),
    .A2(_0206_),
    .Y(_0568_),
    .B1(_3454_));
 sg13g2_o21ai_1 _5094_ (.B1(net2305),
    .Y(_0569_),
    .A1(_3176_),
    .A2(_0209_));
 sg13g2_nand3_1 _5095_ (.B(_0222_),
    .C(_0569_),
    .A(net2379),
    .Y(_0570_));
 sg13g2_nand2b_1 _5096_ (.Y(_0571_),
    .B(_3577_),
    .A_N(_3095_));
 sg13g2_a21oi_1 _5097_ (.A1(_0204_),
    .A2(_0571_),
    .Y(_0572_),
    .B1(net2314));
 sg13g2_nand3_1 _5098_ (.B(net2081),
    .C(net2220),
    .A(net2092),
    .Y(_0573_));
 sg13g2_nand3_1 _5099_ (.B(_3529_),
    .C(_0573_),
    .A(net2421),
    .Y(_0574_));
 sg13g2_nand2b_1 _5100_ (.Y(_0575_),
    .B(net2526),
    .A_N(_0218_));
 sg13g2_a21oi_1 _5101_ (.A1(_0574_),
    .A2(_0575_),
    .Y(_0576_),
    .B1(net2489));
 sg13g2_or4_1 _5102_ (.A(_0568_),
    .B(_0570_),
    .C(_0572_),
    .D(_0576_),
    .X(_0577_));
 sg13g2_o21ai_1 _5103_ (.B1(_0577_),
    .Y(_0578_),
    .A1(_0232_),
    .A2(_0235_));
 sg13g2_nand3_1 _5104_ (.B(net2195),
    .C(_3295_),
    .A(net2021),
    .Y(_0579_));
 sg13g2_nand3b_1 _5105_ (.B(_0579_),
    .C(net2300),
    .Y(_0580_),
    .A_N(_0198_));
 sg13g2_nor2_1 _5106_ (.A(net2509),
    .B(_3278_),
    .Y(_0581_));
 sg13g2_a21oi_1 _5107_ (.A1(net2509),
    .A2(_3272_),
    .Y(_0582_),
    .B1(_0581_));
 sg13g2_a21oi_1 _5108_ (.A1(net2381),
    .A2(_0582_),
    .Y(_0583_),
    .B1(_0580_));
 sg13g2_a21oi_1 _5109_ (.A1(net2294),
    .A2(_0578_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_nand3_1 _5110_ (.B(net2348),
    .C(_2691_),
    .A(net2115),
    .Y(_0585_));
 sg13g2_o21ai_1 _5111_ (.B1(net2163),
    .Y(_0586_),
    .A1(_3019_),
    .A2(net2065));
 sg13g2_and3_1 _5112_ (.X(_0587_),
    .A(_0474_),
    .B(_0585_),
    .C(_0586_));
 sg13g2_a21oi_1 _5113_ (.A1(net2601),
    .A2(_0168_),
    .Y(_0588_),
    .B1(net2532));
 sg13g2_nand2_1 _5114_ (.Y(_0589_),
    .A(net2276),
    .B(_2982_));
 sg13g2_a21oi_1 _5115_ (.A1(_2647_),
    .A2(_2982_),
    .Y(_0590_),
    .B1(_3467_));
 sg13g2_a221oi_1 _5116_ (.B2(_0586_),
    .C1(net2496),
    .B1(_0590_),
    .A1(_0587_),
    .Y(_0591_),
    .A2(_0588_));
 sg13g2_nand2_1 _5117_ (.Y(_0592_),
    .A(net2218),
    .B(net2073));
 sg13g2_o21ai_1 _5118_ (.B1(net2105),
    .Y(_0593_),
    .A1(_3274_),
    .A2(_0471_));
 sg13g2_a22oi_1 _5119_ (.Y(_0594_),
    .B1(_0159_),
    .B2(_0592_),
    .A2(_2836_),
    .A1(net2584));
 sg13g2_a21oi_1 _5120_ (.A1(_0593_),
    .A2(_0594_),
    .Y(_0595_),
    .B1(net2314));
 sg13g2_o21ai_1 _5121_ (.B1(net2153),
    .Y(_0596_),
    .A1(net2241),
    .A2(_2570_));
 sg13g2_a21oi_1 _5122_ (.A1(_0593_),
    .A2(_0596_),
    .Y(_0597_),
    .B1(_3454_));
 sg13g2_nand2b_1 _5123_ (.Y(_0598_),
    .B(net2076),
    .A_N(_2031_));
 sg13g2_o21ai_1 _5124_ (.B1(net2309),
    .Y(_0599_),
    .A1(net2146),
    .A2(_0598_));
 sg13g2_a21oi_1 _5125_ (.A1(_0376_),
    .A2(_0598_),
    .Y(_0600_),
    .B1(_0599_));
 sg13g2_nor4_1 _5126_ (.A(_0591_),
    .B(_0595_),
    .C(_0597_),
    .D(_0600_),
    .Y(_0601_));
 sg13g2_a221oi_1 _5127_ (.B2(net2341),
    .C1(_2416_),
    .B1(_0149_),
    .A1(_2647_),
    .Y(_0602_),
    .A2(net2215));
 sg13g2_a22oi_1 _5128_ (.Y(_0603_),
    .B1(_0602_),
    .B2(_0482_),
    .A2(_0587_),
    .A1(net2477));
 sg13g2_o21ai_1 _5129_ (.B1(net2152),
    .Y(_0604_),
    .A1(_3154_),
    .A2(_3425_));
 sg13g2_o21ai_1 _5130_ (.B1(_0604_),
    .Y(_0605_),
    .A1(net2463),
    .A2(_3354_));
 sg13g2_a22oi_1 _5131_ (.Y(_0606_),
    .B1(_3559_),
    .B2(_0150_),
    .A2(_3262_),
    .A1(net2523));
 sg13g2_o21ai_1 _5132_ (.B1(_0606_),
    .Y(_0607_),
    .A1(net2474),
    .A2(_0474_));
 sg13g2_o21ai_1 _5133_ (.B1(net2202),
    .Y(_0608_),
    .A1(_0605_),
    .A2(_0607_));
 sg13g2_o21ai_1 _5134_ (.B1(_0608_),
    .Y(_0609_),
    .A1(net2390),
    .A2(_0601_));
 sg13g2_a21o_1 _5135_ (.A2(_0603_),
    .A1(net2196),
    .B1(_0609_),
    .X(_0610_));
 sg13g2_a221oi_1 _5136_ (.B2(net2038),
    .C1(_0203_),
    .B1(_0610_),
    .A1(net1981),
    .Y(_0611_),
    .A2(_0584_));
 sg13g2_nor3_1 _5137_ (.A(net1976),
    .B(_0567_),
    .C(_0611_),
    .Y(_0612_));
 sg13g2_nor3_1 _5138_ (.A(_3505_),
    .B(_0443_),
    .C(_0612_),
    .Y(_0613_));
 sg13g2_o21ai_1 _5139_ (.B1(_1085_),
    .Y(_0614_),
    .A1(_0241_),
    .A2(_0613_));
 sg13g2_xnor2_1 _5140_ (.Y(_0615_),
    .A(_1459_),
    .B(_1525_));
 sg13g2_xnor2_1 _5141_ (.Y(_0616_),
    .A(_1470_),
    .B(_1525_));
 sg13g2_nand2_2 _5142_ (.Y(_0617_),
    .A(_3136_),
    .B(_3590_));
 sg13g2_nor2_2 _5143_ (.A(net2284),
    .B(_2982_),
    .Y(_0618_));
 sg13g2_a21oi_1 _5144_ (.A1(net2351),
    .A2(_0618_),
    .Y(_0619_),
    .B1(_3172_));
 sg13g2_o21ai_1 _5145_ (.B1(_3129_),
    .Y(_0620_),
    .A1(net2238),
    .A2(_2826_));
 sg13g2_a221oi_1 _5146_ (.B2(net2033),
    .C1(net2522),
    .B1(_0620_),
    .A1(net2040),
    .Y(_0621_),
    .A2(_0619_));
 sg13g2_nor4_2 _5147_ (.A(net2160),
    .B(net2248),
    .C(_2826_),
    .Y(_0622_),
    .D(_2948_));
 sg13g2_or2_1 _5148_ (.X(_0623_),
    .B(_0622_),
    .A(net2029));
 sg13g2_o21ai_1 _5149_ (.B1(net2570),
    .Y(_0624_),
    .A1(_0617_),
    .A2(_0623_));
 sg13g2_nand3_1 _5150_ (.B(net2282),
    .C(_3421_),
    .A(net2096),
    .Y(_0625_));
 sg13g2_nand2_1 _5151_ (.Y(_0626_),
    .A(_3150_),
    .B(_0625_));
 sg13g2_nand3_1 _5152_ (.B(_3150_),
    .C(_0625_),
    .A(net2581),
    .Y(_0627_));
 sg13g2_o21ai_1 _5153_ (.B1(_0627_),
    .Y(_0628_),
    .A1(net2582),
    .A2(_3158_));
 sg13g2_nor2_1 _5154_ (.A(net2542),
    .B(net2028),
    .Y(_0629_));
 sg13g2_a221oi_1 _5155_ (.B2(_0629_),
    .C1(net2199),
    .B1(_0628_),
    .A1(_0621_),
    .Y(_0630_),
    .A2(_0624_));
 sg13g2_nand2_1 _5156_ (.Y(_0631_),
    .A(net2345),
    .B(net2073));
 sg13g2_a21o_1 _5157_ (.A2(_0631_),
    .A1(net2041),
    .B1(_2482_),
    .X(_0632_));
 sg13g2_a21oi_1 _5158_ (.A1(_3192_),
    .A2(_0399_),
    .Y(_0633_),
    .B1(net2330));
 sg13g2_nand2_1 _5159_ (.Y(_0634_),
    .A(net2050),
    .B(_2863_));
 sg13g2_a221oi_1 _5160_ (.B2(net2306),
    .C1(_0633_),
    .B1(_0634_),
    .A1(net2319),
    .Y(_0635_),
    .A2(_0632_));
 sg13g2_mux2_2 _5161_ (.A0(net2244),
    .A1(net2235),
    .S(net2266),
    .X(_0637_));
 sg13g2_nor2_2 _5162_ (.A(net2124),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_nand2b_2 _5163_ (.Y(_0639_),
    .B(net2170),
    .A_N(_0637_));
 sg13g2_nand2_1 _5164_ (.Y(_0640_),
    .A(net2155),
    .B(net2082));
 sg13g2_nand2_2 _5165_ (.Y(_0641_),
    .A(_0639_),
    .B(net1995));
 sg13g2_nand3_1 _5166_ (.B(_0639_),
    .C(net1995),
    .A(_3192_),
    .Y(_0642_));
 sg13g2_nand3_1 _5167_ (.B(net2080),
    .C(net2222),
    .A(net2090),
    .Y(_0643_));
 sg13g2_a21oi_1 _5168_ (.A1(_2339_),
    .A2(_0643_),
    .Y(_0644_),
    .B1(_3411_));
 sg13g2_a221oi_1 _5169_ (.B2(_0642_),
    .C1(_0644_),
    .B1(_0426_),
    .A1(_0221_),
    .Y(_0645_),
    .A2(_0381_));
 sg13g2_a21o_1 _5170_ (.A2(_0645_),
    .A1(_0635_),
    .B1(net2388),
    .X(_0646_));
 sg13g2_nor3_2 _5171_ (.A(net2158),
    .B(net2353),
    .C(_3124_),
    .Y(_0648_));
 sg13g2_o21ai_1 _5172_ (.B1(net2561),
    .Y(_0649_),
    .A1(_3194_),
    .A2(_0648_));
 sg13g2_o21ai_1 _5173_ (.B1(net2582),
    .Y(_0650_),
    .A1(_2394_),
    .A2(_2713_));
 sg13g2_nand3_1 _5174_ (.B(_0649_),
    .C(_0650_),
    .A(_2636_),
    .Y(_0651_));
 sg13g2_and2_1 _5175_ (.A(_3459_),
    .B(_0651_),
    .X(_0652_));
 sg13g2_nor4_2 _5176_ (.A(net2295),
    .B(_0394_),
    .C(_0630_),
    .Y(_0653_),
    .D(_0652_));
 sg13g2_nor3_1 _5177_ (.A(net2563),
    .B(net2045),
    .C(_3054_),
    .Y(_0654_));
 sg13g2_o21ai_1 _5178_ (.B1(net2101),
    .Y(_0655_),
    .A1(net2244),
    .A2(net2080));
 sg13g2_a21oi_2 _5179_ (.B1(net2148),
    .Y(_0656_),
    .A2(net2081),
    .A1(net2241));
 sg13g2_nor3_1 _5180_ (.A(net2585),
    .B(net2045),
    .C(_0656_),
    .Y(_0657_));
 sg13g2_or3_1 _5181_ (.A(net2325),
    .B(_0654_),
    .C(_0657_),
    .X(_0659_));
 sg13g2_o21ai_1 _5182_ (.B1(net2318),
    .Y(_0660_),
    .A1(_3054_),
    .A2(_3056_));
 sg13g2_o21ai_1 _5183_ (.B1(_3410_),
    .Y(_0661_),
    .A1(_3044_),
    .A2(_0656_));
 sg13g2_nand3_1 _5184_ (.B(_0660_),
    .C(_0661_),
    .A(_0659_),
    .Y(_0662_));
 sg13g2_a22oi_1 _5185_ (.Y(_0663_),
    .B1(_3330_),
    .B2(net2421),
    .A2(_3259_),
    .A1(net2407));
 sg13g2_nand2_1 _5186_ (.Y(_0664_),
    .A(net2173),
    .B(_3022_));
 sg13g2_o21ai_1 _5187_ (.B1(net2439),
    .Y(_0665_),
    .A1(_3026_),
    .A2(_3093_));
 sg13g2_o21ai_1 _5188_ (.B1(_0665_),
    .Y(_0666_),
    .A1(_3293_),
    .A2(_0663_));
 sg13g2_a22oi_1 _5189_ (.Y(_0667_),
    .B1(_0666_),
    .B2(_0124_),
    .A2(_0662_),
    .A1(net2376));
 sg13g2_o21ai_1 _5190_ (.B1(net2089),
    .Y(_0668_),
    .A1(net2250),
    .A2(net2228));
 sg13g2_nand2_1 _5191_ (.Y(_0670_),
    .A(net2560),
    .B(_3088_));
 sg13g2_nand3_1 _5192_ (.B(_3088_),
    .C(_0668_),
    .A(net2440),
    .Y(_0671_));
 sg13g2_o21ai_1 _5193_ (.B1(net2439),
    .Y(_0672_),
    .A1(_1888_),
    .A2(_3104_));
 sg13g2_nand3_1 _5194_ (.B(_2734_),
    .C(_3086_),
    .A(net2421),
    .Y(_0673_));
 sg13g2_nand3_1 _5195_ (.B(_0672_),
    .C(_0673_),
    .A(_3108_),
    .Y(_0674_));
 sg13g2_a221oi_1 _5196_ (.B2(net2202),
    .C1(net2301),
    .B1(_0674_),
    .A1(_0415_),
    .Y(_0675_),
    .A2(_0671_));
 sg13g2_a221oi_1 _5197_ (.B2(_0675_),
    .C1(net2035),
    .B1(_0667_),
    .A1(_0646_),
    .Y(_0676_),
    .A2(_0653_));
 sg13g2_nand3_1 _5198_ (.B(_3265_),
    .C(_3296_),
    .A(net2462),
    .Y(_0677_));
 sg13g2_nand2_1 _5199_ (.Y(_0678_),
    .A(net2294),
    .B(_0677_));
 sg13g2_nand3_1 _5200_ (.B(_3091_),
    .C(_3478_),
    .A(net2338),
    .Y(_0679_));
 sg13g2_o21ai_1 _5201_ (.B1(net2442),
    .Y(_0681_),
    .A1(_3054_),
    .A2(_3238_));
 sg13g2_o21ai_1 _5202_ (.B1(net2305),
    .Y(_0682_),
    .A1(_3054_),
    .A2(_3238_));
 sg13g2_o21ai_1 _5203_ (.B1(net2328),
    .Y(_0683_),
    .A1(net2020),
    .A2(_0434_));
 sg13g2_mux2_2 _5204_ (.A0(_3245_),
    .A1(_0169_),
    .S(net2106),
    .X(_0684_));
 sg13g2_nand2_1 _5205_ (.Y(_0685_),
    .A(net2564),
    .B(_0684_));
 sg13g2_nand2b_1 _5206_ (.Y(_0686_),
    .B(_0685_),
    .A_N(_0190_));
 sg13g2_nand2_2 _5207_ (.Y(_0687_),
    .A(_2816_),
    .B(net2055));
 sg13g2_nand2_2 _5208_ (.Y(_0688_),
    .A(_3297_),
    .B(_0687_));
 sg13g2_nand3_1 _5209_ (.B(_0681_),
    .C(_0688_),
    .A(_3240_),
    .Y(_0689_));
 sg13g2_nand3_1 _5210_ (.B(_0679_),
    .C(_0683_),
    .A(net2391),
    .Y(_0690_));
 sg13g2_a221oi_1 _5211_ (.B2(net2509),
    .C1(_0690_),
    .B1(_0689_),
    .A1(net2319),
    .Y(_0692_),
    .A2(_0686_));
 sg13g2_nor2_1 _5212_ (.A(net2564),
    .B(_3272_),
    .Y(_0693_));
 sg13g2_nand2_1 _5213_ (.Y(_0694_),
    .A(_3255_),
    .B(_3277_));
 sg13g2_a21oi_1 _5214_ (.A1(_3255_),
    .A2(_3277_),
    .Y(_0695_),
    .B1(net2587));
 sg13g2_o21ai_1 _5215_ (.B1(net2338),
    .Y(_0696_),
    .A1(_0693_),
    .A2(_0695_));
 sg13g2_o21ai_1 _5216_ (.B1(net2378),
    .Y(_0697_),
    .A1(net2508),
    .A2(_3272_));
 sg13g2_a21oi_1 _5217_ (.A1(net2332),
    .A2(_3278_),
    .Y(_0698_),
    .B1(_0697_));
 sg13g2_nand3_1 _5218_ (.B(_0696_),
    .C(_0698_),
    .A(_0425_),
    .Y(_0699_));
 sg13g2_nand3b_1 _5219_ (.B(_0699_),
    .C(net2300),
    .Y(_0700_),
    .A_N(_0692_));
 sg13g2_a21oi_1 _5220_ (.A1(_0678_),
    .A2(_0700_),
    .Y(_0701_),
    .B1(net2037));
 sg13g2_nor3_2 _5221_ (.A(net1979),
    .B(_0676_),
    .C(_0701_),
    .Y(_0703_));
 sg13g2_o21ai_1 _5222_ (.B1(_0365_),
    .Y(_0704_),
    .A1(net2404),
    .A2(_3457_));
 sg13g2_a22oi_1 _5223_ (.Y(_0705_),
    .B1(_0561_),
    .B2(_0322_),
    .A2(_0370_),
    .A1(_3048_));
 sg13g2_nor2_1 _5224_ (.A(net2400),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_nand3_1 _5225_ (.B(_3456_),
    .C(net2000),
    .A(_3441_),
    .Y(_0707_));
 sg13g2_a21oi_1 _5226_ (.A1(net2197),
    .A2(_0704_),
    .Y(_0708_),
    .B1(_0706_));
 sg13g2_a21oi_1 _5227_ (.A1(_3459_),
    .A2(_0707_),
    .Y(_0709_),
    .B1(_0362_));
 sg13g2_nand4_1 _5228_ (.B(net2019),
    .C(net2010),
    .A(_3367_),
    .Y(_0710_),
    .D(_0339_));
 sg13g2_nand2_1 _5229_ (.Y(_0711_),
    .A(net2556),
    .B(_0710_));
 sg13g2_a221oi_1 _5230_ (.B2(net2436),
    .C1(_0344_),
    .B1(_0367_),
    .A1(net2481),
    .Y(_0712_),
    .A2(_0366_));
 sg13g2_a21o_1 _5231_ (.A2(_0712_),
    .A1(_0711_),
    .B1(net2384),
    .X(_0714_));
 sg13g2_o21ai_1 _5232_ (.B1(net2327),
    .Y(_0715_),
    .A1(_3407_),
    .A2(_0354_));
 sg13g2_a221oi_1 _5233_ (.B2(_0715_),
    .C1(net2397),
    .B1(_0353_),
    .A1(_0349_),
    .Y(_0716_),
    .A2(_0351_));
 sg13g2_nor2_1 _5234_ (.A(_0357_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_a221oi_1 _5235_ (.B2(_0717_),
    .C1(net2036),
    .B1(_0714_),
    .A1(_0708_),
    .Y(_0718_),
    .A2(_0709_));
 sg13g2_a22oi_1 _5236_ (.Y(_0719_),
    .B1(_0623_),
    .B2(net2411),
    .A2(_0617_),
    .A1(net2531));
 sg13g2_nand3_1 _5237_ (.B(net2219),
    .C(_3320_),
    .A(net2112),
    .Y(_0720_));
 sg13g2_nand4_1 _5238_ (.B(_3138_),
    .C(_3590_),
    .A(_3136_),
    .Y(_0721_),
    .D(_0720_));
 sg13g2_nand2_1 _5239_ (.Y(_0722_),
    .A(_3129_),
    .B(_0174_));
 sg13g2_a21oi_1 _5240_ (.A1(_3606_),
    .A2(_0722_),
    .Y(_0723_),
    .B1(net2513));
 sg13g2_nand2_2 _5241_ (.Y(_0725_),
    .A(net2113),
    .B(_0618_));
 sg13g2_nand4_1 _5242_ (.B(_3575_),
    .C(_0282_),
    .A(_3132_),
    .Y(_0726_),
    .D(_0725_));
 sg13g2_a22oi_1 _5243_ (.Y(_0727_),
    .B1(_0726_),
    .B2(net2443),
    .A2(_0721_),
    .A1(net2425));
 sg13g2_nand3_1 _5244_ (.B(_0723_),
    .C(_0727_),
    .A(_0719_),
    .Y(_0728_));
 sg13g2_a21oi_2 _5245_ (.B1(net2259),
    .Y(_0729_),
    .A2(net2236),
    .A1(net2373));
 sg13g2_nand3_1 _5246_ (.B(net2241),
    .C(_0729_),
    .A(net2099),
    .Y(_0730_));
 sg13g2_o21ai_1 _5247_ (.B1(net2168),
    .Y(_0731_),
    .A1(net2085),
    .A2(_3022_));
 sg13g2_a21oi_1 _5248_ (.A1(net2084),
    .A2(_3023_),
    .Y(_0732_),
    .B1(net2124));
 sg13g2_nand3_1 _5249_ (.B(_0730_),
    .C(net1994),
    .A(net2005),
    .Y(_0733_));
 sg13g2_nand2_1 _5250_ (.Y(_0734_),
    .A(net2426),
    .B(_0733_));
 sg13g2_nor2_2 _5251_ (.A(net2256),
    .B(net2241),
    .Y(_0736_));
 sg13g2_nand2_1 _5252_ (.Y(_0737_),
    .A(net2286),
    .B(net2244));
 sg13g2_nand2_2 _5253_ (.Y(_0738_),
    .A(net2182),
    .B(net2052));
 sg13g2_nor2_1 _5254_ (.A(_2251_),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_nor3_2 _5255_ (.A(net2158),
    .B(net2215),
    .C(_3235_),
    .Y(_0740_));
 sg13g2_o21ai_1 _5256_ (.B1(net2445),
    .Y(_0741_),
    .A1(_0739_),
    .A2(_0740_));
 sg13g2_a21oi_2 _5257_ (.B1(_3078_),
    .Y(_0742_),
    .A2(net2208),
    .A1(net2284));
 sg13g2_nand2_1 _5258_ (.Y(_0743_),
    .A(net2118),
    .B(_0742_));
 sg13g2_o21ai_1 _5259_ (.B1(net2119),
    .Y(_0744_),
    .A1(_1712_),
    .A2(_0742_));
 sg13g2_nand3_1 _5260_ (.B(_0282_),
    .C(_0744_),
    .A(net2512),
    .Y(_0745_));
 sg13g2_nand2_1 _5261_ (.Y(_0747_),
    .A(net2331),
    .B(_0745_));
 sg13g2_nand3_1 _5262_ (.B(_0741_),
    .C(_0747_),
    .A(_0734_),
    .Y(_0748_));
 sg13g2_nand3_1 _5263_ (.B(_0728_),
    .C(_0748_),
    .A(net2387),
    .Y(_0749_));
 sg13g2_o21ai_1 _5264_ (.B1(net2171),
    .Y(_0750_),
    .A1(net2086),
    .A2(_3147_));
 sg13g2_a21oi_1 _5265_ (.A1(net2084),
    .A2(_3148_),
    .Y(_0751_),
    .B1(net2123));
 sg13g2_nand3_1 _5266_ (.B(_0255_),
    .C(net1993),
    .A(net2016),
    .Y(_0752_));
 sg13g2_nand2_1 _5267_ (.Y(_0753_),
    .A(net2550),
    .B(_0752_));
 sg13g2_nor2_2 _5268_ (.A(_3380_),
    .B(net2001),
    .Y(_0754_));
 sg13g2_nor2_2 _5269_ (.A(net2064),
    .B(_3397_),
    .Y(_0755_));
 sg13g2_nor2_1 _5270_ (.A(_3028_),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_o21ai_1 _5271_ (.B1(net2343),
    .Y(_0758_),
    .A1(_0754_),
    .A2(_0756_));
 sg13g2_o21ai_1 _5272_ (.B1(_3606_),
    .Y(_0759_),
    .A1(net2069),
    .A2(_0258_));
 sg13g2_a22oi_1 _5273_ (.Y(_0760_),
    .B1(_0638_),
    .B2(net2479),
    .A2(_3241_),
    .A1(net2082));
 sg13g2_nand4_1 _5274_ (.B(_0758_),
    .C(_0759_),
    .A(_0753_),
    .Y(_0761_),
    .D(_0760_));
 sg13g2_a22oi_1 _5275_ (.Y(_0762_),
    .B1(_3352_),
    .B2(net2084),
    .A2(_3076_),
    .A1(_3033_));
 sg13g2_a22oi_1 _5276_ (.Y(_0763_),
    .B1(_0762_),
    .B2(net2444),
    .A2(_0249_),
    .A1(net2427));
 sg13g2_nor2_1 _5277_ (.A(_3220_),
    .B(_0738_),
    .Y(_0764_));
 sg13g2_nor2_1 _5278_ (.A(net2594),
    .B(_3204_),
    .Y(_0765_));
 sg13g2_o21ai_1 _5279_ (.B1(net2434),
    .Y(_0766_),
    .A1(_0764_),
    .A2(_0765_));
 sg13g2_a21oi_1 _5280_ (.A1(_0763_),
    .A2(_0766_),
    .Y(_0767_),
    .B1(net2193));
 sg13g2_a221oi_1 _5281_ (.B2(net2207),
    .C1(_0767_),
    .B1(_0761_),
    .A1(_3459_),
    .Y(_0769_),
    .A2(_0740_));
 sg13g2_a21oi_2 _5282_ (.B1(net1983),
    .Y(_0770_),
    .A2(_0769_),
    .A1(_0749_));
 sg13g2_nand2_1 _5283_ (.Y(_0771_),
    .A(_3132_),
    .B(_3484_));
 sg13g2_nor3_2 _5284_ (.A(net2270),
    .B(net2359),
    .C(net2224),
    .Y(_0772_));
 sg13g2_or2_2 _5285_ (.X(_0773_),
    .B(_0772_),
    .A(net2179));
 sg13g2_nor2_2 _5286_ (.A(net2002),
    .B(_0772_),
    .Y(_0774_));
 sg13g2_or3_2 _5287_ (.A(net2184),
    .B(net2058),
    .C(_0772_),
    .X(_0775_));
 sg13g2_nand2_2 _5288_ (.Y(_0776_),
    .A(net2515),
    .B(_0775_));
 sg13g2_a221oi_1 _5289_ (.B2(net2574),
    .C1(_0776_),
    .B1(_0771_),
    .A1(_3232_),
    .Y(_0777_),
    .A2(_3353_));
 sg13g2_a21oi_1 _5290_ (.A1(_3416_),
    .A2(_0307_),
    .Y(_0778_),
    .B1(net2597));
 sg13g2_o21ai_1 _5291_ (.B1(net2068),
    .Y(_0780_),
    .A1(net2084),
    .A2(net2229));
 sg13g2_a21oi_1 _5292_ (.A1(net2270),
    .A2(net2209),
    .Y(_0781_),
    .B1(net2232));
 sg13g2_a221oi_1 _5293_ (.B2(_3024_),
    .C1(net2515),
    .B1(_0781_),
    .A1(net2033),
    .Y(_0782_),
    .A2(_0780_));
 sg13g2_nor2_1 _5294_ (.A(net2149),
    .B(_3517_),
    .Y(_0783_));
 sg13g2_nand3_1 _5295_ (.B(net2126),
    .C(_3518_),
    .A(net2574),
    .Y(_0784_));
 sg13g2_o21ai_1 _5296_ (.B1(_0782_),
    .Y(_0785_),
    .A1(net2058),
    .A2(_0784_));
 sg13g2_o21ai_1 _5297_ (.B1(net2554),
    .Y(_0786_),
    .A1(_0778_),
    .A2(_0785_));
 sg13g2_nand2_1 _5298_ (.Y(_0787_),
    .A(net1996),
    .B(_0750_));
 sg13g2_nand3_1 _5299_ (.B(net1995),
    .C(net1993),
    .A(net1996),
    .Y(_0788_));
 sg13g2_nand2_2 _5300_ (.Y(_0789_),
    .A(net2096),
    .B(_3604_));
 sg13g2_o21ai_1 _5301_ (.B1(net2097),
    .Y(_0791_),
    .A1(net2069),
    .A2(_3604_));
 sg13g2_nand3_1 _5302_ (.B(_0307_),
    .C(_0791_),
    .A(_3416_),
    .Y(_0792_));
 sg13g2_o21ai_1 _5303_ (.B1(net2385),
    .Y(_0793_),
    .A1(_2826_),
    .A2(_3062_));
 sg13g2_a221oi_1 _5304_ (.B2(net2340),
    .C1(_0793_),
    .B1(_0792_),
    .A1(net2322),
    .Y(_0794_),
    .A2(_0788_));
 sg13g2_o21ai_1 _5305_ (.B1(_0794_),
    .Y(_0795_),
    .A1(_0777_),
    .A2(_0786_));
 sg13g2_o21ai_1 _5306_ (.B1(net2322),
    .Y(_0796_),
    .A1(_0324_),
    .A2(_0771_));
 sg13g2_nand2_1 _5307_ (.Y(_0797_),
    .A(net2012),
    .B(net2010));
 sg13g2_a22oi_1 _5308_ (.Y(_0798_),
    .B1(_0797_),
    .B2(net2305),
    .A2(_0707_),
    .A1(net2335));
 sg13g2_o21ai_1 _5309_ (.B1(net2040),
    .Y(_0799_),
    .A1(_2691_),
    .A2(_3402_));
 sg13g2_a21o_1 _5310_ (.A2(_0799_),
    .A1(_0326_),
    .B1(net2327),
    .X(_0800_));
 sg13g2_nand4_1 _5311_ (.B(_0796_),
    .C(_0798_),
    .A(_0332_),
    .Y(_0802_),
    .D(_0800_));
 sg13g2_and3_1 _5312_ (.X(_0803_),
    .A(_3300_),
    .B(_0795_),
    .C(_0802_));
 sg13g2_nor4_2 _5313_ (.A(net1977),
    .B(_0718_),
    .C(_0770_),
    .Y(_0804_),
    .D(_0803_));
 sg13g2_nor3_1 _5314_ (.A(_3308_),
    .B(_0703_),
    .C(_0804_),
    .Y(_0805_));
 sg13g2_nor2_1 _5315_ (.A(_3493_),
    .B(net2001),
    .Y(_0806_));
 sg13g2_or3_2 _5316_ (.A(net2182),
    .B(net2059),
    .C(_3493_),
    .X(_0807_));
 sg13g2_nand3_1 _5317_ (.B(net2351),
    .C(net2077),
    .A(net2173),
    .Y(_0808_));
 sg13g2_a21oi_1 _5318_ (.A1(_0807_),
    .A2(_0808_),
    .Y(_0809_),
    .B1(net2436));
 sg13g2_a21oi_1 _5319_ (.A1(_3118_),
    .A2(_0514_),
    .Y(_0810_),
    .B1(net2468));
 sg13g2_nand2_1 _5320_ (.Y(_0811_),
    .A(net2498),
    .B(_3416_));
 sg13g2_o21ai_1 _5321_ (.B1(net2414),
    .Y(_0813_),
    .A1(_3436_),
    .A2(_3473_));
 sg13g2_nand3_1 _5322_ (.B(_3101_),
    .C(net2055),
    .A(net2182),
    .Y(_0814_));
 sg13g2_nand3_1 _5323_ (.B(net2057),
    .C(_3414_),
    .A(net2129),
    .Y(_0815_));
 sg13g2_a21oi_1 _5324_ (.A1(_0814_),
    .A2(_0815_),
    .Y(_0816_),
    .B1(net2418));
 sg13g2_nor4_1 _5325_ (.A(_0809_),
    .B(_0810_),
    .C(_0811_),
    .D(_0816_),
    .Y(_0817_));
 sg13g2_o21ai_1 _5326_ (.B1(net2181),
    .Y(_0818_),
    .A1(net2085),
    .A2(net2055));
 sg13g2_o21ai_1 _5327_ (.B1(_0818_),
    .Y(_0819_),
    .A1(net2058),
    .A2(_0271_));
 sg13g2_nor2_2 _5328_ (.A(net2575),
    .B(net2230),
    .Y(_0820_));
 sg13g2_a22oi_1 _5329_ (.Y(_0821_),
    .B1(_0820_),
    .B2(net2270),
    .A2(_0543_),
    .A1(net2180));
 sg13g2_a21oi_1 _5330_ (.A1(_0807_),
    .A2(_0821_),
    .Y(_0822_),
    .B1(net2554));
 sg13g2_nor2_2 _5331_ (.A(_0157_),
    .B(net2002),
    .Y(_0824_));
 sg13g2_nand3_1 _5332_ (.B(net2057),
    .C(_0158_),
    .A(net2129),
    .Y(_0825_));
 sg13g2_o21ai_1 _5333_ (.B1(_0825_),
    .Y(_0826_),
    .A1(_2306_),
    .A2(_3631_));
 sg13g2_a221oi_1 _5334_ (.B2(net2448),
    .C1(_0822_),
    .B1(_0826_),
    .A1(net2428),
    .Y(_0827_),
    .A2(_0819_));
 sg13g2_nand2_1 _5335_ (.Y(_0828_),
    .A(net2515),
    .B(_0827_));
 sg13g2_a21oi_1 _5336_ (.A1(_0813_),
    .A2(_0817_),
    .Y(_0829_),
    .B1(net2399));
 sg13g2_nand2_1 _5337_ (.Y(_0830_),
    .A(_0828_),
    .B(_0829_));
 sg13g2_o21ai_1 _5338_ (.B1(net2530),
    .Y(_0831_),
    .A1(_3253_),
    .A2(_3338_));
 sg13g2_a21oi_2 _5339_ (.B1(net2572),
    .Y(_0832_),
    .A2(_0242_),
    .A1(net2018));
 sg13g2_nor4_2 _5340_ (.A(net2571),
    .B(net2123),
    .C(_0138_),
    .Y(_0833_),
    .D(_0139_));
 sg13g2_nand2b_1 _5341_ (.Y(_0835_),
    .B(net2551),
    .A_N(_0833_));
 sg13g2_o21ai_1 _5342_ (.B1(_0831_),
    .Y(_0836_),
    .A1(_0832_),
    .A2(_0835_));
 sg13g2_nand3_1 _5343_ (.B(_0098_),
    .C(_0529_),
    .A(net2030),
    .Y(_0837_));
 sg13g2_nor2_2 _5344_ (.A(net2123),
    .B(_0138_),
    .Y(_0838_));
 sg13g2_nand2b_1 _5345_ (.Y(_0839_),
    .B(net2170),
    .A_N(_0138_));
 sg13g2_o21ai_1 _5346_ (.B1(net2446),
    .Y(_0840_),
    .A1(_0740_),
    .A2(_0838_));
 sg13g2_nand2_1 _5347_ (.Y(_0841_),
    .A(net2030),
    .B(_0132_));
 sg13g2_a22oi_1 _5348_ (.Y(_0842_),
    .B1(_0841_),
    .B2(net2412),
    .A2(_0837_),
    .A1(net2478));
 sg13g2_nand3_1 _5349_ (.B(_0840_),
    .C(_0842_),
    .A(_0836_),
    .Y(_0843_));
 sg13g2_nand2_2 _5350_ (.Y(_0844_),
    .A(_3343_),
    .B(_3398_));
 sg13g2_a22oi_1 _5351_ (.Y(_0846_),
    .B1(_0844_),
    .B2(net2040),
    .A2(_0530_),
    .A1(net2594));
 sg13g2_nand2_2 _5352_ (.Y(_0847_),
    .A(net2182),
    .B(_0311_));
 sg13g2_nand2_1 _5353_ (.Y(_0848_),
    .A(_0529_),
    .B(_0847_));
 sg13g2_o21ai_1 _5354_ (.B1(net2180),
    .Y(_0849_),
    .A1(_2559_),
    .A2(_0311_));
 sg13g2_a21oi_1 _5355_ (.A1(_0529_),
    .A2(_0849_),
    .Y(_0850_),
    .B1(net2436));
 sg13g2_nand3_1 _5356_ (.B(net1995),
    .C(_0847_),
    .A(_0529_),
    .Y(_0851_));
 sg13g2_a21oi_1 _5357_ (.A1(net2344),
    .A2(_0851_),
    .Y(_0852_),
    .B1(_0850_));
 sg13g2_o21ai_1 _5358_ (.B1(_0852_),
    .Y(_0853_),
    .A1(net2550),
    .A2(_0846_));
 sg13g2_a221oi_1 _5359_ (.B2(net2197),
    .C1(net2298),
    .B1(_0853_),
    .A1(net2207),
    .Y(_0854_),
    .A2(_0843_));
 sg13g2_a22oi_1 _5360_ (.Y(_0855_),
    .B1(_0710_),
    .B2(net2535),
    .A2(_0562_),
    .A1(net2481));
 sg13g2_o21ai_1 _5361_ (.B1(_0514_),
    .Y(_0857_),
    .A1(_3231_),
    .A2(_3631_));
 sg13g2_nand2_1 _5362_ (.Y(_0858_),
    .A(net2554),
    .B(_0857_));
 sg13g2_a221oi_1 _5363_ (.B2(_0518_),
    .C1(net2385),
    .B1(_0858_),
    .A1(_0512_),
    .Y(_0859_),
    .A2(_0855_));
 sg13g2_nor2_1 _5364_ (.A(_0366_),
    .B(_0562_),
    .Y(_0860_));
 sg13g2_nor2_1 _5365_ (.A(net2316),
    .B(_0710_),
    .Y(_0861_));
 sg13g2_a21oi_1 _5366_ (.A1(net2315),
    .A2(_0860_),
    .Y(_0862_),
    .B1(_0861_));
 sg13g2_a21oi_1 _5367_ (.A1(net2385),
    .A2(_0862_),
    .Y(_0863_),
    .B1(_0859_));
 sg13g2_a221oi_1 _5368_ (.B2(net2297),
    .C1(net2039),
    .B1(_0863_),
    .A1(_0830_),
    .Y(_0864_),
    .A2(_0854_));
 sg13g2_nand4_1 _5369_ (.B(net2046),
    .C(net2044),
    .A(net2485),
    .Y(_0865_),
    .D(_3546_));
 sg13g2_nor2_2 _5370_ (.A(net2268),
    .B(net2351),
    .Y(_0866_));
 sg13g2_nor2_2 _5371_ (.A(net2264),
    .B(_0224_),
    .Y(_0868_));
 sg13g2_a21oi_2 _5372_ (.B1(net2141),
    .Y(_0869_),
    .A2(_3542_),
    .A1(_3146_));
 sg13g2_nor3_1 _5373_ (.A(_0450_),
    .B(_0868_),
    .C(_0869_),
    .Y(_0870_));
 sg13g2_o21ai_1 _5374_ (.B1(net2408),
    .Y(_0871_),
    .A1(_3544_),
    .A2(_0450_));
 sg13g2_o21ai_1 _5375_ (.B1(_0871_),
    .Y(_0872_),
    .A1(net2522),
    .A2(_0870_));
 sg13g2_a21o_1 _5376_ (.A2(_0865_),
    .A1(_1371_),
    .B1(_0872_),
    .X(_0873_));
 sg13g2_a21oi_1 _5377_ (.A1(net2220),
    .A2(_3169_),
    .Y(_0874_),
    .B1(_3607_));
 sg13g2_nor2_1 _5378_ (.A(_2086_),
    .B(_3605_),
    .Y(_0875_));
 sg13g2_a21oi_1 _5379_ (.A1(_3160_),
    .A2(net2022),
    .Y(_0876_),
    .B1(net2337));
 sg13g2_a22oi_1 _5380_ (.Y(_0877_),
    .B1(_0876_),
    .B2(_2339_),
    .A2(_0875_),
    .A1(net2334));
 sg13g2_o21ai_1 _5381_ (.B1(_0873_),
    .Y(_0879_),
    .A1(_0874_),
    .A2(_0877_));
 sg13g2_o21ai_1 _5382_ (.B1(net2580),
    .Y(_0880_),
    .A1(net2091),
    .A2(net2075));
 sg13g2_a21oi_1 _5383_ (.A1(_0670_),
    .A2(_0880_),
    .Y(_0881_),
    .B1(_0445_));
 sg13g2_o21ai_1 _5384_ (.B1(_3580_),
    .Y(_0882_),
    .A1(net2540),
    .A2(_0881_));
 sg13g2_o21ai_1 _5385_ (.B1(net2440),
    .Y(_0883_),
    .A1(net2034),
    .A2(_0445_));
 sg13g2_a221oi_1 _5386_ (.B2(net2366),
    .C1(net2137),
    .B1(net2356),
    .A1(net2273),
    .Y(_0884_),
    .A2(net2358));
 sg13g2_o21ai_1 _5387_ (.B1(net2407),
    .Y(_0885_),
    .A1(_0464_),
    .A2(_0884_));
 sg13g2_a21oi_2 _5388_ (.B1(net2092),
    .Y(_0886_),
    .A2(net2075),
    .A1(net2240));
 sg13g2_o21ai_1 _5389_ (.B1(net2146),
    .Y(_0887_),
    .A1(net2244),
    .A2(_2912_));
 sg13g2_o21ai_1 _5390_ (.B1(net2422),
    .Y(_0888_),
    .A1(_3587_),
    .A2(_0886_));
 sg13g2_a21oi_2 _5391_ (.B1(net2090),
    .Y(_0890_),
    .A2(net2345),
    .A1(net2250));
 sg13g2_a221oi_1 _5392_ (.B2(net2470),
    .C1(net2502),
    .B1(_0890_),
    .A1(_3160_),
    .Y(_0891_),
    .A2(_3606_));
 sg13g2_nand4_1 _5393_ (.B(_0885_),
    .C(_0888_),
    .A(_0883_),
    .Y(_0892_),
    .D(_0891_));
 sg13g2_and2_1 _5394_ (.A(net2388),
    .B(_0892_),
    .X(_0893_));
 sg13g2_a21oi_1 _5395_ (.A1(_0882_),
    .A2(_0893_),
    .Y(_0894_),
    .B1(net2295));
 sg13g2_o21ai_1 _5396_ (.B1(_0894_),
    .Y(_0895_),
    .A1(net2390),
    .A2(_0879_));
 sg13g2_nand3_1 _5397_ (.B(net2006),
    .C(net1994),
    .A(_3575_),
    .Y(_0896_));
 sg13g2_nor3_2 _5398_ (.A(net2265),
    .B(net2356),
    .C(net2233),
    .Y(_0897_));
 sg13g2_nand2_2 _5399_ (.Y(_0898_),
    .A(net2120),
    .B(_0897_));
 sg13g2_o21ai_1 _5400_ (.B1(net2120),
    .Y(_0899_),
    .A1(net2054),
    .A2(_0897_));
 sg13g2_nand2_1 _5401_ (.Y(_0901_),
    .A(_0282_),
    .B(_0899_));
 sg13g2_a221oi_1 _5402_ (.B2(net2266),
    .C1(net2124),
    .B1(net2224),
    .A1(net2084),
    .Y(_0902_),
    .A2(net2076));
 sg13g2_or2_1 _5403_ (.X(_0903_),
    .B(_0902_),
    .A(_0740_));
 sg13g2_o21ai_1 _5404_ (.B1(net2529),
    .Y(_0904_),
    .A1(_0833_),
    .A2(_0903_));
 sg13g2_a221oi_1 _5405_ (.B2(net2445),
    .C1(net2512),
    .B1(_0901_),
    .A1(net2426),
    .Y(_0905_),
    .A2(_0896_));
 sg13g2_xnor2_1 _5406_ (.Y(_0906_),
    .A(net2118),
    .B(_3340_));
 sg13g2_a21oi_1 _5407_ (.A1(_3612_),
    .A2(_0906_),
    .Y(_0907_),
    .B1(net2418));
 sg13g2_nor2_1 _5408_ (.A(_0618_),
    .B(_0897_),
    .Y(_0908_));
 sg13g2_nand2_1 _5409_ (.Y(_0909_),
    .A(net2146),
    .B(_3513_));
 sg13g2_a221oi_1 _5410_ (.B2(net2113),
    .C1(net2404),
    .B1(_0908_),
    .A1(_3125_),
    .Y(_0910_),
    .A2(_3513_));
 sg13g2_o21ai_1 _5411_ (.B1(net2118),
    .Y(_0912_),
    .A1(net2064),
    .A2(_3350_));
 sg13g2_nand3_1 _5412_ (.B(_2207_),
    .C(_3122_),
    .A(net2262),
    .Y(_0913_));
 sg13g2_nand2_1 _5413_ (.Y(_0914_),
    .A(_0481_),
    .B(_0913_));
 sg13g2_a21oi_1 _5414_ (.A1(_0912_),
    .A2(_0914_),
    .Y(_0915_),
    .B1(net2434));
 sg13g2_nor3_2 _5415_ (.A(_0907_),
    .B(_0910_),
    .C(_0915_),
    .Y(_0916_));
 sg13g2_a21oi_1 _5416_ (.A1(net2478),
    .A2(_0901_),
    .Y(_0917_),
    .B1(net2494));
 sg13g2_a221oi_1 _5417_ (.B2(_0917_),
    .C1(net2396),
    .B1(_0916_),
    .A1(_0904_),
    .Y(_0918_),
    .A2(_0905_));
 sg13g2_o21ai_1 _5418_ (.B1(net2176),
    .Y(_0919_),
    .A1(net2372),
    .A2(_3102_));
 sg13g2_a221oi_1 _5419_ (.B2(net2061),
    .C1(net2110),
    .B1(net2062),
    .A1(net2363),
    .Y(_0920_),
    .A2(_3101_));
 sg13g2_or2_1 _5420_ (.X(_0921_),
    .B(_0920_),
    .A(_3170_));
 sg13g2_nand4_1 _5421_ (.B(_3167_),
    .C(_3595_),
    .A(net2048),
    .Y(_0923_),
    .D(_3596_));
 sg13g2_a22oi_1 _5422_ (.Y(_0924_),
    .B1(_0923_),
    .B2(net2443),
    .A2(_0921_),
    .A1(net2476));
 sg13g2_a21oi_1 _5423_ (.A1(_0476_),
    .A2(_0924_),
    .Y(_0925_),
    .B1(net2200));
 sg13g2_nand3_1 _5424_ (.B(_3569_),
    .C(_0912_),
    .A(net2012),
    .Y(_0926_));
 sg13g2_nand4_1 _5425_ (.B(_3550_),
    .C(_3551_),
    .A(net2026),
    .Y(_0927_),
    .D(net1997));
 sg13g2_a22oi_1 _5426_ (.Y(_0928_),
    .B1(_0927_),
    .B2(net2207),
    .A2(_0926_),
    .A1(net2197));
 sg13g2_a221oi_1 _5427_ (.B2(net2570),
    .C1(_3135_),
    .B1(_0452_),
    .A1(_3085_),
    .Y(_0929_),
    .A2(net2055));
 sg13g2_a21oi_1 _5428_ (.A1(_0912_),
    .A2(_0929_),
    .Y(_0930_),
    .B1(_3460_));
 sg13g2_nand3_1 _5429_ (.B(net2246),
    .C(_3079_),
    .A(net2284),
    .Y(_0931_));
 sg13g2_a21o_1 _5430_ (.A2(_0931_),
    .A1(_3148_),
    .B1(net2160),
    .X(_0932_));
 sg13g2_nand2b_1 _5431_ (.Y(_0934_),
    .B(_0932_),
    .A_N(_3181_));
 sg13g2_a21oi_1 _5432_ (.A1(_3451_),
    .A2(_0934_),
    .Y(_0935_),
    .B1(net2302));
 sg13g2_nor2b_1 _5433_ (.A(_0930_),
    .B_N(_0935_),
    .Y(_0936_));
 sg13g2_o21ai_1 _5434_ (.B1(_0936_),
    .Y(_0937_),
    .A1(net2419),
    .A2(_0928_));
 sg13g2_or3_1 _5435_ (.A(_0918_),
    .B(_0925_),
    .C(_0937_),
    .X(_0938_));
 sg13g2_nand3_1 _5436_ (.B(_0895_),
    .C(_0938_),
    .A(net2038),
    .Y(_0939_));
 sg13g2_nor2_1 _5437_ (.A(net1978),
    .B(_0864_),
    .Y(_0940_));
 sg13g2_nor3_2 _5438_ (.A(net2461),
    .B(_3095_),
    .C(net2009),
    .Y(_0941_));
 sg13g2_nor3_1 _5439_ (.A(net2539),
    .B(_3526_),
    .C(net2009),
    .Y(_0942_));
 sg13g2_nand3_1 _5440_ (.B(net2249),
    .C(net2422),
    .A(net2093),
    .Y(_0943_));
 sg13g2_o21ai_1 _5441_ (.B1(_0943_),
    .Y(_0945_),
    .A1(net2520),
    .A2(_0218_));
 sg13g2_nor4_2 _5442_ (.A(net2503),
    .B(_0941_),
    .C(_0942_),
    .Y(_0946_),
    .D(_0945_));
 sg13g2_nand3_1 _5443_ (.B(net2247),
    .C(net2226),
    .A(net2250),
    .Y(_0947_));
 sg13g2_nand2_2 _5444_ (.Y(_0948_),
    .A(net2135),
    .B(_0947_));
 sg13g2_a21oi_1 _5445_ (.A1(_3053_),
    .A2(_0948_),
    .Y(_0949_),
    .B1(net2416));
 sg13g2_nor3_2 _5446_ (.A(net2453),
    .B(net2277),
    .C(net2228),
    .Y(_0950_));
 sg13g2_nand2b_2 _5447_ (.Y(_0951_),
    .B(net2149),
    .A_N(_0950_));
 sg13g2_and2_2 _5448_ (.A(net2101),
    .B(_3230_),
    .X(_0952_));
 sg13g2_nand2_1 _5449_ (.Y(_0953_),
    .A(net2101),
    .B(_3230_));
 sg13g2_a21oi_1 _5450_ (.A1(_0951_),
    .A2(_0953_),
    .Y(_0954_),
    .B1(net2431));
 sg13g2_nand2_1 _5451_ (.Y(_0956_),
    .A(net2506),
    .B(_0575_));
 sg13g2_nor3_1 _5452_ (.A(_0949_),
    .B(_0954_),
    .C(_0956_),
    .Y(_0957_));
 sg13g2_o21ai_1 _5453_ (.B1(net2379),
    .Y(_0958_),
    .A1(_0946_),
    .A2(_0957_));
 sg13g2_o21ai_1 _5454_ (.B1(_0919_),
    .Y(_0959_),
    .A1(net2601),
    .A2(_2991_));
 sg13g2_o21ai_1 _5455_ (.B1(net2318),
    .Y(_0960_),
    .A1(_0209_),
    .A2(_0959_));
 sg13g2_nand2_1 _5456_ (.Y(_0961_),
    .A(_3286_),
    .B(_0227_));
 sg13g2_a21oi_1 _5457_ (.A1(net2328),
    .A2(_0961_),
    .Y(_0962_),
    .B1(net2378));
 sg13g2_nand2_1 _5458_ (.Y(_0963_),
    .A(net2431),
    .B(_0235_));
 sg13g2_nand4_1 _5459_ (.B(_0960_),
    .C(_0962_),
    .A(_0228_),
    .Y(_0964_),
    .D(_0963_));
 sg13g2_nand2_1 _5460_ (.Y(_0965_),
    .A(_3283_),
    .B(_0230_));
 sg13g2_a221oi_1 _5461_ (.B2(net2203),
    .C1(net2300),
    .B1(_0965_),
    .A1(_0958_),
    .Y(_0967_),
    .A2(_0964_));
 sg13g2_o21ai_1 _5462_ (.B1(net2328),
    .Y(_0968_),
    .A1(_0190_),
    .A2(_0695_));
 sg13g2_o21ai_1 _5463_ (.B1(_0582_),
    .Y(_0969_),
    .A1(net2332),
    .A2(net2318));
 sg13g2_mux2_2 _5464_ (.A0(_3266_),
    .A1(_0427_),
    .S(net2108),
    .X(_0970_));
 sg13g2_o21ai_1 _5465_ (.B1(_0970_),
    .Y(_0971_),
    .A1(_3250_),
    .A2(_3253_));
 sg13g2_nand2_1 _5466_ (.Y(_0972_),
    .A(net2510),
    .B(_0971_));
 sg13g2_nand3_1 _5467_ (.B(_0969_),
    .C(_0972_),
    .A(_0968_),
    .Y(_0973_));
 sg13g2_a221oi_1 _5468_ (.B2(net2379),
    .C1(_0580_),
    .B1(_0973_),
    .A1(net2021),
    .Y(_0974_),
    .A2(_3451_));
 sg13g2_or3_1 _5469_ (.A(net2037),
    .B(_0967_),
    .C(_0974_),
    .X(_0975_));
 sg13g2_o21ai_1 _5470_ (.B1(net2258),
    .Y(_0976_),
    .A1(net2209),
    .A2(_3151_));
 sg13g2_nand2_2 _5471_ (.Y(_0978_),
    .A(net2173),
    .B(_0976_));
 sg13g2_a21oi_1 _5472_ (.A1(net2033),
    .A2(net2209),
    .Y(_0979_),
    .B1(_3467_));
 sg13g2_o21ai_1 _5473_ (.B1(_0979_),
    .Y(_0980_),
    .A1(net2565),
    .A2(_0978_));
 sg13g2_o21ai_1 _5474_ (.B1(net2259),
    .Y(_0981_),
    .A1(_2948_),
    .A2(_3151_));
 sg13g2_nand3_1 _5475_ (.B(net2078),
    .C(_0981_),
    .A(net2152),
    .Y(_0982_));
 sg13g2_nor4_1 _5476_ (.A(net2588),
    .B(net2152),
    .C(net2259),
    .D(_3224_),
    .Y(_0983_));
 sg13g2_nor3_1 _5477_ (.A(net2528),
    .B(_0473_),
    .C(_0983_),
    .Y(_0984_));
 sg13g2_o21ai_1 _5478_ (.B1(_0984_),
    .Y(_0985_),
    .A1(net2588),
    .A2(_0982_));
 sg13g2_a22oi_1 _5479_ (.Y(_0986_),
    .B1(_0981_),
    .B2(net2152),
    .A2(_3169_),
    .A1(net2216));
 sg13g2_o21ai_1 _5480_ (.B1(net2510),
    .Y(_0987_),
    .A1(net2341),
    .A2(_0986_));
 sg13g2_a21o_1 _5481_ (.A2(_0985_),
    .A1(_0980_),
    .B1(_0987_),
    .X(_0989_));
 sg13g2_nor2_1 _5482_ (.A(net2313),
    .B(_0820_),
    .Y(_0990_));
 sg13g2_nand3_1 _5483_ (.B(_0604_),
    .C(_0990_),
    .A(_0593_),
    .Y(_0991_));
 sg13g2_nor3_1 _5484_ (.A(net2325),
    .B(_3274_),
    .C(_0471_),
    .Y(_0992_));
 sg13g2_o21ai_1 _5485_ (.B1(_0992_),
    .Y(_0993_),
    .A1(net2033),
    .A2(_3354_));
 sg13g2_nand4_1 _5486_ (.B(_0989_),
    .C(_0991_),
    .A(net2380),
    .Y(_0994_),
    .D(_0993_));
 sg13g2_nor2_1 _5487_ (.A(net2245),
    .B(_0729_),
    .Y(_0995_));
 sg13g2_o21ai_1 _5488_ (.B1(net2033),
    .Y(_0996_),
    .A1(_3223_),
    .A2(_0471_));
 sg13g2_a22oi_1 _5489_ (.Y(_0997_),
    .B1(_0995_),
    .B2(net2023),
    .A2(_0981_),
    .A1(net2152));
 sg13g2_nand2_1 _5490_ (.Y(_0998_),
    .A(_0996_),
    .B(_0997_));
 sg13g2_o21ai_1 _5491_ (.B1(net2588),
    .Y(_0999_),
    .A1(_2273_),
    .A2(net2216));
 sg13g2_o21ai_1 _5492_ (.B1(net2565),
    .Y(_1000_),
    .A1(net2259),
    .A2(net2228));
 sg13g2_nand4_1 _5493_ (.B(net2106),
    .C(_0999_),
    .A(net2545),
    .Y(_1001_),
    .D(_1000_));
 sg13g2_nand3_1 _5494_ (.B(_0604_),
    .C(_1001_),
    .A(_0474_),
    .Y(_1002_));
 sg13g2_nor2_1 _5495_ (.A(net2126),
    .B(_0976_),
    .Y(_1003_));
 sg13g2_nand2_1 _5496_ (.Y(_1004_),
    .A(net2175),
    .B(_0452_));
 sg13g2_nor3_1 _5497_ (.A(_3354_),
    .B(_3455_),
    .C(_1003_),
    .Y(_1005_));
 sg13g2_nor4_1 _5498_ (.A(net2386),
    .B(_3354_),
    .C(_3419_),
    .D(_0561_),
    .Y(_1006_));
 sg13g2_a21oi_2 _5499_ (.B1(_1005_),
    .Y(_1007_),
    .A2(_1006_),
    .A1(_1004_));
 sg13g2_a22oi_1 _5500_ (.Y(_1008_),
    .B1(_1002_),
    .B2(net2203),
    .A2(_0998_),
    .A1(_3459_));
 sg13g2_nand4_1 _5501_ (.B(_0994_),
    .C(_1007_),
    .A(net2294),
    .Y(_1010_),
    .D(_1008_));
 sg13g2_a21oi_1 _5502_ (.A1(net2038),
    .A2(_1010_),
    .Y(_1011_),
    .B1(net1977));
 sg13g2_a221oi_1 _5503_ (.B2(_1011_),
    .C1(net1976),
    .B1(_0975_),
    .A1(_0939_),
    .Y(_1012_),
    .A2(_0940_));
 sg13g2_o21ai_1 _5504_ (.B1(_3505_),
    .Y(_1013_),
    .A1(_0805_),
    .A2(_1012_));
 sg13g2_nand2_1 _5505_ (.Y(_1014_),
    .A(net2120),
    .B(_3493_));
 sg13g2_nand4_1 _5506_ (.B(net2005),
    .C(net1994),
    .A(_0224_),
    .Y(_1015_),
    .D(_1014_));
 sg13g2_a22oi_1 _5507_ (.Y(_1016_),
    .B1(_1015_),
    .B2(net2549),
    .A2(_0287_),
    .A1(net2478));
 sg13g2_nand2_1 _5508_ (.Y(_1017_),
    .A(_0747_),
    .B(_1016_));
 sg13g2_mux2_1 _5509_ (.A0(net2234),
    .A1(_3182_),
    .S(net2282),
    .X(_1018_));
 sg13g2_a21oi_2 _5510_ (.B1(net2570),
    .Y(_1019_),
    .A2(_1018_),
    .A1(net2112));
 sg13g2_o21ai_1 _5511_ (.B1(net2571),
    .Y(_1021_),
    .A1(net2284),
    .A2(net2235));
 sg13g2_a21oi_1 _5512_ (.A1(_3011_),
    .A2(_3397_),
    .Y(_1022_),
    .B1(_1021_));
 sg13g2_o21ai_1 _5513_ (.B1(net2529),
    .Y(_1023_),
    .A1(_1019_),
    .A2(_1022_));
 sg13g2_nor2_1 _5514_ (.A(net2110),
    .B(net2341),
    .Y(_1024_));
 sg13g2_nor3_1 _5515_ (.A(net2418),
    .B(_2853_),
    .C(net2072),
    .Y(_1025_));
 sg13g2_a221oi_1 _5516_ (.B2(net2445),
    .C1(_1025_),
    .B1(_0744_),
    .A1(net2166),
    .Y(_1026_),
    .A2(net2343));
 sg13g2_nand2_1 _5517_ (.Y(_1027_),
    .A(_1023_),
    .B(_1026_));
 sg13g2_nor2_1 _5518_ (.A(net2512),
    .B(_0617_),
    .Y(_1028_));
 sg13g2_a21oi_1 _5519_ (.A1(_1027_),
    .A2(_1028_),
    .Y(_1029_),
    .B1(net2396));
 sg13g2_a21oi_1 _5520_ (.A1(_3018_),
    .A2(_0754_),
    .Y(_1030_),
    .B1(_0638_));
 sg13g2_nor2_2 _5521_ (.A(net2546),
    .B(net2105),
    .Y(_1032_));
 sg13g2_a221oi_1 _5522_ (.B2(net2550),
    .C1(net2495),
    .B1(_0752_),
    .A1(net2412),
    .Y(_1033_),
    .A2(_0167_));
 sg13g2_o21ai_1 _5523_ (.B1(_1033_),
    .Y(_1034_),
    .A1(net2550),
    .A2(_1030_));
 sg13g2_nand3_1 _5524_ (.B(net2006),
    .C(_0731_),
    .A(net2025),
    .Y(_1035_));
 sg13g2_nor3_2 _5525_ (.A(net2164),
    .B(net2067),
    .C(_0258_),
    .Y(_1036_));
 sg13g2_a21oi_1 _5526_ (.A1(net2084),
    .A2(_3352_),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_nor3_2 _5527_ (.A(net2138),
    .B(net2250),
    .C(net2356),
    .Y(_1038_));
 sg13g2_nand2_2 _5528_ (.Y(_1039_),
    .A(net2098),
    .B(_0300_));
 sg13g2_o21ai_1 _5529_ (.B1(net2486),
    .Y(_1040_),
    .A1(net2417),
    .A2(_1039_));
 sg13g2_a221oi_1 _5530_ (.B2(net2408),
    .C1(_1040_),
    .B1(_1038_),
    .A1(net2441),
    .Y(_1041_),
    .A2(_1037_));
 sg13g2_o21ai_1 _5531_ (.B1(net2018),
    .Y(_1042_),
    .A1(_3220_),
    .A2(_0738_));
 sg13g2_a22oi_1 _5532_ (.Y(_1043_),
    .B1(_1042_),
    .B2(net2343),
    .A2(_1035_),
    .A1(net2478));
 sg13g2_a21oi_1 _5533_ (.A1(_1041_),
    .A2(_1043_),
    .Y(_1044_),
    .B1(net2382));
 sg13g2_a221oi_1 _5534_ (.B2(_1044_),
    .C1(net2302),
    .B1(_1034_),
    .A1(_1017_),
    .Y(_1045_),
    .A2(_1029_));
 sg13g2_a21oi_2 _5535_ (.B1(net2576),
    .Y(_1046_),
    .A2(net1993),
    .A1(net1996));
 sg13g2_nand3_1 _5536_ (.B(_3553_),
    .C(net1993),
    .A(net2015),
    .Y(_1047_));
 sg13g2_o21ai_1 _5537_ (.B1(net2321),
    .Y(_1048_),
    .A1(_1046_),
    .A2(_1047_));
 sg13g2_o21ai_1 _5538_ (.B1(net2181),
    .Y(_1049_),
    .A1(net2086),
    .A2(_0306_));
 sg13g2_o21ai_1 _5539_ (.B1(_1049_),
    .Y(_1050_),
    .A1(_3576_),
    .A2(net2002));
 sg13g2_nand3_1 _5540_ (.B(_3079_),
    .C(_3161_),
    .A(net2269),
    .Y(_1051_));
 sg13g2_nand3_1 _5541_ (.B(net2052),
    .C(_1051_),
    .A(net2180),
    .Y(_1053_));
 sg13g2_o21ai_1 _5542_ (.B1(_1053_),
    .Y(_1054_),
    .A1(_3035_),
    .A2(net2058));
 sg13g2_a22oi_1 _5543_ (.Y(_1055_),
    .B1(_1054_),
    .B2(net2307),
    .A2(_1050_),
    .A1(net2310));
 sg13g2_a21oi_1 _5544_ (.A1(_1048_),
    .A2(_1055_),
    .Y(_1056_),
    .B1(net2397));
 sg13g2_nand3_1 _5545_ (.B(_3245_),
    .C(net2053),
    .A(net2177),
    .Y(_1057_));
 sg13g2_nor2_2 _5546_ (.A(_3235_),
    .B(net1992),
    .Y(_1058_));
 sg13g2_nor2_1 _5547_ (.A(_0320_),
    .B(_1058_),
    .Y(_1059_));
 sg13g2_o21ai_1 _5548_ (.B1(net2577),
    .Y(_1060_),
    .A1(_0320_),
    .A2(_1058_));
 sg13g2_nor3_1 _5549_ (.A(net2558),
    .B(_0329_),
    .C(_1058_),
    .Y(_1061_));
 sg13g2_a21oi_1 _5550_ (.A1(_3248_),
    .A2(_3313_),
    .Y(_1062_),
    .B1(net2532));
 sg13g2_a221oi_1 _5551_ (.B2(_1059_),
    .C1(net2201),
    .B1(_1062_),
    .A1(_1060_),
    .Y(_1064_),
    .A2(_1061_));
 sg13g2_or3_2 _5552_ (.A(net2154),
    .B(net2060),
    .C(_0427_),
    .X(_1065_));
 sg13g2_nor2_1 _5553_ (.A(net2574),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_nor2_1 _5554_ (.A(_3266_),
    .B(_3509_),
    .Y(_1067_));
 sg13g2_nand3_1 _5555_ (.B(net2242),
    .C(_3267_),
    .A(net2179),
    .Y(_1068_));
 sg13g2_nor3_1 _5556_ (.A(_0296_),
    .B(_1066_),
    .C(_1067_),
    .Y(_1069_));
 sg13g2_nand3_1 _5557_ (.B(net2242),
    .C(_2691_),
    .A(net2184),
    .Y(_1070_));
 sg13g2_nand3_1 _5558_ (.B(net2271),
    .C(_2991_),
    .A(net2178),
    .Y(_1071_));
 sg13g2_nand4_1 _5559_ (.B(net2003),
    .C(_1070_),
    .A(net2013),
    .Y(_1072_),
    .D(_1071_));
 sg13g2_a21oi_1 _5560_ (.A1(_3289_),
    .A2(_1072_),
    .Y(_1073_),
    .B1(net2296));
 sg13g2_o21ai_1 _5561_ (.B1(_1073_),
    .Y(_1075_),
    .A1(_3460_),
    .A2(_1069_));
 sg13g2_nand3_1 _5562_ (.B(net1998),
    .C(_1049_),
    .A(net2014),
    .Y(_1076_));
 sg13g2_o21ai_1 _5563_ (.B1(net2183),
    .Y(_1077_),
    .A1(net2085),
    .A2(_2218_));
 sg13g2_a21oi_1 _5564_ (.A1(_1065_),
    .A2(_1077_),
    .Y(_1078_),
    .B1(net2437));
 sg13g2_a221oi_1 _5565_ (.B2(net2342),
    .C1(_1078_),
    .B1(_1076_),
    .A1(net2480),
    .Y(_1079_),
    .A2(_1050_));
 sg13g2_nor2b_1 _5566_ (.A(_1079_),
    .B_N(_0124_),
    .Y(_1080_));
 sg13g2_nor4_1 _5567_ (.A(_1056_),
    .B(_1064_),
    .C(_1075_),
    .D(_1080_),
    .Y(_1081_));
 sg13g2_nor3_1 _5568_ (.A(net2039),
    .B(_1045_),
    .C(_1081_),
    .Y(_1082_));
 sg13g2_nand4_1 _5569_ (.B(net2003),
    .C(net1995),
    .A(net2017),
    .Y(_1083_),
    .D(_1077_));
 sg13g2_o21ai_1 _5570_ (.B1(net2032),
    .Y(_1084_),
    .A1(net2082),
    .A2(_3088_));
 sg13g2_o21ai_1 _5571_ (.B1(net2342),
    .Y(_1086_),
    .A1(_0318_),
    .A2(_1084_));
 sg13g2_nand3_1 _5572_ (.B(_3245_),
    .C(_0166_),
    .A(net2177),
    .Y(_1087_));
 sg13g2_nand2_1 _5573_ (.Y(_1088_),
    .A(_0319_),
    .B(_1087_));
 sg13g2_a221oi_1 _5574_ (.B2(net2449),
    .C1(net2500),
    .B1(_1088_),
    .A1(net2480),
    .Y(_1089_),
    .A2(_1083_));
 sg13g2_nand3_1 _5575_ (.B(net2078),
    .C(_3267_),
    .A(net2178),
    .Y(_1090_));
 sg13g2_nand4_1 _5576_ (.B(net2017),
    .C(net2003),
    .A(net2500),
    .Y(_1091_),
    .D(_1090_));
 sg13g2_a21oi_1 _5577_ (.A1(net2533),
    .A2(_0354_),
    .Y(_1092_),
    .B1(_1091_));
 sg13g2_a21oi_1 _5578_ (.A1(_1086_),
    .A2(_1089_),
    .Y(_1093_),
    .B1(_1092_));
 sg13g2_nor2_1 _5579_ (.A(net2518),
    .B(_1088_),
    .Y(_1094_));
 sg13g2_nand3_1 _5580_ (.B(net2260),
    .C(_3222_),
    .A(net2474),
    .Y(_1095_));
 sg13g2_nand4_1 _5581_ (.B(net2000),
    .C(net1992),
    .A(net2518),
    .Y(_1097_),
    .D(_1095_));
 sg13g2_nor2_1 _5582_ (.A(net2383),
    .B(_1094_),
    .Y(_1098_));
 sg13g2_a221oi_1 _5583_ (.B2(_1098_),
    .C1(net2294),
    .B1(_1097_),
    .A1(net2383),
    .Y(_1099_),
    .A2(_1093_));
 sg13g2_o21ai_1 _5584_ (.B1(net2000),
    .Y(_1100_),
    .A1(_3247_),
    .A2(_3312_));
 sg13g2_a221oi_1 _5585_ (.B2(net2601),
    .C1(net2518),
    .B1(_1100_),
    .A1(net2533),
    .Y(_1101_),
    .A2(_0165_));
 sg13g2_a221oi_1 _5586_ (.B2(_1101_),
    .C1(net2397),
    .B1(_1060_),
    .A1(net2518),
    .Y(_1102_),
    .A2(_1059_));
 sg13g2_o21ai_1 _5587_ (.B1(net2000),
    .Y(_1103_),
    .A1(_2306_),
    .A2(_3247_));
 sg13g2_nor2_1 _5588_ (.A(net2341),
    .B(net2192),
    .Y(_1104_));
 sg13g2_a21oi_1 _5589_ (.A1(_1103_),
    .A2(_1104_),
    .Y(_1105_),
    .B1(net2303));
 sg13g2_o21ai_1 _5590_ (.B1(_1105_),
    .Y(_1106_),
    .A1(_3460_),
    .A2(_1059_));
 sg13g2_nand3_1 _5591_ (.B(net1999),
    .C(_1090_),
    .A(net2017),
    .Y(_1108_));
 sg13g2_and3_1 _5592_ (.X(_1109_),
    .A(net2467),
    .B(net2205),
    .C(_1108_));
 sg13g2_a21oi_1 _5593_ (.A1(net2230),
    .A2(_3256_),
    .Y(_1110_),
    .B1(_0324_));
 sg13g2_nor4_1 _5594_ (.A(net2383),
    .B(_3419_),
    .C(_0561_),
    .D(_1110_),
    .Y(_1111_));
 sg13g2_nor4_1 _5595_ (.A(_1102_),
    .B(_1106_),
    .C(_1109_),
    .D(_1111_),
    .Y(_1112_));
 sg13g2_nor3_1 _5596_ (.A(net2036),
    .B(_1099_),
    .C(_1112_),
    .Y(_1113_));
 sg13g2_o21ai_1 _5597_ (.B1(net1980),
    .Y(_1114_),
    .A1(_1082_),
    .A2(_1113_));
 sg13g2_nand2_1 _5598_ (.Y(_1115_),
    .A(net2050),
    .B(_3192_));
 sg13g2_a21oi_1 _5599_ (.A1(net2050),
    .A2(_3192_),
    .Y(_1116_),
    .B1(net2538));
 sg13g2_nand3_1 _5600_ (.B(_2892_),
    .C(net2025),
    .A(net2046),
    .Y(_1117_));
 sg13g2_nand3_1 _5601_ (.B(_2750_),
    .C(_3192_),
    .A(net2578),
    .Y(_1119_));
 sg13g2_and3_1 _5602_ (.X(_1120_),
    .A(net2538),
    .B(_1117_),
    .C(_1119_));
 sg13g2_o21ai_1 _5603_ (.B1(net2501),
    .Y(_1121_),
    .A1(_1116_),
    .A2(_1120_));
 sg13g2_nand2_1 _5604_ (.Y(_1122_),
    .A(net2579),
    .B(_2449_));
 sg13g2_mux2_1 _5605_ (.A0(_2449_),
    .A1(_0643_),
    .S(net2559),
    .X(_1123_));
 sg13g2_a21o_1 _5606_ (.A2(_1123_),
    .A1(net2050),
    .B1(net2521),
    .X(_1124_));
 sg13g2_a21oi_1 _5607_ (.A1(net2050),
    .A2(_2863_),
    .Y(_1125_),
    .B1(_3062_));
 sg13g2_nor3_1 _5608_ (.A(net2133),
    .B(net2240),
    .C(net2308),
    .Y(_1126_));
 sg13g2_o21ai_1 _5609_ (.B1(net2470),
    .Y(_1127_),
    .A1(_2460_),
    .A2(_3104_));
 sg13g2_a21oi_1 _5610_ (.A1(_1124_),
    .A2(_1127_),
    .Y(_1128_),
    .B1(net2502));
 sg13g2_nor4_1 _5611_ (.A(net2388),
    .B(_1125_),
    .C(_1126_),
    .D(_1128_),
    .Y(_1130_));
 sg13g2_or2_1 _5612_ (.X(_1131_),
    .B(_0177_),
    .A(net2029));
 sg13g2_nor3_1 _5613_ (.A(net2581),
    .B(net2029),
    .C(_0177_),
    .Y(_1132_));
 sg13g2_o21ai_1 _5614_ (.B1(_0627_),
    .Y(_1133_),
    .A1(net2581),
    .A2(_1131_));
 sg13g2_nor2_1 _5615_ (.A(net2417),
    .B(net2029),
    .Y(_1134_));
 sg13g2_a22oi_1 _5616_ (.Y(_1135_),
    .B1(_1134_),
    .B2(_3577_),
    .A2(_1133_),
    .A1(net2524));
 sg13g2_nand2_1 _5617_ (.Y(_1136_),
    .A(_3146_),
    .B(net2061));
 sg13g2_a22oi_1 _5618_ (.Y(_1137_),
    .B1(_3509_),
    .B2(_3132_),
    .A2(net2061),
    .A1(_3146_));
 sg13g2_nor3_1 _5619_ (.A(net2435),
    .B(_0623_),
    .C(_1137_),
    .Y(_1138_));
 sg13g2_nor2_1 _5620_ (.A(net2493),
    .B(_1138_),
    .Y(_1139_));
 sg13g2_o21ai_1 _5621_ (.B1(_1139_),
    .Y(_1141_),
    .A1(_0920_),
    .A2(_1135_));
 sg13g2_a21oi_1 _5622_ (.A1(net2044),
    .A2(_0649_),
    .Y(_1142_),
    .B1(net2314));
 sg13g2_or2_1 _5623_ (.X(_1143_),
    .B(_0648_),
    .A(_3149_));
 sg13g2_nand3_1 _5624_ (.B(_3077_),
    .C(net2208),
    .A(net2374),
    .Y(_1144_));
 sg13g2_a21o_1 _5625_ (.A2(_1144_),
    .A1(_3085_),
    .B1(_3594_),
    .X(_1145_));
 sg13g2_o21ai_1 _5626_ (.B1(net2306),
    .Y(_1146_),
    .A1(_1143_),
    .A2(_1145_));
 sg13g2_nor2_1 _5627_ (.A(_3052_),
    .B(_0396_),
    .Y(_1147_));
 sg13g2_a21oi_1 _5628_ (.A1(_3176_),
    .A2(_3200_),
    .Y(_1148_),
    .B1(_0626_));
 sg13g2_o21ai_1 _5629_ (.B1(_1146_),
    .Y(_1149_),
    .A1(net2308),
    .A2(_1148_));
 sg13g2_nor4_2 _5630_ (.A(net2377),
    .B(_1142_),
    .C(_1147_),
    .Y(_1150_),
    .D(_1149_));
 sg13g2_a22oi_1 _5631_ (.Y(_1152_),
    .B1(_1141_),
    .B2(_1150_),
    .A2(_1130_),
    .A1(_1121_));
 sg13g2_mux2_2 _5632_ (.A0(_3266_),
    .A1(_3274_),
    .S(net2107),
    .X(_1153_));
 sg13g2_nand2b_2 _5633_ (.Y(_1154_),
    .B(_3277_),
    .A_N(_3269_));
 sg13g2_nor2_1 _5634_ (.A(net2587),
    .B(_1153_),
    .Y(_1155_));
 sg13g2_nand2_1 _5635_ (.Y(_1156_),
    .A(net2566),
    .B(_1154_));
 sg13g2_o21ai_1 _5636_ (.B1(_0970_),
    .Y(_1157_),
    .A1(net2587),
    .A2(_1153_));
 sg13g2_nor3_2 _5637_ (.A(net2313),
    .B(_3270_),
    .C(_3294_),
    .Y(_1158_));
 sg13g2_a21oi_1 _5638_ (.A1(net2338),
    .A2(_1157_),
    .Y(_1159_),
    .B1(_1158_));
 sg13g2_nor2_1 _5639_ (.A(_0697_),
    .B(_1158_),
    .Y(_1160_));
 sg13g2_and2_1 _5640_ (.A(_0698_),
    .B(_1159_),
    .X(_1161_));
 sg13g2_and2_1 _5641_ (.A(net2104),
    .B(_0170_),
    .X(_1163_));
 sg13g2_o21ai_1 _5642_ (.B1(_3410_),
    .Y(_1164_),
    .A1(net2020),
    .A2(_1163_));
 sg13g2_a21oi_2 _5643_ (.B1(net2378),
    .Y(_1165_),
    .A2(_0684_),
    .A1(net2318));
 sg13g2_nand2b_1 _5644_ (.Y(_1166_),
    .B(_3478_),
    .A_N(_0266_));
 sg13g2_nand2_1 _5645_ (.Y(_1167_),
    .A(_0682_),
    .B(_1166_));
 sg13g2_nand2_1 _5646_ (.Y(_1168_),
    .A(_3478_),
    .B(_0426_));
 sg13g2_nand4_1 _5647_ (.B(_1164_),
    .C(_1165_),
    .A(_0683_),
    .Y(_1169_),
    .D(_1168_));
 sg13g2_o21ai_1 _5648_ (.B1(net2300),
    .Y(_1170_),
    .A1(_1167_),
    .A2(_1169_));
 sg13g2_a21oi_1 _5649_ (.A1(net2294),
    .A2(_0677_),
    .Y(_1171_),
    .B1(net2037));
 sg13g2_o21ai_1 _5650_ (.B1(_1171_),
    .Y(_1172_),
    .A1(_1161_),
    .A2(_1170_));
 sg13g2_o21ai_1 _5651_ (.B1(net2306),
    .Y(_1174_),
    .A1(_3030_),
    .A2(_3080_));
 sg13g2_nand3_1 _5652_ (.B(_3096_),
    .C(_1174_),
    .A(net2389),
    .Y(_1175_));
 sg13g2_nand2_1 _5653_ (.Y(_1176_),
    .A(_2449_),
    .B(_3075_));
 sg13g2_o21ai_1 _5654_ (.B1(net2439),
    .Y(_1177_),
    .A1(_2460_),
    .A2(net2034));
 sg13g2_a21oi_1 _5655_ (.A1(_0673_),
    .A2(_1177_),
    .Y(_1178_),
    .B1(net2483));
 sg13g2_nand3_1 _5656_ (.B(_2273_),
    .C(net2053),
    .A(net2098),
    .Y(_1179_));
 sg13g2_a21oi_2 _5657_ (.B1(net2520),
    .Y(_1180_),
    .A2(_1179_),
    .A1(_3031_));
 sg13g2_a21oi_1 _5658_ (.A1(_3031_),
    .A2(_1179_),
    .Y(_1181_),
    .B1(net2308));
 sg13g2_nor3_1 _5659_ (.A(net2041),
    .B(net2034),
    .C(_3097_),
    .Y(_1182_));
 sg13g2_nor3_1 _5660_ (.A(_3025_),
    .B(net2070),
    .C(_3174_),
    .Y(_1183_));
 sg13g2_nor3_1 _5661_ (.A(net2336),
    .B(_1182_),
    .C(_1183_),
    .Y(_1185_));
 sg13g2_nor4_2 _5662_ (.A(_1175_),
    .B(_1178_),
    .C(_1181_),
    .Y(_1186_),
    .D(_1185_));
 sg13g2_nor3_1 _5663_ (.A(net2544),
    .B(_3044_),
    .C(_0656_),
    .Y(_1187_));
 sg13g2_nor3_1 _5664_ (.A(net2429),
    .B(_3044_),
    .C(_3093_),
    .Y(_1188_));
 sg13g2_a21oi_2 _5665_ (.B1(net2148),
    .Y(_1189_),
    .A2(net2087),
    .A1(net2357));
 sg13g2_nor3_1 _5666_ (.A(net2416),
    .B(_3044_),
    .C(_1189_),
    .Y(_1190_));
 sg13g2_nor4_1 _5667_ (.A(net2484),
    .B(_1187_),
    .C(_1188_),
    .D(_1190_),
    .Y(_1191_));
 sg13g2_a22oi_1 _5668_ (.Y(_1192_),
    .B1(net2041),
    .B2(_3055_),
    .A2(net2045),
    .A1(net2563));
 sg13g2_a21oi_1 _5669_ (.A1(_0655_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(net2325));
 sg13g2_mux2_1 _5670_ (.A0(_3055_),
    .A1(_3230_),
    .S(net2101),
    .X(_1194_));
 sg13g2_a21o_1 _5671_ (.A2(_1194_),
    .A1(_3061_),
    .B1(net2391),
    .X(_1196_));
 sg13g2_nor4_1 _5672_ (.A(_3059_),
    .B(_1191_),
    .C(_1193_),
    .D(_1196_),
    .Y(_1197_));
 sg13g2_o21ai_1 _5673_ (.B1(_3431_),
    .Y(_1198_),
    .A1(_1186_),
    .A2(_1197_));
 sg13g2_and3_1 _5674_ (.X(_1199_),
    .A(net1977),
    .B(_1172_),
    .C(_1198_));
 sg13g2_o21ai_1 _5675_ (.B1(_1199_),
    .Y(_1200_),
    .A1(_3375_),
    .A2(_1152_));
 sg13g2_nand3_1 _5676_ (.B(_1114_),
    .C(_1200_),
    .A(_3309_),
    .Y(_1201_));
 sg13g2_and2_1 _5677_ (.A(_3115_),
    .B(net2016),
    .X(_1202_));
 sg13g2_a21oi_2 _5678_ (.B1(net2182),
    .Y(_1203_),
    .A2(_3117_),
    .A1(_3114_));
 sg13g2_a21oi_2 _5679_ (.B1(_0452_),
    .Y(_1204_),
    .A2(net2032),
    .A1(_3118_));
 sg13g2_a21oi_1 _5680_ (.A1(net2576),
    .A2(_1202_),
    .Y(_1205_),
    .B1(_2185_));
 sg13g2_o21ai_1 _5681_ (.B1(_1205_),
    .Y(_1207_),
    .A1(_1203_),
    .A2(_1204_));
 sg13g2_a21oi_1 _5682_ (.A1(_0807_),
    .A2(_0814_),
    .Y(_1208_),
    .B1(net2468));
 sg13g2_nor2_1 _5683_ (.A(net2404),
    .B(_0385_),
    .Y(_1209_));
 sg13g2_o21ai_1 _5684_ (.B1(net2515),
    .Y(_1210_),
    .A1(net2554),
    .A2(net2031));
 sg13g2_a21oi_1 _5685_ (.A1(_0825_),
    .A2(_0847_),
    .Y(_1211_),
    .B1(net2436));
 sg13g2_nor4_1 _5686_ (.A(_1208_),
    .B(_1209_),
    .C(_1210_),
    .D(_1211_),
    .Y(_1212_));
 sg13g2_o21ai_1 _5687_ (.B1(net2415),
    .Y(_1213_),
    .A1(_3436_),
    .A2(_1204_));
 sg13g2_nor3_1 _5688_ (.A(net2597),
    .B(net2245),
    .C(net2239),
    .Y(_1214_));
 sg13g2_a21oi_1 _5689_ (.A1(_3018_),
    .A2(_3161_),
    .Y(_1215_),
    .B1(net2575));
 sg13g2_o21ai_1 _5690_ (.B1(_3085_),
    .Y(_1216_),
    .A1(_1214_),
    .A2(_1215_));
 sg13g2_nand4_1 _5691_ (.B(net2030),
    .C(_0514_),
    .A(net2498),
    .Y(_1218_),
    .D(_1216_));
 sg13g2_a221oi_1 _5692_ (.B2(net2315),
    .C1(_0810_),
    .B1(_1218_),
    .A1(net2481),
    .Y(_1219_),
    .A2(_3133_));
 sg13g2_a221oi_1 _5693_ (.B2(_1219_),
    .C1(net2399),
    .B1(_1213_),
    .A1(_1207_),
    .Y(_1220_),
    .A2(_1212_));
 sg13g2_o21ai_1 _5694_ (.B1(net2182),
    .Y(_1221_),
    .A1(_2901_),
    .A2(_0311_));
 sg13g2_a21oi_1 _5695_ (.A1(_0825_),
    .A2(_1221_),
    .Y(_1222_),
    .B1(net2468));
 sg13g2_a21oi_1 _5696_ (.A1(net2415),
    .A2(_0848_),
    .Y(_1223_),
    .B1(_1222_));
 sg13g2_a21oi_1 _5697_ (.A1(net2554),
    .A2(_0848_),
    .Y(_1224_),
    .B1(_0850_));
 sg13g2_a21oi_1 _5698_ (.A1(_1223_),
    .A2(_1224_),
    .Y(_1225_),
    .B1(net2192));
 sg13g2_nor3_2 _5699_ (.A(net2594),
    .B(net2123),
    .C(_0138_),
    .Y(_1226_));
 sg13g2_o21ai_1 _5700_ (.B1(net2121),
    .Y(_1227_),
    .A1(net2067),
    .A2(_0328_));
 sg13g2_a21oi_1 _5701_ (.A1(_0839_),
    .A2(_1227_),
    .Y(_1229_),
    .B1(net2594));
 sg13g2_nor3_1 _5702_ (.A(_0832_),
    .B(_0835_),
    .C(_1229_),
    .Y(_1230_));
 sg13g2_a221oi_1 _5703_ (.B2(_0140_),
    .C1(_0831_),
    .B1(net2052),
    .A1(net2594),
    .Y(_1231_),
    .A2(_0530_));
 sg13g2_nor3_1 _5704_ (.A(net2200),
    .B(_1230_),
    .C(_1231_),
    .Y(_1232_));
 sg13g2_or4_2 _5705_ (.A(net1985),
    .B(_1220_),
    .C(_1225_),
    .D(_1232_),
    .X(_1233_));
 sg13g2_a21oi_1 _5706_ (.A1(net2240),
    .A2(net2073),
    .Y(_1234_),
    .B1(_3025_));
 sg13g2_o21ai_1 _5707_ (.B1(net2520),
    .Y(_1235_),
    .A1(_0445_),
    .A2(_1234_));
 sg13g2_a22oi_1 _5708_ (.Y(_1236_),
    .B1(_3276_),
    .B2(net2421),
    .A2(_3030_),
    .A1(net2344));
 sg13g2_nand3_1 _5709_ (.B(_1235_),
    .C(_1236_),
    .A(_3580_),
    .Y(_1237_));
 sg13g2_nand2_1 _5710_ (.Y(_1238_),
    .A(_3195_),
    .B(_3575_));
 sg13g2_o21ai_1 _5711_ (.B1(net2471),
    .Y(_1240_),
    .A1(_0464_),
    .A2(_1238_));
 sg13g2_o21ai_1 _5712_ (.B1(net2407),
    .Y(_1241_),
    .A1(_0209_),
    .A2(_0886_));
 sg13g2_a21oi_1 _5713_ (.A1(_2570_),
    .A2(_2982_),
    .Y(_1242_),
    .B1(net2138));
 sg13g2_o21ai_1 _5714_ (.B1(net2539),
    .Y(_1243_),
    .A1(_0886_),
    .A2(_1242_));
 sg13g2_a21oi_1 _5715_ (.A1(net2081),
    .A2(net2440),
    .Y(_1244_),
    .B1(net2503));
 sg13g2_nand4_1 _5716_ (.B(_1241_),
    .C(_1243_),
    .A(_1240_),
    .Y(_1245_),
    .D(_1244_));
 sg13g2_nand3_1 _5717_ (.B(_1237_),
    .C(_1245_),
    .A(net2389),
    .Y(_1246_));
 sg13g2_a21oi_1 _5718_ (.A1(net2046),
    .A2(_0625_),
    .Y(_1247_),
    .B1(net2561));
 sg13g2_a21oi_1 _5719_ (.A1(net2583),
    .A2(_3610_),
    .Y(_1248_),
    .B1(_1247_));
 sg13g2_nand2_1 _5720_ (.Y(_1249_),
    .A(_3195_),
    .B(net2025));
 sg13g2_nand3_1 _5721_ (.B(_3195_),
    .C(net2025),
    .A(net2522),
    .Y(_1251_));
 sg13g2_o21ai_1 _5722_ (.B1(net2464),
    .Y(_1252_),
    .A1(_3610_),
    .A2(_1251_));
 sg13g2_nand2_1 _5723_ (.Y(_1253_),
    .A(net2540),
    .B(_3600_));
 sg13g2_nor2_1 _5724_ (.A(net2087),
    .B(net2212),
    .Y(_1254_));
 sg13g2_a21o_1 _5725_ (.A2(_3549_),
    .A1(net2083),
    .B1(_3028_),
    .X(_1255_));
 sg13g2_nor2_1 _5726_ (.A(_0869_),
    .B(_1253_),
    .Y(_1256_));
 sg13g2_a221oi_1 _5727_ (.B2(_1256_),
    .C1(net2504),
    .B1(_1255_),
    .A1(_1248_),
    .Y(_1257_),
    .A2(_1252_));
 sg13g2_nand2_1 _5728_ (.Y(_1258_),
    .A(net2561),
    .B(_3260_));
 sg13g2_nand4_1 _5729_ (.B(_3195_),
    .C(_3575_),
    .A(net2542),
    .Y(_1259_),
    .D(_1258_));
 sg13g2_o21ai_1 _5730_ (.B1(net2522),
    .Y(_1260_),
    .A1(net2583),
    .A2(_3122_));
 sg13g2_o21ai_1 _5731_ (.B1(_1259_),
    .Y(_1262_),
    .A1(_0869_),
    .A2(_1260_));
 sg13g2_a21oi_1 _5732_ (.A1(net2051),
    .A2(_1262_),
    .Y(_1263_),
    .B1(net2485));
 sg13g2_o21ai_1 _5733_ (.B1(net2377),
    .Y(_1264_),
    .A1(_1257_),
    .A2(_1263_));
 sg13g2_nand3_1 _5734_ (.B(_1246_),
    .C(_1264_),
    .A(net1982),
    .Y(_1265_));
 sg13g2_nand3_1 _5735_ (.B(net2263),
    .C(_3377_),
    .A(net2166),
    .Y(_1266_));
 sg13g2_nand3_1 _5736_ (.B(_0912_),
    .C(_1266_),
    .A(net2012),
    .Y(_1267_));
 sg13g2_or2_1 _5737_ (.X(_1268_),
    .B(_3578_),
    .A(net2029));
 sg13g2_or3_2 _5738_ (.A(net2029),
    .B(net2028),
    .C(_3578_),
    .X(_1269_));
 sg13g2_a21oi_1 _5739_ (.A1(net2071),
    .A2(_3351_),
    .Y(_1270_),
    .B1(_3607_));
 sg13g2_a221oi_1 _5740_ (.B2(net2476),
    .C1(_1270_),
    .B1(_0617_),
    .A1(net2425),
    .Y(_1271_),
    .A2(net2223));
 sg13g2_a22oi_1 _5741_ (.Y(_1273_),
    .B1(_1269_),
    .B2(net2548),
    .A2(_1267_),
    .A1(net2412));
 sg13g2_a21oi_1 _5742_ (.A1(_1271_),
    .A2(_1273_),
    .Y(_1274_),
    .B1(net2193));
 sg13g2_nand4_1 _5743_ (.B(net2048),
    .C(net2044),
    .A(net2561),
    .Y(_1275_),
    .D(_3167_));
 sg13g2_nand3_1 _5744_ (.B(_3173_),
    .C(_3221_),
    .A(net2282),
    .Y(_1276_));
 sg13g2_nand3_1 _5745_ (.B(_0548_),
    .C(_1276_),
    .A(net2110),
    .Y(_1277_));
 sg13g2_nand4_1 _5746_ (.B(net2026),
    .C(_3596_),
    .A(net2581),
    .Y(_1278_),
    .D(_1277_));
 sg13g2_nand3_1 _5747_ (.B(_1275_),
    .C(_1278_),
    .A(net2548),
    .Y(_1279_));
 sg13g2_nand2b_1 _5748_ (.Y(_1280_),
    .B(_0932_),
    .A_N(_0920_));
 sg13g2_a22oi_1 _5749_ (.Y(_1281_),
    .B1(_1280_),
    .B2(net2476),
    .A2(_0927_),
    .A1(net2410));
 sg13g2_a21oi_1 _5750_ (.A1(_1279_),
    .A2(_1281_),
    .Y(_1282_),
    .B1(net2200));
 sg13g2_a21oi_1 _5751_ (.A1(net2170),
    .A2(_3512_),
    .Y(_1284_),
    .B1(net2596));
 sg13g2_nand3_1 _5752_ (.B(_0899_),
    .C(_1284_),
    .A(net2030),
    .Y(_1285_));
 sg13g2_nand2_1 _5753_ (.Y(_1286_),
    .A(net2266),
    .B(_3020_));
 sg13g2_nand3_1 _5754_ (.B(net2052),
    .C(_1286_),
    .A(net2171),
    .Y(_1287_));
 sg13g2_nand3_1 _5755_ (.B(net2276),
    .C(_2240_),
    .A(net2097),
    .Y(_1288_));
 sg13g2_nand4_1 _5756_ (.B(net2005),
    .C(_1287_),
    .A(net2595),
    .Y(_1289_),
    .D(_1288_));
 sg13g2_nand3_1 _5757_ (.B(_1285_),
    .C(_1289_),
    .A(net2329),
    .Y(_1290_));
 sg13g2_nor2_1 _5758_ (.A(_3062_),
    .B(_1287_),
    .Y(_1291_));
 sg13g2_a221oi_1 _5759_ (.B2(net2595),
    .C1(net2549),
    .B1(_3510_),
    .A1(net2167),
    .Y(_1292_),
    .A2(_3340_));
 sg13g2_a22oi_1 _5760_ (.Y(_1293_),
    .B1(_3321_),
    .B2(net2071),
    .A2(_3124_),
    .A1(net2168));
 sg13g2_nand3b_1 _5761_ (.B(net2549),
    .C(_0260_),
    .Y(_1295_),
    .A_N(_1293_));
 sg13g2_a21oi_1 _5762_ (.A1(_0899_),
    .A2(_1292_),
    .Y(_1296_),
    .B1(net2494));
 sg13g2_a221oi_1 _5763_ (.B2(_1296_),
    .C1(_1291_),
    .B1(_1295_),
    .A1(net2323),
    .Y(_1297_),
    .A2(_0903_));
 sg13g2_a21oi_2 _5764_ (.B1(net2396),
    .Y(_1298_),
    .A2(_1297_),
    .A1(_1290_));
 sg13g2_nor4_2 _5765_ (.A(_3432_),
    .B(_1274_),
    .C(_1282_),
    .Y(_1299_),
    .D(_1298_));
 sg13g2_nand3_1 _5766_ (.B(_0339_),
    .C(_1057_),
    .A(net2008),
    .Y(_1300_));
 sg13g2_a21oi_1 _5767_ (.A1(net2599),
    .A2(_0311_),
    .Y(_1301_),
    .B1(net2556));
 sg13g2_nand4_1 _5768_ (.B(net1998),
    .C(_1077_),
    .A(net2013),
    .Y(_1302_),
    .D(_1301_));
 sg13g2_a21oi_1 _5769_ (.A1(net2184),
    .A2(net2052),
    .Y(_1303_),
    .B1(net2534));
 sg13g2_a21oi_1 _5770_ (.A1(_0514_),
    .A2(_1303_),
    .Y(_1304_),
    .B1(net2499));
 sg13g2_nor2b_1 _5771_ (.A(_0340_),
    .B_N(net1992),
    .Y(_1306_));
 sg13g2_a22oi_1 _5772_ (.Y(_1307_),
    .B1(_1302_),
    .B2(_1304_),
    .A2(_1300_),
    .A1(net2311));
 sg13g2_o21ai_1 _5773_ (.B1(_1307_),
    .Y(_1308_),
    .A1(_3062_),
    .A2(_1306_));
 sg13g2_nand4_1 _5774_ (.B(net2019),
    .C(_0339_),
    .A(net2311),
    .Y(_1309_),
    .D(net1992));
 sg13g2_o21ai_1 _5775_ (.B1(_1309_),
    .Y(_1310_),
    .A1(net2311),
    .A2(_1300_));
 sg13g2_o21ai_1 _5776_ (.B1(net2000),
    .Y(_1311_),
    .A1(net2574),
    .A2(net1992));
 sg13g2_nor2_1 _5777_ (.A(_3088_),
    .B(_0736_),
    .Y(_1312_));
 sg13g2_a221oi_1 _5778_ (.B2(_3451_),
    .C1(net1983),
    .B1(_1312_),
    .A1(_3289_),
    .Y(_1313_),
    .A2(_1311_));
 sg13g2_o21ai_1 _5779_ (.B1(_1313_),
    .Y(_1314_),
    .A1(net2400),
    .A2(_1310_));
 sg13g2_a21oi_1 _5780_ (.A1(net2400),
    .A2(_1308_),
    .Y(_1315_),
    .B1(_1314_));
 sg13g2_nor3_2 _5781_ (.A(net1980),
    .B(_1299_),
    .C(_1315_),
    .Y(_1317_));
 sg13g2_nand3_1 _5782_ (.B(_1265_),
    .C(_1317_),
    .A(_1233_),
    .Y(_1318_));
 sg13g2_a21oi_1 _5783_ (.A1(_3035_),
    .A2(_0217_),
    .Y(_1319_),
    .B1(net2429));
 sg13g2_and3_1 _5784_ (.X(_1320_),
    .A(net2407),
    .B(_3142_),
    .C(_3575_));
 sg13g2_nor4_2 _5785_ (.A(net2503),
    .B(_0941_),
    .C(_1319_),
    .Y(_1321_),
    .D(_1320_));
 sg13g2_mux2_1 _5786_ (.A0(net2082),
    .A1(_0950_),
    .S(net2149),
    .X(_1322_));
 sg13g2_nand2_1 _5787_ (.Y(_1323_),
    .A(_3053_),
    .B(_0951_));
 sg13g2_a21oi_1 _5788_ (.A1(_3053_),
    .A2(_0951_),
    .Y(_1324_),
    .B1(net2431));
 sg13g2_a21oi_1 _5789_ (.A1(_3034_),
    .A2(_0948_),
    .Y(_1325_),
    .B1(net2585));
 sg13g2_o21ai_1 _5790_ (.B1(net2507),
    .Y(_1326_),
    .A1(net2526),
    .A2(_1322_));
 sg13g2_nor4_1 _5791_ (.A(_0219_),
    .B(_1324_),
    .C(_1325_),
    .D(_1326_),
    .Y(_1328_));
 sg13g2_mux2_2 _5792_ (.A0(_3171_),
    .A1(_3565_),
    .S(net2135),
    .X(_1329_));
 sg13g2_and2_1 _5793_ (.A(_3271_),
    .B(_1329_),
    .X(_1330_));
 sg13g2_a21oi_1 _5794_ (.A1(net2306),
    .A2(_1330_),
    .Y(_1331_),
    .B1(net2391));
 sg13g2_o21ai_1 _5795_ (.B1(_1331_),
    .Y(_1332_),
    .A1(_1321_),
    .A2(_1328_));
 sg13g2_nand2_2 _5796_ (.Y(_1333_),
    .A(net2024),
    .B(_0230_));
 sg13g2_a21oi_1 _5797_ (.A1(net2024),
    .A2(_0230_),
    .Y(_1334_),
    .B1(net2587));
 sg13g2_o21ai_1 _5798_ (.B1(net2332),
    .Y(_1335_),
    .A1(_0233_),
    .A2(_1334_));
 sg13g2_a21o_2 _5799_ (.A2(_0950_),
    .A1(net2236),
    .B1(net2102),
    .X(_1336_));
 sg13g2_nor2_1 _5800_ (.A(net2585),
    .B(_1336_),
    .Y(_1337_));
 sg13g2_nand2_1 _5801_ (.Y(_1339_),
    .A(_0208_),
    .B(_0951_));
 sg13g2_o21ai_1 _5802_ (.B1(net2318),
    .Y(_1340_),
    .A1(_1337_),
    .A2(_1339_));
 sg13g2_nand4_1 _5803_ (.B(_0962_),
    .C(_1335_),
    .A(_0236_),
    .Y(_1341_),
    .D(_1340_));
 sg13g2_a21oi_2 _5804_ (.B1(net1983),
    .Y(_1342_),
    .A2(_1341_),
    .A1(_1332_));
 sg13g2_nand3_1 _5805_ (.B(net2289),
    .C(net2216),
    .A(net2105),
    .Y(_1343_));
 sg13g2_nand3_1 _5806_ (.B(_0982_),
    .C(_1343_),
    .A(_3150_),
    .Y(_1344_));
 sg13g2_a21oi_1 _5807_ (.A1(net2601),
    .A2(_3017_),
    .Y(_1345_),
    .B1(net2532));
 sg13g2_nand4_1 _5808_ (.B(_0982_),
    .C(_1343_),
    .A(_3150_),
    .Y(_1346_),
    .D(_1345_));
 sg13g2_nor4_2 _5809_ (.A(net2145),
    .B(net2248),
    .C(net2063),
    .Y(_1347_),
    .D(net2210));
 sg13g2_a21oi_2 _5810_ (.B1(net2105),
    .Y(_1348_),
    .A2(_0976_),
    .A1(net2078));
 sg13g2_o21ai_1 _5811_ (.B1(_0485_),
    .Y(_1350_),
    .A1(_1347_),
    .A2(_1348_));
 sg13g2_nand3_1 _5812_ (.B(_1346_),
    .C(_1350_),
    .A(net2510),
    .Y(_1351_));
 sg13g2_nand3_1 _5813_ (.B(net1997),
    .C(_0730_),
    .A(_0416_),
    .Y(_1352_));
 sg13g2_nor3_1 _5814_ (.A(net2308),
    .B(_1347_),
    .C(_1348_),
    .Y(_1353_));
 sg13g2_nand3_1 _5815_ (.B(net2121),
    .C(_3493_),
    .A(net2571),
    .Y(_1354_));
 sg13g2_or4_1 _5816_ (.A(net2569),
    .B(net2162),
    .C(net2262),
    .D(_3020_),
    .X(_1355_));
 sg13g2_nand4_1 _5817_ (.B(_0604_),
    .C(_1354_),
    .A(net1997),
    .Y(_1356_),
    .D(_1355_));
 sg13g2_a221oi_1 _5818_ (.B2(net2320),
    .C1(_1353_),
    .B1(_1356_),
    .A1(net2307),
    .Y(_1357_),
    .A2(_1352_));
 sg13g2_a21oi_1 _5819_ (.A1(_1351_),
    .A2(_1357_),
    .Y(_1358_),
    .B1(net2393));
 sg13g2_nand2_1 _5820_ (.Y(_1359_),
    .A(net2474),
    .B(_1344_));
 sg13g2_nand2_1 _5821_ (.Y(_1361_),
    .A(net2078),
    .B(_0981_));
 sg13g2_a221oi_1 _5822_ (.B2(net2173),
    .C1(net2403),
    .B1(_1361_),
    .A1(net2217),
    .Y(_1362_),
    .A2(_3130_));
 sg13g2_and4_1 _5823_ (.A(net2545),
    .B(net2152),
    .C(net2078),
    .D(_0981_),
    .X(_1363_));
 sg13g2_nor3_1 _5824_ (.A(net2088),
    .B(net2212),
    .C(_0149_),
    .Y(_1364_));
 sg13g2_nor3_1 _5825_ (.A(_1362_),
    .B(_1363_),
    .C(_1364_),
    .Y(_1365_));
 sg13g2_a21oi_1 _5826_ (.A1(_1359_),
    .A2(_1365_),
    .Y(_1366_),
    .B1(net2194));
 sg13g2_nand3_1 _5827_ (.B(net2088),
    .C(_3077_),
    .A(net2117),
    .Y(_1367_));
 sg13g2_nand3_1 _5828_ (.B(_0604_),
    .C(_1367_),
    .A(net1997),
    .Y(_1368_));
 sg13g2_nand2_1 _5829_ (.Y(_1369_),
    .A(net2289),
    .B(net2211));
 sg13g2_nand3_1 _5830_ (.B(_0288_),
    .C(_1369_),
    .A(net2126),
    .Y(_1370_));
 sg13g2_a21oi_1 _5831_ (.A1(_0978_),
    .A2(_1370_),
    .Y(_1372_),
    .B1(net2467));
 sg13g2_a21oi_1 _5832_ (.A1(net2087),
    .A2(net2234),
    .Y(_1373_),
    .B1(net2148));
 sg13g2_o21ai_1 _5833_ (.B1(net2098),
    .Y(_1374_),
    .A1(net2083),
    .A2(net2235));
 sg13g2_a221oi_1 _5834_ (.B2(net2253),
    .C1(net2145),
    .B1(_3222_),
    .A1(net2087),
    .Y(_1375_),
    .A2(net2234));
 sg13g2_nand2b_1 _5835_ (.Y(_1376_),
    .B(_0604_),
    .A_N(_1375_));
 sg13g2_a221oi_1 _5836_ (.B2(net2545),
    .C1(_1372_),
    .B1(_1376_),
    .A1(net2414),
    .Y(_1377_),
    .A2(_1368_));
 sg13g2_o21ai_1 _5837_ (.B1(_3431_),
    .Y(_1378_),
    .A1(net2199),
    .A2(_1377_));
 sg13g2_nor3_2 _5838_ (.A(_1358_),
    .B(_1366_),
    .C(_1378_),
    .Y(_1379_));
 sg13g2_and2_1 _5839_ (.A(_3295_),
    .B(_0152_),
    .X(_1380_));
 sg13g2_o21ai_1 _5840_ (.B1(net2333),
    .Y(_1381_),
    .A1(_0693_),
    .A2(_1380_));
 sg13g2_o21ai_1 _5841_ (.B1(net2328),
    .Y(_1383_),
    .A1(_0190_),
    .A2(_1155_));
 sg13g2_o21ai_1 _5842_ (.B1(net2590),
    .Y(_1384_),
    .A1(_3246_),
    .A2(_0229_));
 sg13g2_nand2_1 _5843_ (.Y(_1385_),
    .A(net2564),
    .B(_3278_));
 sg13g2_a21oi_1 _5844_ (.A1(_1384_),
    .A2(_1385_),
    .Y(_1386_),
    .B1(net2313));
 sg13g2_a21o_1 _5845_ (.A2(_1385_),
    .A1(_1384_),
    .B1(net2313),
    .X(_1387_));
 sg13g2_nand4_1 _5846_ (.B(_1381_),
    .C(_1383_),
    .A(_0972_),
    .Y(_1388_),
    .D(_1387_));
 sg13g2_nand4_1 _5847_ (.B(_3271_),
    .C(net2196),
    .A(net2589),
    .Y(_1389_),
    .D(_3295_));
 sg13g2_nand4_1 _5848_ (.B(net2260),
    .C(net2432),
    .A(net2154),
    .Y(_1390_),
    .D(net2232));
 sg13g2_nand4_1 _5849_ (.B(net2021),
    .C(net2198),
    .A(net2463),
    .Y(_1391_),
    .D(_1390_));
 sg13g2_nand3_1 _5850_ (.B(_1389_),
    .C(_1391_),
    .A(_3300_),
    .Y(_1392_));
 sg13g2_nand3_1 _5851_ (.B(_3153_),
    .C(_3358_),
    .A(_2778_),
    .Y(_1394_));
 sg13g2_a221oi_1 _5852_ (.B2(net2203),
    .C1(_1392_),
    .B1(_1394_),
    .A1(net2380),
    .Y(_1395_),
    .A2(_1388_));
 sg13g2_nor4_2 _5853_ (.A(net1977),
    .B(_1342_),
    .C(_1379_),
    .Y(_1396_),
    .D(_1395_));
 sg13g2_nor2_1 _5854_ (.A(_3309_),
    .B(_1396_),
    .Y(_1397_));
 sg13g2_a21oi_1 _5855_ (.A1(_1318_),
    .A2(_1397_),
    .Y(_1398_),
    .B1(_3505_));
 sg13g2_a21oi_1 _5856_ (.A1(_1201_),
    .A2(_1398_),
    .Y(_1399_),
    .B1(_1085_));
 sg13g2_a21oi_1 _5857_ (.A1(_1013_),
    .A2(_1399_),
    .Y(_1400_),
    .B1(_0615_));
 sg13g2_o21ai_1 _5858_ (.B1(net2168),
    .Y(_1401_),
    .A1(_3022_),
    .A2(net2065));
 sg13g2_inv_1 _5859_ (.Y(_1402_),
    .A(_1401_));
 sg13g2_nand2_1 _5860_ (.Y(_1403_),
    .A(net2005),
    .B(_1401_));
 sg13g2_nand3_1 _5861_ (.B(net2006),
    .C(_1401_),
    .A(_2724_),
    .Y(_1405_));
 sg13g2_nand3_1 _5862_ (.B(_1855_),
    .C(_2691_),
    .A(net2115),
    .Y(_1406_));
 sg13g2_and4_1 _5863_ (.A(net2571),
    .B(net2005),
    .C(_1401_),
    .D(_1406_),
    .X(_1407_));
 sg13g2_nor3_1 _5864_ (.A(net2166),
    .B(net2263),
    .C(net2219),
    .Y(_1408_));
 sg13g2_a221oi_1 _5865_ (.B2(_0308_),
    .C1(_1408_),
    .B1(_0880_),
    .A1(net2118),
    .Y(_1409_),
    .A2(_0742_));
 sg13g2_or3_1 _5866_ (.A(net2549),
    .B(_1407_),
    .C(_1409_),
    .X(_1410_));
 sg13g2_a21oi_2 _5867_ (.B1(net2077),
    .Y(_1411_),
    .A2(_3081_),
    .A1(net2288));
 sg13g2_o21ai_1 _5868_ (.B1(_0731_),
    .Y(_1412_),
    .A1(net2001),
    .A2(_1411_));
 sg13g2_a221oi_1 _5869_ (.B2(net2445),
    .C1(net2494),
    .B1(_1412_),
    .A1(net2426),
    .Y(_1413_),
    .A2(_1405_));
 sg13g2_a21oi_2 _5870_ (.B1(net2457),
    .Y(_1414_),
    .A2(net2242),
    .A1(net2287));
 sg13g2_nand2_2 _5871_ (.Y(_1416_),
    .A(net2246),
    .B(_1414_));
 sg13g2_a21o_1 _5872_ (.A2(_1414_),
    .A1(net2247),
    .B1(net2118),
    .X(_1417_));
 sg13g2_nor3_1 _5873_ (.A(net2167),
    .B(_1844_),
    .C(_3321_),
    .Y(_1418_));
 sg13g2_nand4_1 _5874_ (.B(_3560_),
    .C(net2005),
    .A(net2494),
    .Y(_1419_),
    .D(_1417_));
 sg13g2_o21ai_1 _5875_ (.B1(net2316),
    .Y(_1420_),
    .A1(_1418_),
    .A2(_1419_));
 sg13g2_o21ai_1 _5876_ (.B1(net2112),
    .Y(_1421_),
    .A1(_3092_),
    .A2(net2054));
 sg13g2_nand2_1 _5877_ (.Y(_1422_),
    .A(_1417_),
    .B(_1421_));
 sg13g2_nand3_1 _5878_ (.B(net2254),
    .C(_2680_),
    .A(net2140),
    .Y(_1423_));
 sg13g2_nor3_2 _5879_ (.A(net2254),
    .B(net2347),
    .C(net2229),
    .Y(_1424_));
 sg13g2_o21ai_1 _5880_ (.B1(net2095),
    .Y(_1425_),
    .A1(net2073),
    .A2(_1424_));
 sg13g2_nand3_1 _5881_ (.B(_1423_),
    .C(_1425_),
    .A(net2011),
    .Y(_1427_));
 sg13g2_a22oi_1 _5882_ (.Y(_1428_),
    .B1(_1427_),
    .B2(net2478),
    .A2(_1422_),
    .A1(net2412));
 sg13g2_a221oi_1 _5883_ (.B2(_1428_),
    .C1(net2396),
    .B1(_1420_),
    .A1(_1410_),
    .Y(_1429_),
    .A2(_1413_));
 sg13g2_nor2_2 _5884_ (.A(net2373),
    .B(net2252),
    .Y(_1430_));
 sg13g2_o21ai_1 _5885_ (.B1(_3076_),
    .Y(_1431_),
    .A1(net2373),
    .A2(net2262));
 sg13g2_nand3_1 _5886_ (.B(net2124),
    .C(_1431_),
    .A(net2596),
    .Y(_1432_));
 sg13g2_nand4_1 _5887_ (.B(net1994),
    .C(net1991),
    .A(net2018),
    .Y(_1433_),
    .D(_1432_));
 sg13g2_mux2_1 _5888_ (.A0(net2068),
    .A1(_0637_),
    .S(net2170),
    .X(_1434_));
 sg13g2_a21oi_2 _5889_ (.B1(net2168),
    .Y(_1435_),
    .A2(_0931_),
    .A1(net2068));
 sg13g2_nand2b_1 _5890_ (.Y(_1436_),
    .B(_0639_),
    .A_N(_1435_));
 sg13g2_a22oi_1 _5891_ (.Y(_1438_),
    .B1(_1436_),
    .B2(_3289_),
    .A2(_1433_),
    .A1(_3459_));
 sg13g2_nor4_2 _5892_ (.A(net2170),
    .B(net2059),
    .C(_3260_),
    .Y(_1439_),
    .D(_3380_));
 sg13g2_nand4_1 _5893_ (.B(net2056),
    .C(_3261_),
    .A(net2115),
    .Y(_1440_),
    .D(_3381_));
 sg13g2_a21oi_1 _5894_ (.A1(_0639_),
    .A2(_1440_),
    .Y(_1441_),
    .B1(net2465));
 sg13g2_a21oi_1 _5895_ (.A1(_0555_),
    .A2(_0639_),
    .Y(_1442_),
    .B1(net2418));
 sg13g2_nand2_1 _5896_ (.Y(_1443_),
    .A(_0898_),
    .B(_1434_));
 sg13g2_a21oi_1 _5897_ (.A1(_0898_),
    .A2(_1434_),
    .Y(_1444_),
    .B1(net2405));
 sg13g2_a21oi_1 _5898_ (.A1(_0514_),
    .A2(_0839_),
    .Y(_1445_),
    .B1(net2434));
 sg13g2_nor4_1 _5899_ (.A(_1441_),
    .B(_1442_),
    .C(_1444_),
    .D(_1445_),
    .Y(_1446_));
 sg13g2_o21ai_1 _5900_ (.B1(_1438_),
    .Y(_1447_),
    .A1(net2200),
    .A2(_1446_));
 sg13g2_o21ai_1 _5901_ (.B1(net1984),
    .Y(_1449_),
    .A1(_1429_),
    .A2(_1447_));
 sg13g2_nor3_2 _5902_ (.A(net2131),
    .B(_3022_),
    .C(_0736_),
    .Y(_1450_));
 sg13g2_nand3_1 _5903_ (.B(_3023_),
    .C(net2053),
    .A(net2170),
    .Y(_1451_));
 sg13g2_nor2_1 _5904_ (.A(_0296_),
    .B(_1450_),
    .Y(_1452_));
 sg13g2_nor2_1 _5905_ (.A(net2555),
    .B(_1450_),
    .Y(_1453_));
 sg13g2_nor2b_1 _5906_ (.A(_0296_),
    .B_N(_1453_),
    .Y(_1454_));
 sg13g2_nor2b_2 _5907_ (.A(_0738_),
    .B_N(_0102_),
    .Y(_1455_));
 sg13g2_nand3_1 _5908_ (.B(_0102_),
    .C(net2052),
    .A(net2175),
    .Y(_1456_));
 sg13g2_o21ai_1 _5909_ (.B1(net2576),
    .Y(_1457_),
    .A1(_0774_),
    .A2(_1455_));
 sg13g2_a21oi_1 _5910_ (.A1(net2598),
    .A2(_0774_),
    .Y(_1458_),
    .B1(net2535));
 sg13g2_nor2_2 _5911_ (.A(_3509_),
    .B(_0451_),
    .Y(_1460_));
 sg13g2_nor2_1 _5912_ (.A(_0296_),
    .B(_1460_),
    .Y(_1461_));
 sg13g2_a221oi_1 _5913_ (.B2(_1461_),
    .C1(net2386),
    .B1(_1458_),
    .A1(_1454_),
    .Y(_1462_),
    .A2(_1457_));
 sg13g2_a21oi_2 _5914_ (.B1(net2597),
    .Y(_1463_),
    .A2(net1993),
    .A1(_0529_));
 sg13g2_nor3_1 _5915_ (.A(net2555),
    .B(_1047_),
    .C(_1463_),
    .Y(_1464_));
 sg13g2_nor2_1 _5916_ (.A(net2576),
    .B(_1053_),
    .Y(_1465_));
 sg13g2_nand3_1 _5917_ (.B(_0302_),
    .C(_1451_),
    .A(net2555),
    .Y(_1466_));
 sg13g2_o21ai_1 _5918_ (.B1(net2384),
    .Y(_1467_),
    .A1(_1465_),
    .A2(_1466_));
 sg13g2_o21ai_1 _5919_ (.B1(net2498),
    .Y(_1468_),
    .A1(_1464_),
    .A2(_1467_));
 sg13g2_or3_1 _5920_ (.A(net2185),
    .B(net2058),
    .C(_0866_),
    .X(_1469_));
 sg13g2_nand3_1 _5921_ (.B(_3101_),
    .C(_3122_),
    .A(net2183),
    .Y(_1471_));
 sg13g2_nand3_1 _5922_ (.B(net1990),
    .C(_1471_),
    .A(_3322_),
    .Y(_1472_));
 sg13g2_nand2_2 _5923_ (.Y(_1473_),
    .A(_2262_),
    .B(net2219));
 sg13g2_nand2_1 _5924_ (.Y(_1474_),
    .A(_1070_),
    .B(net1988));
 sg13g2_a221oi_1 _5925_ (.B2(_0298_),
    .C1(_1474_),
    .B1(_1473_),
    .A1(net2556),
    .Y(_1475_),
    .A2(_1472_));
 sg13g2_a221oi_1 _5926_ (.B2(net2206),
    .C1(net1985),
    .B1(_1475_),
    .A1(_0124_),
    .Y(_1476_),
    .A2(_1452_));
 sg13g2_o21ai_1 _5927_ (.B1(_1476_),
    .Y(_1477_),
    .A1(_1462_),
    .A2(_1468_));
 sg13g2_a21oi_2 _5928_ (.B1(net2126),
    .Y(_1478_),
    .A2(_3102_),
    .A1(net2083));
 sg13g2_o21ai_1 _5929_ (.B1(net2183),
    .Y(_1479_),
    .A1(net2086),
    .A2(_3101_));
 sg13g2_nand3_1 _5930_ (.B(net1989),
    .C(_1479_),
    .A(net1995),
    .Y(_1480_));
 sg13g2_o21ai_1 _5931_ (.B1(net2181),
    .Y(_1482_),
    .A1(net2085),
    .A2(_0101_));
 sg13g2_a22oi_1 _5932_ (.Y(_1483_),
    .B1(_0775_),
    .B2(_1482_),
    .A2(_3450_),
    .A1(_3411_));
 sg13g2_a21oi_2 _5933_ (.B1(net2289),
    .Y(_1484_),
    .A2(net2219),
    .A1(net2234));
 sg13g2_nor2_1 _5934_ (.A(_0773_),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_o21ai_1 _5935_ (.B1(_1482_),
    .Y(_1486_),
    .A1(_0773_),
    .A2(_1484_));
 sg13g2_a221oi_1 _5936_ (.B2(_3419_),
    .C1(_1483_),
    .B1(_1486_),
    .A1(net2307),
    .Y(_1487_),
    .A2(_1480_));
 sg13g2_and2_1 _5937_ (.A(net2399),
    .B(_1487_),
    .X(_1488_));
 sg13g2_nand2_2 _5938_ (.Y(_1489_),
    .A(net2031),
    .B(net1988));
 sg13g2_nand3_1 _5939_ (.B(net1990),
    .C(net1988),
    .A(net2031),
    .Y(_1490_));
 sg13g2_nand2_1 _5940_ (.Y(_1491_),
    .A(net2322),
    .B(_1490_));
 sg13g2_nand3_1 _5941_ (.B(_1487_),
    .C(_1491_),
    .A(net2400),
    .Y(_1493_));
 sg13g2_nand3_1 _5942_ (.B(net1990),
    .C(net1988),
    .A(_1070_),
    .Y(_1494_));
 sg13g2_nor2_2 _5943_ (.A(net2438),
    .B(net2031),
    .Y(_1495_));
 sg13g2_o21ai_1 _5944_ (.B1(net2517),
    .Y(_1496_),
    .A1(_1494_),
    .A2(_1495_));
 sg13g2_a21oi_1 _5945_ (.A1(_3420_),
    .A2(_1472_),
    .Y(_1497_),
    .B1(net2400));
 sg13g2_a21oi_1 _5946_ (.A1(_1496_),
    .A2(_1497_),
    .Y(_1498_),
    .B1(_3432_));
 sg13g2_a21oi_1 _5947_ (.A1(_1493_),
    .A2(_1498_),
    .Y(_1499_),
    .B1(net1977));
 sg13g2_mux2_1 _5948_ (.A0(_2273_),
    .A1(_0866_),
    .S(net2127),
    .X(_1500_));
 sg13g2_o21ai_1 _5949_ (.B1(_3132_),
    .Y(_1501_),
    .A1(net2185),
    .A2(_0866_));
 sg13g2_nor3_2 _5950_ (.A(net2130),
    .B(_3512_),
    .C(_0736_),
    .Y(_1502_));
 sg13g2_mux2_1 _5951_ (.A0(net1987),
    .A1(_1502_),
    .S(net2597),
    .X(_1504_));
 sg13g2_o21ai_1 _5952_ (.B1(_3015_),
    .Y(_1505_),
    .A1(_1501_),
    .A2(_1504_));
 sg13g2_nand4_1 _5953_ (.B(net2004),
    .C(net1995),
    .A(net2017),
    .Y(_1506_),
    .D(_1451_));
 sg13g2_a21oi_1 _5954_ (.A1(net2553),
    .A2(_0755_),
    .Y(_1507_),
    .B1(net2515));
 sg13g2_a221oi_1 _5955_ (.B2(_1500_),
    .C1(net2337),
    .B1(_1451_),
    .A1(_1129_),
    .Y(_1508_),
    .A2(_1294_));
 sg13g2_a221oi_1 _5956_ (.B2(_1486_),
    .C1(_1508_),
    .B1(_1507_),
    .A1(_3410_),
    .Y(_1509_),
    .A2(_1506_));
 sg13g2_a21oi_1 _5957_ (.A1(_1505_),
    .A2(_1509_),
    .Y(_1510_),
    .B1(net2400));
 sg13g2_nand4_1 _5958_ (.B(net2031),
    .C(net1989),
    .A(net2467),
    .Y(_1511_),
    .D(net1988));
 sg13g2_a22oi_1 _5959_ (.Y(_1512_),
    .B1(_1511_),
    .B2(net2205),
    .A2(_1489_),
    .A1(_3289_));
 sg13g2_nand3_1 _5960_ (.B(_3183_),
    .C(_3388_),
    .A(net2481),
    .Y(_1513_));
 sg13g2_nor2_1 _5961_ (.A(_1489_),
    .B(_1513_),
    .Y(_1515_));
 sg13g2_a22oi_1 _5962_ (.Y(_1516_),
    .B1(_1501_),
    .B2(net2197),
    .A2(_1478_),
    .A1(_3459_));
 sg13g2_o21ai_1 _5963_ (.B1(_1516_),
    .Y(_1517_),
    .A1(_1512_),
    .A2(_1515_));
 sg13g2_o21ai_1 _5964_ (.B1(_3374_),
    .Y(_1518_),
    .A1(_1510_),
    .A2(_1517_));
 sg13g2_and4_2 _5965_ (.A(_1449_),
    .B(_1477_),
    .C(_1499_),
    .D(_1518_),
    .X(_1519_));
 sg13g2_a221oi_1 _5966_ (.B2(_0152_),
    .C1(net2199),
    .B1(_3295_),
    .A1(net2432),
    .Y(_1520_),
    .A2(_3263_));
 sg13g2_nor2_1 _5967_ (.A(net1983),
    .B(_1520_),
    .Y(_1521_));
 sg13g2_nor2_1 _5968_ (.A(net1979),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_a221oi_1 _5969_ (.B2(net2095),
    .C1(_3196_),
    .B1(_3147_),
    .A1(_2548_),
    .Y(_1523_),
    .A2(_2625_));
 sg13g2_a21oi_1 _5970_ (.A1(_3298_),
    .A2(_1523_),
    .Y(_1524_),
    .B1(net2542));
 sg13g2_a21oi_1 _5971_ (.A1(_3168_),
    .A2(_0399_),
    .Y(_1526_),
    .B1(net2417));
 sg13g2_and2_1 _5972_ (.A(net2142),
    .B(_0480_),
    .X(_1527_));
 sg13g2_nor3_1 _5973_ (.A(_3170_),
    .B(_3594_),
    .C(_1527_),
    .Y(_1528_));
 sg13g2_o21ai_1 _5974_ (.B1(net2485),
    .Y(_1529_),
    .A1(net2430),
    .A2(_1528_));
 sg13g2_nor3_1 _5975_ (.A(_1524_),
    .B(_1526_),
    .C(_1529_),
    .Y(_1530_));
 sg13g2_nand3_1 _5976_ (.B(net2254),
    .C(_3549_),
    .A(net2142),
    .Y(_1531_));
 sg13g2_and2_1 _5977_ (.A(net2026),
    .B(_1531_),
    .X(_1532_));
 sg13g2_nand2_1 _5978_ (.Y(_1533_),
    .A(net2026),
    .B(_1531_));
 sg13g2_a21oi_1 _5979_ (.A1(net2581),
    .A2(_3235_),
    .Y(_1534_),
    .B1(net2337));
 sg13g2_nand2_1 _5980_ (.Y(_1535_),
    .A(_1532_),
    .B(_1534_));
 sg13g2_a21o_2 _5981_ (.A2(_0170_),
    .A1(net2070),
    .B1(net2142),
    .X(_1537_));
 sg13g2_nand2_2 _5982_ (.Y(_1538_),
    .A(_3393_),
    .B(_0171_));
 sg13g2_and2_1 _5983_ (.A(net2011),
    .B(_1531_),
    .X(_1539_));
 sg13g2_nand3_1 _5984_ (.B(_1537_),
    .C(_1539_),
    .A(net2334),
    .Y(_1540_));
 sg13g2_o21ai_1 _5985_ (.B1(_1540_),
    .Y(_1541_),
    .A1(_1268_),
    .A2(_1535_));
 sg13g2_o21ai_1 _5986_ (.B1(net2390),
    .Y(_1542_),
    .A1(_1530_),
    .A2(_1541_));
 sg13g2_a21oi_1 _5987_ (.A1(_2449_),
    .A2(_3075_),
    .Y(_1543_),
    .B1(net2559));
 sg13g2_a21oi_1 _5988_ (.A1(_2863_),
    .A2(_3075_),
    .Y(_1544_),
    .B1(net2578));
 sg13g2_o21ai_1 _5989_ (.B1(net2319),
    .Y(_1545_),
    .A1(_1543_),
    .A2(_1544_));
 sg13g2_nand3_1 _5990_ (.B(_3195_),
    .C(_0789_),
    .A(_2750_),
    .Y(_1546_));
 sg13g2_mux2_1 _5991_ (.A0(net2240),
    .A1(_2251_),
    .S(net2133),
    .X(_1548_));
 sg13g2_a21oi_1 _5992_ (.A1(_0643_),
    .A2(_1548_),
    .Y(_1549_),
    .B1(_3454_));
 sg13g2_a221oi_1 _5993_ (.B2(net2305),
    .C1(_1549_),
    .B1(_1546_),
    .A1(_3410_),
    .Y(_1550_),
    .A2(_1115_));
 sg13g2_nor2_2 _5994_ (.A(net2490),
    .B(net2341),
    .Y(_1551_));
 sg13g2_nand3_1 _5995_ (.B(net2047),
    .C(_2734_),
    .A(net2051),
    .Y(_1552_));
 sg13g2_a221oi_1 _5996_ (.B2(_1552_),
    .C1(net2388),
    .B1(_1551_),
    .A1(net2309),
    .Y(_1553_),
    .A2(_1115_));
 sg13g2_nand3_1 _5997_ (.B(_1550_),
    .C(_1553_),
    .A(_1545_),
    .Y(_1554_));
 sg13g2_and2_1 _5998_ (.A(net1982),
    .B(_1554_),
    .X(_1555_));
 sg13g2_nor2_1 _5999_ (.A(net2510),
    .B(_0970_),
    .Y(_1556_));
 sg13g2_nor3_1 _6000_ (.A(_3270_),
    .B(_3294_),
    .C(_0560_),
    .Y(_1557_));
 sg13g2_a21oi_2 _6001_ (.B1(net2431),
    .Y(_1559_),
    .A2(_0169_),
    .A1(net2104));
 sg13g2_a221oi_1 _6002_ (.B2(net2024),
    .C1(net2491),
    .B1(_1559_),
    .A1(net2432),
    .Y(_1560_),
    .A2(_1153_));
 sg13g2_or3_1 _6003_ (.A(_1556_),
    .B(_1557_),
    .C(_1560_),
    .X(_1561_));
 sg13g2_nand3_1 _6004_ (.B(net2450),
    .C(_3231_),
    .A(net2107),
    .Y(_1562_));
 sg13g2_mux2_1 _6005_ (.A0(_3227_),
    .A1(_0166_),
    .S(net2102),
    .X(_1563_));
 sg13g2_a21oi_1 _6006_ (.A1(net2526),
    .A2(_1563_),
    .Y(_1564_),
    .B1(_3285_));
 sg13g2_a21oi_1 _6007_ (.A1(_3042_),
    .A2(_1564_),
    .Y(_1565_),
    .B1(net2201));
 sg13g2_o21ai_1 _6008_ (.B1(_3451_),
    .Y(_1566_),
    .A1(net2020),
    .A2(_1163_));
 sg13g2_nand3_1 _6009_ (.B(net2195),
    .C(_0684_),
    .A(net2432),
    .Y(_1567_));
 sg13g2_nand2_1 _6010_ (.Y(_1568_),
    .A(_1566_),
    .B(_1567_));
 sg13g2_a221oi_1 _6011_ (.B2(_1565_),
    .C1(_1568_),
    .B1(_1562_),
    .A1(net2381),
    .Y(_1570_),
    .A2(_1561_));
 sg13g2_a21oi_2 _6012_ (.B1(net2330),
    .Y(_1571_),
    .A2(_3083_),
    .A1(_3045_));
 sg13g2_o21ai_1 _6013_ (.B1(net2473),
    .Y(_1572_),
    .A1(_3238_),
    .A2(_0952_));
 sg13g2_nand3_1 _6014_ (.B(_0655_),
    .C(_1572_),
    .A(_3057_),
    .Y(_1573_));
 sg13g2_a21oi_1 _6015_ (.A1(_3239_),
    .A2(_0953_),
    .Y(_1574_),
    .B1(_3052_));
 sg13g2_a21oi_1 _6016_ (.A1(_3057_),
    .A2(_0655_),
    .Y(_1575_),
    .B1(net2506));
 sg13g2_o21ai_1 _6017_ (.B1(net2585),
    .Y(_1576_),
    .A1(net2045),
    .A2(_0656_));
 sg13g2_nand3b_1 _6018_ (.B(_1576_),
    .C(_3045_),
    .Y(_1577_),
    .A_N(_1189_));
 sg13g2_a221oi_1 _6019_ (.B2(net2338),
    .C1(_1571_),
    .B1(_1577_),
    .A1(net2484),
    .Y(_1578_),
    .A2(_1573_));
 sg13g2_o21ai_1 _6020_ (.B1(net2407),
    .Y(_1579_),
    .A1(_2229_),
    .A2(_3477_));
 sg13g2_o21ai_1 _6021_ (.B1(net2470),
    .Y(_1581_),
    .A1(_3044_),
    .A2(_3093_));
 sg13g2_nand3b_1 _6022_ (.B(_1579_),
    .C(_1581_),
    .Y(_1582_),
    .A_N(_1180_));
 sg13g2_a21oi_1 _6023_ (.A1(_3031_),
    .A2(_1179_),
    .Y(_1583_),
    .B1(net2560));
 sg13g2_a21oi_1 _6024_ (.A1(_3031_),
    .A2(_1179_),
    .Y(_1584_),
    .B1(net2461));
 sg13g2_a21oi_2 _6025_ (.B1(net2520),
    .Y(_1585_),
    .A2(_3075_),
    .A1(_2449_));
 sg13g2_a21oi_1 _6026_ (.A1(_1877_),
    .A2(_3088_),
    .Y(_1586_),
    .B1(net2402));
 sg13g2_or3_1 _6027_ (.A(_1584_),
    .B(_1585_),
    .C(_1586_),
    .X(_1587_));
 sg13g2_a22oi_1 _6028_ (.Y(_1588_),
    .B1(_1587_),
    .B2(net2202),
    .A2(_1582_),
    .A1(net2196));
 sg13g2_o21ai_1 _6029_ (.B1(_1588_),
    .Y(_1589_),
    .A1(net2389),
    .A2(_1578_));
 sg13g2_o21ai_1 _6030_ (.B1(_1522_),
    .Y(_1590_),
    .A1(net1985),
    .A2(_1570_));
 sg13g2_a221oi_1 _6031_ (.B2(_3431_),
    .C1(_1590_),
    .B1(_1589_),
    .A1(_1542_),
    .Y(_1592_),
    .A2(_1555_));
 sg13g2_o21ai_1 _6032_ (.B1(net1976),
    .Y(_1593_),
    .A1(_1519_),
    .A2(_1592_));
 sg13g2_or3_2 _6033_ (.A(net2185),
    .B(_0866_),
    .C(_1484_),
    .X(_1594_));
 sg13g2_nor2b_1 _6034_ (.A(_1489_),
    .B_N(_1594_),
    .Y(_1595_));
 sg13g2_o21ai_1 _6035_ (.B1(net2296),
    .Y(_1596_),
    .A1(net2315),
    .A2(_1595_));
 sg13g2_nor2_2 _6036_ (.A(net2575),
    .B(net1993),
    .Y(_1597_));
 sg13g2_nand3_1 _6037_ (.B(net2242),
    .C(net2074),
    .A(net2181),
    .Y(_1598_));
 sg13g2_nand4_1 _6038_ (.B(net2129),
    .C(net2056),
    .A(net2597),
    .Y(_1599_),
    .D(_0158_));
 sg13g2_nand2_1 _6039_ (.Y(_1600_),
    .A(_1598_),
    .B(_1599_));
 sg13g2_nor3_2 _6040_ (.A(_0776_),
    .B(_1597_),
    .C(_1600_),
    .Y(_1601_));
 sg13g2_o21ai_1 _6041_ (.B1(net2554),
    .Y(_1603_),
    .A1(_0824_),
    .A2(_0838_));
 sg13g2_nand3_1 _6042_ (.B(net2074),
    .C(net2052),
    .A(net2185),
    .Y(_1604_));
 sg13g2_nand3_1 _6043_ (.B(net1989),
    .C(_1604_),
    .A(net2577),
    .Y(_1605_));
 sg13g2_nand4_1 _6044_ (.B(net2031),
    .C(net1989),
    .A(net2598),
    .Y(_1606_),
    .D(net1988));
 sg13g2_nand3_1 _6045_ (.B(_1605_),
    .C(_1606_),
    .A(net2555),
    .Y(_1607_));
 sg13g2_nand2_1 _6046_ (.Y(_1608_),
    .A(_3183_),
    .B(_3393_));
 sg13g2_a21oi_1 _6047_ (.A1(net2481),
    .A2(_1608_),
    .Y(_1609_),
    .B1(net2515));
 sg13g2_a22oi_1 _6048_ (.Y(_1610_),
    .B1(_1607_),
    .B2(_1609_),
    .A2(_1603_),
    .A1(_1601_));
 sg13g2_nor2_1 _6049_ (.A(_1596_),
    .B(_1610_),
    .Y(_1611_));
 sg13g2_o21ai_1 _6050_ (.B1(net2171),
    .Y(_1612_),
    .A1(net2085),
    .A2(_0480_));
 sg13g2_nor2_1 _6051_ (.A(net2594),
    .B(_1612_),
    .Y(_1614_));
 sg13g2_nor2_2 _6052_ (.A(net2265),
    .B(_3421_),
    .Y(_1615_));
 sg13g2_nor2_2 _6053_ (.A(net2169),
    .B(_1615_),
    .Y(_1616_));
 sg13g2_or3_2 _6054_ (.A(net2171),
    .B(net2059),
    .C(_1615_),
    .X(_1617_));
 sg13g2_nand3b_1 _6055_ (.B(_1617_),
    .C(net2514),
    .Y(_1618_),
    .A_N(_0833_));
 sg13g2_o21ai_1 _6056_ (.B1(net2331),
    .Y(_1619_),
    .A1(_1614_),
    .A2(_1618_));
 sg13g2_nand2_1 _6057_ (.Y(_1620_),
    .A(_1612_),
    .B(_1617_));
 sg13g2_nand2b_1 _6058_ (.Y(_1621_),
    .B(_1227_),
    .A_N(_0902_));
 sg13g2_a22oi_1 _6059_ (.Y(_1622_),
    .B1(_1621_),
    .B2(net2446),
    .A2(_1620_),
    .A1(net2427));
 sg13g2_a21oi_1 _6060_ (.A1(_0825_),
    .A2(_0849_),
    .Y(_1623_),
    .B1(net2404));
 sg13g2_a21oi_1 _6061_ (.A1(net1996),
    .A2(_0639_),
    .Y(_1625_),
    .B1(net2468));
 sg13g2_nor3_1 _6062_ (.A(net2515),
    .B(_1623_),
    .C(_1625_),
    .Y(_1626_));
 sg13g2_nand3_1 _6063_ (.B(_0098_),
    .C(_1617_),
    .A(net2030),
    .Y(_1627_));
 sg13g2_nand2_1 _6064_ (.Y(_1628_),
    .A(_0849_),
    .B(_1617_));
 sg13g2_a22oi_1 _6065_ (.Y(_1629_),
    .B1(_1628_),
    .B2(net2428),
    .A2(_1627_),
    .A1(net2448));
 sg13g2_a22oi_1 _6066_ (.Y(_1630_),
    .B1(_1626_),
    .B2(_1629_),
    .A2(_1622_),
    .A1(_1619_));
 sg13g2_nor2_1 _6067_ (.A(net2297),
    .B(_1630_),
    .Y(_1631_));
 sg13g2_o21ai_1 _6068_ (.B1(net2399),
    .Y(_1632_),
    .A1(_1611_),
    .A2(_1631_));
 sg13g2_o21ai_1 _6069_ (.B1(net2575),
    .Y(_1633_),
    .A1(_0546_),
    .A2(_0638_));
 sg13g2_a21oi_1 _6070_ (.A1(net1996),
    .A2(_0639_),
    .Y(_1634_),
    .B1(net2436));
 sg13g2_o21ai_1 _6071_ (.B1(net2516),
    .Y(_1636_),
    .A1(_0806_),
    .A2(_1634_));
 sg13g2_nand2_1 _6072_ (.Y(_1637_),
    .A(_0807_),
    .B(_1451_));
 sg13g2_or2_1 _6073_ (.X(_1638_),
    .B(_1637_),
    .A(_1046_));
 sg13g2_o21ai_1 _6074_ (.B1(net2321),
    .Y(_1639_),
    .A1(_1046_),
    .A2(_1637_));
 sg13g2_nor2_2 _6075_ (.A(net2565),
    .B(_3275_),
    .Y(_1640_));
 sg13g2_o21ai_1 _6076_ (.B1(net2340),
    .Y(_1641_),
    .A1(_1502_),
    .A2(_1640_));
 sg13g2_nand2_1 _6077_ (.Y(_1642_),
    .A(net1993),
    .B(_0807_));
 sg13g2_nor2_1 _6078_ (.A(_0738_),
    .B(_1484_),
    .Y(_1643_));
 sg13g2_a22oi_1 _6079_ (.Y(_1644_),
    .B1(_1643_),
    .B2(net2335),
    .A2(_1642_),
    .A1(net2329));
 sg13g2_nand4_1 _6080_ (.B(_1639_),
    .C(_1641_),
    .A(_1636_),
    .Y(_1645_),
    .D(_1644_));
 sg13g2_a21oi_1 _6081_ (.A1(_3052_),
    .A2(_1608_),
    .Y(_1647_),
    .B1(_1489_));
 sg13g2_o21ai_1 _6082_ (.B1(_1647_),
    .Y(_1648_),
    .A1(_3052_),
    .A2(_1594_));
 sg13g2_a221oi_1 _6083_ (.B2(net1984),
    .C1(_0559_),
    .B1(_1648_),
    .A1(_3300_),
    .Y(_1649_),
    .A2(_1645_));
 sg13g2_inv_1 _6084_ (.Y(_1650_),
    .A(_1649_));
 sg13g2_nor4_1 _6085_ (.A(net2493),
    .B(_3137_),
    .C(_3541_),
    .D(net2009),
    .Y(_1651_));
 sg13g2_or2_1 _6086_ (.X(_1652_),
    .B(_1651_),
    .A(_3419_));
 sg13g2_nor3_2 _6087_ (.A(net2115),
    .B(net2214),
    .C(_3129_),
    .Y(_1653_));
 sg13g2_o21ai_1 _6088_ (.B1(net2410),
    .Y(_1654_),
    .A1(_3594_),
    .A2(_1653_));
 sg13g2_nand2_1 _6089_ (.Y(_1655_),
    .A(_0472_),
    .B(_0931_));
 sg13g2_nand2_1 _6090_ (.Y(_1656_),
    .A(net1997),
    .B(_0625_));
 sg13g2_o21ai_1 _6091_ (.B1(net2441),
    .Y(_1658_),
    .A1(_0450_),
    .A2(_1656_));
 sg13g2_nand2_1 _6092_ (.Y(_1659_),
    .A(_0399_),
    .B(_1277_));
 sg13g2_a22oi_1 _6093_ (.Y(_1660_),
    .B1(_1659_),
    .B2(net2423),
    .A2(_1655_),
    .A1(_3369_));
 sg13g2_nand4_1 _6094_ (.B(_1654_),
    .C(_1658_),
    .A(_1652_),
    .Y(_1661_),
    .D(_1660_));
 sg13g2_nor2b_1 _6095_ (.A(_0919_),
    .B_N(_3200_),
    .Y(_1662_));
 sg13g2_o21ai_1 _6096_ (.B1(net2444),
    .Y(_1663_),
    .A1(_1268_),
    .A2(_1662_));
 sg13g2_nor4_1 _6097_ (.A(_3052_),
    .B(_3392_),
    .C(_3574_),
    .D(_1137_),
    .Y(_1664_));
 sg13g2_nor2_1 _6098_ (.A(net2513),
    .B(_0920_),
    .Y(_1665_));
 sg13g2_nor4_1 _6099_ (.A(_1371_),
    .B(_3392_),
    .C(net2009),
    .D(_0920_),
    .Y(_1666_));
 sg13g2_o21ai_1 _6100_ (.B1(_1663_),
    .Y(_1667_),
    .A1(_1664_),
    .A2(_1666_));
 sg13g2_nand3_1 _6101_ (.B(_1661_),
    .C(_1667_),
    .A(net2295),
    .Y(_1669_));
 sg13g2_nand3_1 _6102_ (.B(_0887_),
    .C(net1991),
    .A(net2049),
    .Y(_1670_));
 sg13g2_nand3_1 _6103_ (.B(_0887_),
    .C(_1039_),
    .A(_3195_),
    .Y(_1671_));
 sg13g2_a221oi_1 _6104_ (.B2(net2471),
    .C1(net2505),
    .B1(_1671_),
    .A1(net2409),
    .Y(_1672_),
    .A2(_1670_));
 sg13g2_a21oi_1 _6105_ (.A1(net2153),
    .A2(net2074),
    .Y(_1673_),
    .B1(net2244));
 sg13g2_nand2_1 _6106_ (.Y(_1674_),
    .A(_3098_),
    .B(_1673_));
 sg13g2_o21ai_1 _6107_ (.B1(_0909_),
    .Y(_1675_),
    .A1(net2251),
    .A2(net2235));
 sg13g2_o21ai_1 _6108_ (.B1(net2330),
    .Y(_1676_),
    .A1(_0183_),
    .A2(_1675_));
 sg13g2_nor2_1 _6109_ (.A(_3514_),
    .B(_3543_),
    .Y(_1677_));
 sg13g2_a21oi_1 _6110_ (.A1(_3098_),
    .A2(_1673_),
    .Y(_1678_),
    .B1(net2564));
 sg13g2_o21ai_1 _6111_ (.B1(net2545),
    .Y(_1680_),
    .A1(_1677_),
    .A2(_1678_));
 sg13g2_a21oi_1 _6112_ (.A1(_1676_),
    .A2(_1680_),
    .Y(_1681_),
    .B1(_1672_));
 sg13g2_nand2_1 _6113_ (.Y(_1682_),
    .A(net2588),
    .B(_1670_));
 sg13g2_o21ai_1 _6114_ (.B1(_0273_),
    .Y(_1683_),
    .A1(net2373),
    .A2(net2258));
 sg13g2_nand2_1 _6115_ (.Y(_1684_),
    .A(net2216),
    .B(net2073));
 sg13g2_a22oi_1 _6116_ (.Y(_1685_),
    .B1(_1684_),
    .B2(_3027_),
    .A2(_1683_),
    .A1(net2022));
 sg13g2_a21oi_1 _6117_ (.A1(_1682_),
    .A2(_1685_),
    .Y(_1686_),
    .B1(net2325));
 sg13g2_o21ai_1 _6118_ (.B1(net2301),
    .Y(_1687_),
    .A1(_1681_),
    .A2(_1686_));
 sg13g2_nand3_1 _6119_ (.B(_1669_),
    .C(_1687_),
    .A(net2398),
    .Y(_1688_));
 sg13g2_o21ai_1 _6120_ (.B1(net2472),
    .Y(_1689_),
    .A1(_3610_),
    .A2(_1656_));
 sg13g2_o21ai_1 _6121_ (.B1(net2096),
    .Y(_1691_),
    .A1(_2680_),
    .A2(net2069));
 sg13g2_a21oi_1 _6122_ (.A1(net2050),
    .A2(_1691_),
    .Y(_1692_),
    .B1(net2584));
 sg13g2_o21ai_1 _6123_ (.B1(_1691_),
    .Y(_1693_),
    .A1(net2584),
    .A2(net2050));
 sg13g2_o21ai_1 _6124_ (.B1(net2097),
    .Y(_1694_),
    .A1(net2077),
    .A2(_3326_));
 sg13g2_inv_1 _6125_ (.Y(_1695_),
    .A(_1694_));
 sg13g2_o21ai_1 _6126_ (.B1(_1694_),
    .Y(_1696_),
    .A1(net2232),
    .A2(_3045_));
 sg13g2_a21oi_1 _6127_ (.A1(net2083),
    .A2(net2346),
    .Y(_1697_),
    .B1(_3266_));
 sg13g2_a21o_1 _6128_ (.A2(_1697_),
    .A1(_3241_),
    .B1(net2504),
    .X(_1698_));
 sg13g2_a221oi_1 _6129_ (.B2(net2409),
    .C1(_1698_),
    .B1(_1696_),
    .A1(net2541),
    .Y(_1699_),
    .A2(_1693_));
 sg13g2_o21ai_1 _6130_ (.B1(net2051),
    .Y(_1700_),
    .A1(_3034_),
    .A2(net2210));
 sg13g2_a21oi_1 _6131_ (.A1(net2525),
    .A2(_1700_),
    .Y(_1702_),
    .B1(net2484));
 sg13g2_and2_1 _6132_ (.A(net2422),
    .B(_0890_),
    .X(_1703_));
 sg13g2_a221oi_1 _6133_ (.B2(net2439),
    .C1(_1703_),
    .B1(_1671_),
    .A1(net2344),
    .Y(_1704_),
    .A2(_1249_));
 sg13g2_a22oi_1 _6134_ (.Y(_1705_),
    .B1(_1702_),
    .B2(_1704_),
    .A2(_1699_),
    .A1(_1689_));
 sg13g2_nand3_1 _6135_ (.B(_3529_),
    .C(net2007),
    .A(_3136_),
    .Y(_1706_));
 sg13g2_o21ai_1 _6136_ (.B1(net2529),
    .Y(_1707_),
    .A1(_3574_),
    .A2(_1706_));
 sg13g2_nand2b_1 _6137_ (.Y(_1708_),
    .B(net2549),
    .A_N(_0899_));
 sg13g2_a21oi_1 _6138_ (.A1(net2242),
    .A2(net2072),
    .Y(_1709_),
    .B1(_2185_));
 sg13g2_a22oi_1 _6139_ (.Y(_1710_),
    .B1(_1709_),
    .B2(_0481_),
    .A2(_1416_),
    .A1(_3358_));
 sg13g2_nand4_1 _6140_ (.B(_1707_),
    .C(_1708_),
    .A(net2513),
    .Y(_1711_),
    .D(_1710_));
 sg13g2_o21ai_1 _6141_ (.B1(net2329),
    .Y(_1713_),
    .A1(net2569),
    .A2(_3261_));
 sg13g2_nor4_1 _6142_ (.A(_3135_),
    .B(_3526_),
    .C(_0740_),
    .D(_1713_),
    .Y(_1714_));
 sg13g2_nor3_2 _6143_ (.A(net2283),
    .B(net2215),
    .C(net2214),
    .Y(_1715_));
 sg13g2_nand3_1 _6144_ (.B(net2030),
    .C(_1227_),
    .A(net2323),
    .Y(_1716_));
 sg13g2_a221oi_1 _6145_ (.B2(_3027_),
    .C1(_1716_),
    .B1(_1715_),
    .A1(net2040),
    .Y(_1717_),
    .A2(_3425_));
 sg13g2_nor3_1 _6146_ (.A(net2302),
    .B(_1714_),
    .C(_1717_),
    .Y(_1718_));
 sg13g2_a221oi_1 _6147_ (.B2(_1718_),
    .C1(net2395),
    .B1(_1711_),
    .A1(net2302),
    .Y(_1719_),
    .A2(_1705_));
 sg13g2_nor2_1 _6148_ (.A(net2036),
    .B(_1719_),
    .Y(_1720_));
 sg13g2_a22oi_1 _6149_ (.Y(_1721_),
    .B1(_1688_),
    .B2(_1720_),
    .A2(_1650_),
    .A1(_1632_));
 sg13g2_a22oi_1 _6150_ (.Y(_1722_),
    .B1(_0288_),
    .B2(net2106),
    .A2(_3176_),
    .A1(net2078));
 sg13g2_nand2_1 _6151_ (.Y(_1724_),
    .A(net2231),
    .B(net2070));
 sg13g2_a22oi_1 _6152_ (.Y(_1725_),
    .B1(_1724_),
    .B2(_1032_),
    .A2(_1722_),
    .A1(net2545));
 sg13g2_a21oi_2 _6153_ (.B1(net2485),
    .Y(_1726_),
    .A2(_3184_),
    .A1(net2408));
 sg13g2_nand2b_1 _6154_ (.Y(_1727_),
    .B(_1726_),
    .A_N(_1725_));
 sg13g2_nand3_1 _6155_ (.B(net2231),
    .C(net2070),
    .A(net2153),
    .Y(_1728_));
 sg13g2_nor3_2 _6156_ (.A(net2104),
    .B(net2238),
    .C(net2075),
    .Y(_1729_));
 sg13g2_nor3_1 _6157_ (.A(net2153),
    .B(net2245),
    .C(_3250_),
    .Y(_1730_));
 sg13g2_nor3_1 _6158_ (.A(net2341),
    .B(_1729_),
    .C(_1730_),
    .Y(_1731_));
 sg13g2_a21o_1 _6159_ (.A2(_1728_),
    .A1(_1559_),
    .B1(_1731_),
    .X(_1732_));
 sg13g2_a22oi_1 _6160_ (.Y(_1733_),
    .B1(_0656_),
    .B2(_1855_),
    .A2(_3352_),
    .A1(net2208));
 sg13g2_a221oi_1 _6161_ (.B2(net2320),
    .C1(net2394),
    .B1(_1733_),
    .A1(net2490),
    .Y(_1735_),
    .A2(_1732_));
 sg13g2_o21ai_1 _6162_ (.B1(net2143),
    .Y(_1736_),
    .A1(_3172_),
    .A2(_3175_));
 sg13g2_o21ai_1 _6163_ (.B1(_3354_),
    .Y(_1737_),
    .A1(_1811_),
    .A2(net2210));
 sg13g2_nand3_1 _6164_ (.B(_1736_),
    .C(_1737_),
    .A(net2441),
    .Y(_1738_));
 sg13g2_nor3_2 _6165_ (.A(net2115),
    .B(_2999_),
    .C(_3101_),
    .Y(_1739_));
 sg13g2_o21ai_1 _6166_ (.B1(net2430),
    .Y(_1740_),
    .A1(_3365_),
    .A2(_1739_));
 sg13g2_nand3_1 _6167_ (.B(_1738_),
    .C(_1740_),
    .A(_3607_),
    .Y(_1741_));
 sg13g2_a21oi_1 _6168_ (.A1(net2565),
    .A2(net2353),
    .Y(_1742_),
    .B1(net2545));
 sg13g2_nand3_1 _6169_ (.B(net2231),
    .C(_3129_),
    .A(net2153),
    .Y(_1743_));
 sg13g2_a221oi_1 _6170_ (.B2(net2104),
    .C1(net2528),
    .B1(_0169_),
    .A1(net2588),
    .Y(_1744_),
    .A2(net2214));
 sg13g2_a221oi_1 _6171_ (.B2(_1744_),
    .C1(net2194),
    .B1(_1743_),
    .A1(_1722_),
    .Y(_1746_),
    .A2(_1742_));
 sg13g2_nand2b_1 _6172_ (.Y(_1747_),
    .B(_3431_),
    .A_N(_1746_));
 sg13g2_a221oi_1 _6173_ (.B2(net2204),
    .C1(_1747_),
    .B1(_1741_),
    .A1(_1727_),
    .Y(_1748_),
    .A2(_1735_));
 sg13g2_a21oi_1 _6174_ (.A1(net2474),
    .A2(_3262_),
    .Y(_1749_),
    .B1(net2491));
 sg13g2_a21o_1 _6175_ (.A2(_1749_),
    .A1(_1562_),
    .B1(_1158_),
    .X(_1750_));
 sg13g2_a221oi_1 _6176_ (.B2(net2393),
    .C1(net1985),
    .B1(_1750_),
    .A1(_3263_),
    .Y(_1751_),
    .A2(_3289_));
 sg13g2_nand3_1 _6177_ (.B(_3271_),
    .C(_3295_),
    .A(net2333),
    .Y(_1752_));
 sg13g2_nand3_1 _6178_ (.B(net2108),
    .C(_3275_),
    .A(net2474),
    .Y(_1753_));
 sg13g2_o21ai_1 _6179_ (.B1(_1753_),
    .Y(_1754_),
    .A1(net2546),
    .A2(_0970_));
 sg13g2_and2_1 _6180_ (.A(net2510),
    .B(_1754_),
    .X(_1755_));
 sg13g2_a22oi_1 _6181_ (.Y(_1757_),
    .B1(_1333_),
    .B2(net2320),
    .A2(_1154_),
    .A1(net2328));
 sg13g2_nand2_1 _6182_ (.Y(_1758_),
    .A(_1752_),
    .B(_1757_));
 sg13g2_o21ai_1 _6183_ (.B1(net2381),
    .Y(_1759_),
    .A1(_1755_),
    .A2(_1758_));
 sg13g2_nand2_1 _6184_ (.Y(_1760_),
    .A(_1751_),
    .B(_1759_));
 sg13g2_o21ai_1 _6185_ (.B1(net2150),
    .Y(_1761_),
    .A1(net2241),
    .A2(_2912_));
 sg13g2_a21oi_2 _6186_ (.B1(net2101),
    .Y(_1762_),
    .A2(net2075),
    .A1(net2244));
 sg13g2_o21ai_1 _6187_ (.B1(net2424),
    .Y(_1763_),
    .A1(_0209_),
    .A2(_1762_));
 sg13g2_nand2_1 _6188_ (.Y(_1764_),
    .A(_0227_),
    .B(_1761_));
 sg13g2_o21ai_1 _6189_ (.B1(net2442),
    .Y(_1765_),
    .A1(_0226_),
    .A2(_1762_));
 sg13g2_a21o_1 _6190_ (.A2(_1336_),
    .A1(_3053_),
    .B1(net2463),
    .X(_1766_));
 sg13g2_nand3_1 _6191_ (.B(_1765_),
    .C(_1766_),
    .A(_1763_),
    .Y(_1768_));
 sg13g2_o21ai_1 _6192_ (.B1(net2409),
    .Y(_1769_),
    .A1(_0209_),
    .A2(_1762_));
 sg13g2_nand2b_1 _6193_ (.Y(_1770_),
    .B(_1769_),
    .A_N(_1768_));
 sg13g2_a21oi_1 _6194_ (.A1(_3271_),
    .A2(_1329_),
    .Y(_1771_),
    .B1(net2507));
 sg13g2_nand2_1 _6195_ (.Y(_1772_),
    .A(net2431),
    .B(_1329_));
 sg13g2_nand2_1 _6196_ (.Y(_1773_),
    .A(_1771_),
    .B(_1772_));
 sg13g2_nor2_1 _6197_ (.A(_3411_),
    .B(_0783_),
    .Y(_1774_));
 sg13g2_a221oi_1 _6198_ (.B2(_0948_),
    .C1(net2391),
    .B1(_1774_),
    .A1(_3419_),
    .Y(_1775_),
    .A2(_1322_));
 sg13g2_a21oi_1 _6199_ (.A1(net2024),
    .A2(_0230_),
    .Y(_1776_),
    .B1(net2527));
 sg13g2_a21oi_1 _6200_ (.A1(net2527),
    .A2(_1764_),
    .Y(_1777_),
    .B1(_1776_));
 sg13g2_o21ai_1 _6201_ (.B1(net1984),
    .Y(_1779_),
    .A1(net2199),
    .A2(_1777_));
 sg13g2_a221oi_1 _6202_ (.B2(_1775_),
    .C1(_1779_),
    .B1(_1773_),
    .A1(net2195),
    .Y(_1780_),
    .A2(_1770_));
 sg13g2_nor3_1 _6203_ (.A(net1977),
    .B(_1748_),
    .C(_1780_),
    .Y(_1781_));
 sg13g2_a21oi_1 _6204_ (.A1(_1760_),
    .A2(_1781_),
    .Y(_1782_),
    .B1(net1976));
 sg13g2_o21ai_1 _6205_ (.B1(_1782_),
    .Y(_1783_),
    .A1(net1980),
    .A2(_1721_));
 sg13g2_and2_1 _6206_ (.A(_3506_),
    .B(_1593_),
    .X(_1784_));
 sg13g2_o21ai_1 _6207_ (.B1(net2446),
    .Y(_1785_),
    .A1(_3574_),
    .A2(_1403_));
 sg13g2_o21ai_1 _6208_ (.B1(_1227_),
    .Y(_1786_),
    .A1(_0156_),
    .A2(_0738_));
 sg13g2_nand2b_1 _6209_ (.Y(_1787_),
    .B(_1287_),
    .A_N(_0740_));
 sg13g2_a221oi_1 _6210_ (.B2(net2412),
    .C1(net2512),
    .B1(_1787_),
    .A1(net2478),
    .Y(_1788_),
    .A2(_1786_));
 sg13g2_nand3_1 _6211_ (.B(net2005),
    .C(net1994),
    .A(_0242_),
    .Y(_1790_));
 sg13g2_nand2_1 _6212_ (.Y(_1791_),
    .A(net2426),
    .B(_1790_));
 sg13g2_nand3_1 _6213_ (.B(_1788_),
    .C(_1791_),
    .A(_1785_),
    .Y(_1792_));
 sg13g2_nand2_1 _6214_ (.Y(_1793_),
    .A(net2230),
    .B(_1254_));
 sg13g2_nand2_1 _6215_ (.Y(_1794_),
    .A(net2083),
    .B(_2592_));
 sg13g2_o21ai_1 _6216_ (.B1(net2513),
    .Y(_1795_),
    .A1(net2466),
    .A2(_3144_));
 sg13g2_a221oi_1 _6217_ (.B2(_3241_),
    .C1(_1795_),
    .B1(_1794_),
    .A1(_1032_),
    .Y(_1796_),
    .A2(_1793_));
 sg13g2_nor2_1 _6218_ (.A(net2434),
    .B(_3392_),
    .Y(_1797_));
 sg13g2_a22oi_1 _6219_ (.Y(_1798_),
    .B1(_1797_),
    .B2(_0898_),
    .A2(_0899_),
    .A1(net2434));
 sg13g2_nand2b_1 _6220_ (.Y(_1799_),
    .B(_1796_),
    .A_N(_1798_));
 sg13g2_nand3_1 _6221_ (.B(_2548_),
    .C(_0947_),
    .A(net2142),
    .Y(_1801_));
 sg13g2_nand3_1 _6222_ (.B(_1277_),
    .C(_1801_),
    .A(net2581),
    .Y(_1802_));
 sg13g2_nand4_1 _6223_ (.B(net2044),
    .C(net1997),
    .A(net2561),
    .Y(_1803_),
    .D(_0625_));
 sg13g2_nand3_1 _6224_ (.B(_1802_),
    .C(_1803_),
    .A(net2542),
    .Y(_1804_));
 sg13g2_nand3_1 _6225_ (.B(_0932_),
    .C(_1531_),
    .A(net2027),
    .Y(_1805_));
 sg13g2_a22oi_1 _6226_ (.Y(_1806_),
    .B1(_0318_),
    .B2(_0472_),
    .A2(_3540_),
    .A1(net2158));
 sg13g2_a22oi_1 _6227_ (.Y(_1807_),
    .B1(_1806_),
    .B2(net2410),
    .A2(_1805_),
    .A1(net2476));
 sg13g2_a21oi_1 _6228_ (.A1(_1804_),
    .A2(_1807_),
    .Y(_1808_),
    .B1(net2493));
 sg13g2_nand4_1 _6229_ (.B(net2593),
    .C(net2548),
    .A(net2493),
    .Y(_1809_),
    .D(_1269_));
 sg13g2_o21ai_1 _6230_ (.B1(net2310),
    .Y(_1810_),
    .A1(_0920_),
    .A2(_1268_));
 sg13g2_nand2_1 _6231_ (.Y(_1812_),
    .A(_0398_),
    .B(_0952_));
 sg13g2_a22oi_1 _6232_ (.Y(_1813_),
    .B1(_1416_),
    .B2(net2040),
    .A2(_0619_),
    .A1(_3027_));
 sg13g2_a21o_1 _6233_ (.A2(_1813_),
    .A1(_1812_),
    .B1(net2316),
    .X(_1814_));
 sg13g2_nand3_1 _6234_ (.B(_1810_),
    .C(_1814_),
    .A(_1809_),
    .Y(_1815_));
 sg13g2_o21ai_1 _6235_ (.B1(net2395),
    .Y(_1816_),
    .A1(_1808_),
    .A2(_1815_));
 sg13g2_nand3_1 _6236_ (.B(_1792_),
    .C(_1799_),
    .A(net2382),
    .Y(_1817_));
 sg13g2_nand3_1 _6237_ (.B(_1816_),
    .C(_1817_),
    .A(_3431_),
    .Y(_1818_));
 sg13g2_nand2_2 _6238_ (.Y(_1819_),
    .A(net2282),
    .B(_3510_));
 sg13g2_nand2_1 _6239_ (.Y(_1820_),
    .A(net2093),
    .B(_1819_));
 sg13g2_and2_2 _6240_ (.A(net2103),
    .B(_1819_),
    .X(_1821_));
 sg13g2_nor2_1 _6241_ (.A(net2585),
    .B(_1820_),
    .Y(_1823_));
 sg13g2_o21ai_1 _6242_ (.B1(_3031_),
    .Y(_1824_),
    .A1(net2560),
    .A2(_0230_));
 sg13g2_o21ai_1 _6243_ (.B1(net2544),
    .Y(_1825_),
    .A1(_1823_),
    .A2(_1824_));
 sg13g2_a21oi_1 _6244_ (.A1(net2042),
    .A2(net1991),
    .Y(_1826_),
    .B1(net2417));
 sg13g2_a221oi_1 _6245_ (.B2(net2439),
    .C1(_1826_),
    .B1(_1242_),
    .A1(net2539),
    .Y(_1827_),
    .A2(_0886_));
 sg13g2_a22oi_1 _6246_ (.Y(_1828_),
    .B1(_1827_),
    .B2(_1672_),
    .A2(_1825_),
    .A1(_1676_));
 sg13g2_o21ai_1 _6247_ (.B1(net2522),
    .Y(_1829_),
    .A1(_3253_),
    .A2(_1411_));
 sg13g2_nor3_1 _6248_ (.A(_3610_),
    .B(_1247_),
    .C(_1829_),
    .Y(_1830_));
 sg13g2_o21ai_1 _6249_ (.B1(net2485),
    .Y(_1831_),
    .A1(_1249_),
    .A2(_1253_));
 sg13g2_a221oi_1 _6250_ (.B2(net2562),
    .C1(net2523),
    .B1(_0300_),
    .A1(net2097),
    .Y(_1832_),
    .A2(_3145_));
 sg13g2_a21oi_1 _6251_ (.A1(net1991),
    .A2(_1832_),
    .Y(_1834_),
    .B1(net2486));
 sg13g2_a221oi_1 _6252_ (.B2(_1834_),
    .C1(net2389),
    .B1(_1251_),
    .A1(_2086_),
    .Y(_1835_),
    .A2(_0560_));
 sg13g2_o21ai_1 _6253_ (.B1(_1835_),
    .Y(_1836_),
    .A1(_1830_),
    .A2(_1831_));
 sg13g2_o21ai_1 _6254_ (.B1(_1836_),
    .Y(_1837_),
    .A1(net2380),
    .A2(_1828_));
 sg13g2_nor2_2 _6255_ (.A(net2354),
    .B(net2068),
    .Y(_1838_));
 sg13g2_nor3_1 _6256_ (.A(net2129),
    .B(net2354),
    .C(net2068),
    .Y(_1839_));
 sg13g2_nor4_1 _6257_ (.A(net2536),
    .B(_3133_),
    .C(_0546_),
    .D(_1839_),
    .Y(_1840_));
 sg13g2_nor4_1 _6258_ (.A(net2557),
    .B(_3335_),
    .C(_3433_),
    .D(_1502_),
    .Y(_1841_));
 sg13g2_a22oi_1 _6259_ (.Y(_1842_),
    .B1(_3274_),
    .B2(net2414),
    .A2(_3141_),
    .A1(net2449));
 sg13g2_o21ai_1 _6260_ (.B1(_1842_),
    .Y(_1843_),
    .A1(_1840_),
    .A2(_1841_));
 sg13g2_nor3_1 _6261_ (.A(_0751_),
    .B(_1203_),
    .C(_1226_),
    .Y(_1845_));
 sg13g2_o21ai_1 _6262_ (.B1(net2385),
    .Y(_1846_),
    .A1(net2327),
    .A2(_1845_));
 sg13g2_a221oi_1 _6263_ (.B2(net2516),
    .C1(_1846_),
    .B1(_1843_),
    .A1(net2321),
    .Y(_1847_),
    .A2(_1638_));
 sg13g2_nand2b_1 _6264_ (.Y(_1848_),
    .B(_1227_),
    .A_N(_1653_));
 sg13g2_nand3_1 _6265_ (.B(net2019),
    .C(_1612_),
    .A(net2025),
    .Y(_1849_));
 sg13g2_a21oi_1 _6266_ (.A1(_0141_),
    .A2(_1617_),
    .Y(_1850_),
    .B1(net2550));
 sg13g2_o21ai_1 _6267_ (.B1(net2207),
    .Y(_1851_),
    .A1(net2465),
    .A2(net2211));
 sg13g2_or3_1 _6268_ (.A(_1495_),
    .B(_1850_),
    .C(_1851_),
    .X(_1852_));
 sg13g2_a221oi_1 _6269_ (.B2(net2426),
    .C1(_1852_),
    .B1(_1849_),
    .A1(net2446),
    .Y(_1853_),
    .A2(_1848_));
 sg13g2_nand2_1 _6270_ (.Y(_1854_),
    .A(net2554),
    .B(_1628_));
 sg13g2_and3_1 _6271_ (.X(_1856_),
    .A(net2197),
    .B(_1223_),
    .C(_1854_));
 sg13g2_or4_2 _6272_ (.A(net2297),
    .B(_1847_),
    .C(_1853_),
    .D(_1856_),
    .X(_1857_));
 sg13g2_nand3_1 _6273_ (.B(_1303_),
    .C(_1599_),
    .A(net1996),
    .Y(_1858_));
 sg13g2_nand3_1 _6274_ (.B(_0775_),
    .C(_1077_),
    .A(net2414),
    .Y(_1859_));
 sg13g2_a21oi_1 _6275_ (.A1(_1858_),
    .A2(_1859_),
    .Y(_1860_),
    .B1(net2200));
 sg13g2_nand4_1 _6276_ (.B(_3410_),
    .C(_0825_),
    .A(net2399),
    .Y(_1861_),
    .D(_0849_));
 sg13g2_nand3_1 _6277_ (.B(net2289),
    .C(_3511_),
    .A(net2126),
    .Y(_1862_));
 sg13g2_nand3_1 _6278_ (.B(net1992),
    .C(_1862_),
    .A(_0725_),
    .Y(_1863_));
 sg13g2_o21ai_1 _6279_ (.B1(net2296),
    .Y(_1864_),
    .A1(_0110_),
    .A2(_1863_));
 sg13g2_nor2b_1 _6280_ (.A(_1864_),
    .B_N(_1861_),
    .Y(_1865_));
 sg13g2_nand3_1 _6281_ (.B(net2056),
    .C(_1819_),
    .A(net2128),
    .Y(_1867_));
 sg13g2_nand2_1 _6282_ (.Y(_1868_),
    .A(net2553),
    .B(_1867_));
 sg13g2_o21ai_1 _6283_ (.B1(net2404),
    .Y(_1869_),
    .A1(_1312_),
    .A2(_1868_));
 sg13g2_nand2_1 _6284_ (.Y(_1870_),
    .A(net1992),
    .B(_1867_));
 sg13g2_a21oi_1 _6285_ (.A1(net2437),
    .A2(_1870_),
    .Y(_1871_),
    .B1(net2192));
 sg13g2_nand2_1 _6286_ (.Y(_1872_),
    .A(net2315),
    .B(_1863_));
 sg13g2_a21oi_1 _6287_ (.A1(net1992),
    .A2(_1867_),
    .Y(_1873_),
    .B1(net2315));
 sg13g2_o21ai_1 _6288_ (.B1(net2383),
    .Y(_1874_),
    .A1(_3062_),
    .A2(_3314_));
 sg13g2_nor2_1 _6289_ (.A(_1873_),
    .B(_1874_),
    .Y(_1875_));
 sg13g2_a221oi_1 _6290_ (.B2(_1875_),
    .C1(_1860_),
    .B1(_1872_),
    .A1(_1869_),
    .Y(_1876_),
    .A2(_1871_));
 sg13g2_a21oi_1 _6291_ (.A1(_1865_),
    .A2(_1876_),
    .Y(_1878_),
    .B1(net2039));
 sg13g2_a221oi_1 _6292_ (.B2(_1878_),
    .C1(net1978),
    .B1(_1857_),
    .A1(net1982),
    .Y(_1879_),
    .A2(_1837_));
 sg13g2_o21ai_1 _6293_ (.B1(_1855_),
    .Y(_1880_),
    .A1(_2394_),
    .A2(_3469_));
 sg13g2_a21oi_1 _6294_ (.A1(net2352),
    .A2(net2069),
    .Y(_1881_),
    .B1(_0157_));
 sg13g2_nor2_1 _6295_ (.A(net2588),
    .B(_3151_),
    .Y(_1882_));
 sg13g2_a221oi_1 _6296_ (.B2(_3352_),
    .C1(net2314),
    .B1(_1882_),
    .A1(net2041),
    .Y(_1883_),
    .A2(_1881_));
 sg13g2_a221oi_1 _6297_ (.B2(net2569),
    .C1(_3531_),
    .B1(_0866_),
    .A1(net2115),
    .Y(_1884_),
    .A2(net2248));
 sg13g2_a22oi_1 _6298_ (.Y(_1885_),
    .B1(_1884_),
    .B2(net2545),
    .A2(_0485_),
    .A1(_1877_));
 sg13g2_o21ai_1 _6299_ (.B1(net2588),
    .Y(_1886_),
    .A1(_0473_),
    .A2(_1729_));
 sg13g2_a221oi_1 _6300_ (.B2(net2033),
    .C1(net2325),
    .B1(_0729_),
    .A1(net2022),
    .Y(_1887_),
    .A2(_0589_));
 sg13g2_a22oi_1 _6301_ (.Y(_1889_),
    .B1(_1886_),
    .B2(_1887_),
    .A2(_1883_),
    .A1(_1880_));
 sg13g2_o21ai_1 _6302_ (.B1(_1889_),
    .Y(_1890_),
    .A1(net2490),
    .A2(_1885_));
 sg13g2_nor2_1 _6303_ (.A(_3182_),
    .B(_3397_),
    .Y(_1891_));
 sg13g2_nor3_1 _6304_ (.A(net2128),
    .B(_0561_),
    .C(_1891_),
    .Y(_1892_));
 sg13g2_nor2_1 _6305_ (.A(net1981),
    .B(_1892_),
    .Y(_1893_));
 sg13g2_a221oi_1 _6306_ (.B2(net2108),
    .C1(_3256_),
    .B1(_3275_),
    .A1(net2565),
    .Y(_1894_),
    .A2(_3269_));
 sg13g2_nor2_1 _6307_ (.A(net2326),
    .B(_1894_),
    .Y(_1895_));
 sg13g2_nor4_1 _6308_ (.A(_1386_),
    .B(_1392_),
    .C(_1755_),
    .D(_1895_),
    .Y(_1896_));
 sg13g2_a22oi_1 _6309_ (.Y(_1897_),
    .B1(_1896_),
    .B2(_1381_),
    .A2(_1893_),
    .A1(_1890_));
 sg13g2_nor2_1 _6310_ (.A(net2393),
    .B(_1897_),
    .Y(_1898_));
 sg13g2_o21ai_1 _6311_ (.B1(net2506),
    .Y(_1900_),
    .A1(_0219_),
    .A2(_1324_));
 sg13g2_nand2_1 _6312_ (.Y(_1901_),
    .A(net2586),
    .B(_1329_));
 sg13g2_a21oi_1 _6313_ (.A1(_0784_),
    .A2(_1901_),
    .Y(_1902_),
    .B1(net2326));
 sg13g2_nand2_2 _6314_ (.Y(_1903_),
    .A(_0216_),
    .B(_0221_));
 sg13g2_o21ai_1 _6315_ (.B1(_1903_),
    .Y(_1904_),
    .A1(_3420_),
    .A2(_1322_));
 sg13g2_a22oi_1 _6316_ (.Y(_1905_),
    .B1(_3171_),
    .B2(net2093),
    .A2(net2041),
    .A1(_3021_));
 sg13g2_nor2_1 _6317_ (.A(net2313),
    .B(_1905_),
    .Y(_1906_));
 sg13g2_nor3_1 _6318_ (.A(_1902_),
    .B(_1904_),
    .C(_1906_),
    .Y(_1907_));
 sg13g2_a21oi_1 _6319_ (.A1(_1900_),
    .A2(_1907_),
    .Y(_1908_),
    .B1(net2391));
 sg13g2_nand2_1 _6320_ (.Y(_1909_),
    .A(_0208_),
    .B(_1336_));
 sg13g2_a22oi_1 _6321_ (.Y(_1911_),
    .B1(_1909_),
    .B2(net2409),
    .A2(_1323_),
    .A1(net2473));
 sg13g2_nand3_1 _6322_ (.B(_1765_),
    .C(_1911_),
    .A(_1763_),
    .Y(_1912_));
 sg13g2_and2_1 _6323_ (.A(net2195),
    .B(_1912_),
    .X(_1913_));
 sg13g2_nand2_1 _6324_ (.Y(_1914_),
    .A(net2544),
    .B(_3249_));
 sg13g2_nor2_1 _6325_ (.A(_0965_),
    .B(_1914_),
    .Y(_1915_));
 sg13g2_nor3_1 _6326_ (.A(net2402),
    .B(net2020),
    .C(_0229_),
    .Y(_1916_));
 sg13g2_o21ai_1 _6327_ (.B1(net2203),
    .Y(_1917_),
    .A1(net2462),
    .A2(_0961_));
 sg13g2_nor3_1 _6328_ (.A(_1915_),
    .B(_1916_),
    .C(_1917_),
    .Y(_1918_));
 sg13g2_nor4_2 _6329_ (.A(net1983),
    .B(_1908_),
    .C(_1913_),
    .Y(_1919_),
    .D(_1918_));
 sg13g2_a21oi_1 _6330_ (.A1(net2022),
    .A2(_0589_),
    .Y(_1920_),
    .B1(_1888_));
 sg13g2_nand2b_1 _6331_ (.Y(_1922_),
    .B(net2543),
    .A_N(_1920_));
 sg13g2_o21ai_1 _6332_ (.B1(_3297_),
    .Y(_1923_),
    .A1(net2064),
    .A2(_0554_));
 sg13g2_a21oi_1 _6333_ (.A1(net2265),
    .A2(net2216),
    .Y(_1924_),
    .B1(net2122));
 sg13g2_a22oi_1 _6334_ (.Y(_1925_),
    .B1(_1924_),
    .B2(net2230),
    .A2(net2213),
    .A1(net2413));
 sg13g2_and3_2 _6335_ (.X(_1926_),
    .A(net2495),
    .B(_1923_),
    .C(_1925_));
 sg13g2_nor4_2 _6336_ (.A(net2522),
    .B(net2095),
    .C(_3172_),
    .Y(_1927_),
    .D(_1838_));
 sg13g2_and2_1 _6337_ (.A(net2523),
    .B(_1739_),
    .X(_1928_));
 sg13g2_o21ai_1 _6338_ (.B1(net2461),
    .Y(_1929_),
    .A1(_1375_),
    .A2(_1928_));
 sg13g2_a221oi_1 _6339_ (.B2(net2161),
    .C1(net2466),
    .B1(_1254_),
    .A1(_2647_),
    .Y(_1930_),
    .A2(net2215));
 sg13g2_nor3_1 _6340_ (.A(net2496),
    .B(_1927_),
    .C(_1930_),
    .Y(_1931_));
 sg13g2_a22oi_1 _6341_ (.Y(_1933_),
    .B1(_1929_),
    .B2(_1931_),
    .A2(_1926_),
    .A1(_1922_));
 sg13g2_or2_1 _6342_ (.X(_1934_),
    .B(_1749_),
    .A(_1392_));
 sg13g2_o21ai_1 _6343_ (.B1(_1934_),
    .Y(_1935_),
    .A1(net1981),
    .A2(_1933_));
 sg13g2_and2_1 _6344_ (.A(net2393),
    .B(_1935_),
    .X(_1936_));
 sg13g2_or4_1 _6345_ (.A(net1977),
    .B(_1898_),
    .C(_1919_),
    .D(_1936_),
    .X(_1937_));
 sg13g2_a21oi_1 _6346_ (.A1(_1818_),
    .A2(_1879_),
    .Y(_1938_),
    .B1(net1976));
 sg13g2_o21ai_1 _6347_ (.B1(net2534),
    .Y(_1939_),
    .A1(_1046_),
    .A2(_1463_));
 sg13g2_a21oi_1 _6348_ (.A1(_0302_),
    .A2(_1049_),
    .Y(_1940_),
    .B1(net2436));
 sg13g2_a21oi_1 _6349_ (.A1(_0791_),
    .A2(_1053_),
    .Y(_1941_),
    .B1(net2418));
 sg13g2_nor3_1 _6350_ (.A(net2519),
    .B(_1940_),
    .C(_1941_),
    .Y(_1942_));
 sg13g2_nand2_1 _6351_ (.Y(_1944_),
    .A(net2519),
    .B(_1049_));
 sg13g2_a21oi_1 _6352_ (.A1(net2436),
    .A2(_0324_),
    .Y(_1945_),
    .B1(_1944_));
 sg13g2_a221oi_1 _6353_ (.B2(_0297_),
    .C1(net2297),
    .B1(_1945_),
    .A1(_1939_),
    .Y(_1946_),
    .A2(_1942_));
 sg13g2_a21oi_1 _6354_ (.A1(net2227),
    .A2(_3320_),
    .Y(_1947_),
    .B1(_1021_));
 sg13g2_a21oi_1 _6355_ (.A1(net2595),
    .A2(_1537_),
    .Y(_1948_),
    .B1(_1947_));
 sg13g2_nor3_1 _6356_ (.A(net2418),
    .B(net2054),
    .C(_0554_),
    .Y(_1949_));
 sg13g2_and2_1 _6357_ (.A(_1866_),
    .B(_0102_),
    .X(_1950_));
 sg13g2_a221oi_1 _6358_ (.B2(_1950_),
    .C1(_1949_),
    .B1(net2445),
    .A1(net2465),
    .Y(_1951_),
    .A2(net2166));
 sg13g2_o21ai_1 _6359_ (.B1(_1951_),
    .Y(_1952_),
    .A1(net2549),
    .A2(_1948_));
 sg13g2_nand3_1 _6360_ (.B(_1417_),
    .C(_1952_),
    .A(net2494),
    .Y(_1953_));
 sg13g2_a221oi_1 _6361_ (.B2(_3081_),
    .C1(net2054),
    .B1(net2286),
    .A1(_1129_),
    .Y(_1955_),
    .A2(_1294_));
 sg13g2_nor2_1 _6362_ (.A(net2572),
    .B(net2054),
    .Y(_1956_));
 sg13g2_nor4_1 _6363_ (.A(net2573),
    .B(_3007_),
    .C(net2054),
    .D(_0100_),
    .Y(_1957_));
 sg13g2_nor3_1 _6364_ (.A(_0149_),
    .B(_1955_),
    .C(_1957_),
    .Y(_1958_));
 sg13g2_nor4_1 _6365_ (.A(net2170),
    .B(net2244),
    .C(net2405),
    .D(_2982_),
    .Y(_1959_));
 sg13g2_nor2_1 _6366_ (.A(net2530),
    .B(net1994),
    .Y(_1960_));
 sg13g2_nand2_1 _6367_ (.Y(_1961_),
    .A(net2119),
    .B(_1950_));
 sg13g2_a21oi_1 _6368_ (.A1(_1414_),
    .A2(_1924_),
    .Y(_1962_),
    .B1(net2465));
 sg13g2_nor4_1 _6369_ (.A(net2495),
    .B(_1958_),
    .C(_1959_),
    .D(_1960_),
    .Y(_1963_));
 sg13g2_a22oi_1 _6370_ (.Y(_1964_),
    .B1(_1961_),
    .B2(_1962_),
    .A2(_1403_),
    .A1(net2413));
 sg13g2_a21oi_2 _6371_ (.B1(net2303),
    .Y(_1966_),
    .A2(_1964_),
    .A1(_1963_));
 sg13g2_a21o_1 _6372_ (.A2(_1966_),
    .A1(_1953_),
    .B1(_1946_),
    .X(_1967_));
 sg13g2_nand3_1 _6373_ (.B(net2018),
    .C(net1994),
    .A(net2025),
    .Y(_1968_));
 sg13g2_nand2_1 _6374_ (.Y(_1969_),
    .A(net2312),
    .B(_1968_));
 sg13g2_nor3_1 _6375_ (.A(_3040_),
    .B(_3380_),
    .C(_1432_),
    .Y(_1970_));
 sg13g2_nand2_1 _6376_ (.Y(_1971_),
    .A(net2337),
    .B(net2308));
 sg13g2_a221oi_1 _6377_ (.B2(_1971_),
    .C1(_1970_),
    .B1(_1436_),
    .A1(_3453_),
    .Y(_1972_),
    .A2(_0764_));
 sg13g2_nand3_1 _6378_ (.B(_0093_),
    .C(net1991),
    .A(net2018),
    .Y(_1973_));
 sg13g2_o21ai_1 _6379_ (.B1(_3061_),
    .Y(_1974_),
    .A1(_3133_),
    .A2(_1973_));
 sg13g2_nand4_1 _6380_ (.B(_1969_),
    .C(_1972_),
    .A(net2298),
    .Y(_1975_),
    .D(_1974_));
 sg13g2_nand2_1 _6381_ (.Y(_1977_),
    .A(net2412),
    .B(_1439_));
 sg13g2_a22oi_1 _6382_ (.Y(_1978_),
    .B1(_1443_),
    .B2(net2427),
    .A2(_0787_),
    .A1(net2445));
 sg13g2_nand4_1 _6383_ (.B(net2013),
    .C(net2003),
    .A(net2428),
    .Y(_1979_),
    .D(_1068_));
 sg13g2_o21ai_1 _6384_ (.B1(net2497),
    .Y(_1980_),
    .A1(_0774_),
    .A2(_1067_));
 sg13g2_o21ai_1 _6385_ (.B1(_1979_),
    .Y(_1981_),
    .A1(net2437),
    .A2(_1072_));
 sg13g2_a21o_1 _6386_ (.A2(_1980_),
    .A1(net2327),
    .B1(_1981_),
    .X(_1982_));
 sg13g2_o21ai_1 _6387_ (.B1(net2518),
    .Y(_1983_),
    .A1(_0329_),
    .A2(_1058_));
 sg13g2_o21ai_1 _6388_ (.B1(_1867_),
    .Y(_1984_),
    .A1(net2024),
    .A2(_3312_));
 sg13g2_a22oi_1 _6389_ (.Y(_1985_),
    .B1(_1984_),
    .B2(net2332),
    .A2(_3226_),
    .A1(net2311));
 sg13g2_nand4_1 _6390_ (.B(_1982_),
    .C(_1983_),
    .A(net2303),
    .Y(_1986_),
    .D(_1985_));
 sg13g2_a21oi_1 _6391_ (.A1(_1977_),
    .A2(_1978_),
    .Y(_1988_),
    .B1(net2200));
 sg13g2_a21o_1 _6392_ (.A2(_1975_),
    .A1(net2395),
    .B1(_1988_),
    .X(_1989_));
 sg13g2_a221oi_1 _6393_ (.B2(_1989_),
    .C1(net2039),
    .B1(_1986_),
    .A1(net2384),
    .Y(_1990_),
    .A2(_1967_));
 sg13g2_nand4_1 _6394_ (.B(net2262),
    .C(_3144_),
    .A(net2162),
    .Y(_1991_),
    .D(net2208));
 sg13g2_a21oi_1 _6395_ (.A1(net2176),
    .A2(net2065),
    .Y(_1992_),
    .B1(net2404));
 sg13g2_a22oi_1 _6396_ (.Y(_1993_),
    .B1(_1991_),
    .B2(_1992_),
    .A2(_1087_),
    .A1(net2449));
 sg13g2_o21ai_1 _6397_ (.B1(_1993_),
    .Y(_1994_),
    .A1(net2419),
    .A2(_1084_));
 sg13g2_nor2_1 _6398_ (.A(net2500),
    .B(_1821_),
    .Y(_1995_));
 sg13g2_a21oi_1 _6399_ (.A1(net2532),
    .A2(_1485_),
    .Y(_1996_),
    .B1(_1091_));
 sg13g2_and4_1 _6400_ (.A(net2017),
    .B(net2003),
    .C(net1995),
    .D(_1049_),
    .X(_1997_));
 sg13g2_a221oi_1 _6401_ (.B2(_3410_),
    .C1(_1996_),
    .B1(_1997_),
    .A1(_1994_),
    .Y(_1999_),
    .A2(_1995_));
 sg13g2_nand2_1 _6402_ (.Y(_2000_),
    .A(net2481),
    .B(_2901_));
 sg13g2_o21ai_1 _6403_ (.B1(net2205),
    .Y(_2001_),
    .A1(net2177),
    .A2(_2000_));
 sg13g2_nor2_1 _6404_ (.A(_1870_),
    .B(_2001_),
    .Y(_2002_));
 sg13g2_nor2_1 _6405_ (.A(net2192),
    .B(_1821_),
    .Y(_2003_));
 sg13g2_a21oi_1 _6406_ (.A1(_1087_),
    .A2(_2003_),
    .Y(_2004_),
    .B1(_2002_));
 sg13g2_o21ai_1 _6407_ (.B1(_2004_),
    .Y(_2005_),
    .A1(net2397),
    .A2(_1999_));
 sg13g2_o21ai_1 _6408_ (.B1(_0775_),
    .Y(_2006_),
    .A1(net2233),
    .A2(_3255_));
 sg13g2_o21ai_1 _6409_ (.B1(_1090_),
    .Y(_2007_),
    .A1(net2467),
    .A2(_0288_));
 sg13g2_o21ai_1 _6410_ (.B1(net2518),
    .Y(_2008_),
    .A1(_1485_),
    .A2(_2007_));
 sg13g2_o21ai_1 _6411_ (.B1(_1867_),
    .Y(_2010_),
    .A1(_2306_),
    .A2(_3247_));
 sg13g2_a21oi_1 _6412_ (.A1(net2307),
    .A2(_2010_),
    .Y(_2011_),
    .B1(_1873_));
 sg13g2_nand3_1 _6413_ (.B(_2008_),
    .C(_2011_),
    .A(net2397),
    .Y(_2012_));
 sg13g2_nor2b_1 _6414_ (.A(_1058_),
    .B_N(_1867_),
    .Y(_2013_));
 sg13g2_a221oi_1 _6415_ (.B2(net2474),
    .C1(net2393),
    .B1(_1984_),
    .A1(net2497),
    .Y(_2014_),
    .A2(_0165_));
 sg13g2_o21ai_1 _6416_ (.B1(_2014_),
    .Y(_2015_),
    .A1(net2480),
    .A2(_2013_));
 sg13g2_a221oi_1 _6417_ (.B2(_2015_),
    .C1(net1981),
    .B1(_2012_),
    .A1(_3451_),
    .Y(_2016_),
    .A2(_2006_));
 sg13g2_a21oi_1 _6418_ (.A1(net1982),
    .A2(_2005_),
    .Y(_2017_),
    .B1(_2016_));
 sg13g2_nand3b_1 _6419_ (.B(_2017_),
    .C(net1978),
    .Y(_2018_),
    .A_N(_1990_));
 sg13g2_nand4_1 _6420_ (.B(net2046),
    .C(_2750_),
    .A(net2580),
    .Y(_2019_),
    .D(net2025));
 sg13g2_nand4_1 _6421_ (.B(net2046),
    .C(net2044),
    .A(net2559),
    .Y(_2021_),
    .D(_1406_));
 sg13g2_nand3_1 _6422_ (.B(_2019_),
    .C(_2021_),
    .A(net2538),
    .Y(_2022_));
 sg13g2_nor2_1 _6423_ (.A(net2483),
    .B(_1116_),
    .Y(_2023_));
 sg13g2_o21ai_1 _6424_ (.B1(_2863_),
    .Y(_2024_),
    .A1(net2090),
    .A2(_1838_));
 sg13g2_a221oi_1 _6425_ (.B2(net2407),
    .C1(net2502),
    .B1(_2024_),
    .A1(net2470),
    .Y(_2025_),
    .A2(_1176_));
 sg13g2_a22oi_1 _6426_ (.Y(_2026_),
    .B1(_2025_),
    .B2(_1124_),
    .A2(_2023_),
    .A1(_2022_));
 sg13g2_nand3_1 _6427_ (.B(_1423_),
    .C(_1537_),
    .A(net2011),
    .Y(_2027_));
 sg13g2_and2_1 _6428_ (.A(net2305),
    .B(_2027_),
    .X(_2028_));
 sg13g2_a21oi_1 _6429_ (.A1(_3176_),
    .A2(_0398_),
    .Y(_2029_),
    .B1(_1143_));
 sg13g2_nand2_1 _6430_ (.Y(_2030_),
    .A(net2095),
    .B(_0277_));
 sg13g2_a21oi_1 _6431_ (.A1(_1539_),
    .A2(_2030_),
    .Y(_2032_),
    .B1(_0266_));
 sg13g2_a21oi_1 _6432_ (.A1(_0395_),
    .A2(_1523_),
    .Y(_2033_),
    .B1(net2314));
 sg13g2_nand3_1 _6433_ (.B(_3011_),
    .C(net2064),
    .A(net2166),
    .Y(_2034_));
 sg13g2_nand2_1 _6434_ (.Y(_2035_),
    .A(net2026),
    .B(_2034_));
 sg13g2_o21ai_1 _6435_ (.B1(net2309),
    .Y(_2036_),
    .A1(_0626_),
    .A2(_2035_));
 sg13g2_nor2_1 _6436_ (.A(net2562),
    .B(_3158_),
    .Y(_2037_));
 sg13g2_a221oi_1 _6437_ (.B2(_1532_),
    .C1(net2336),
    .B1(_2037_),
    .A1(_1132_),
    .Y(_2038_),
    .A2(_1539_));
 sg13g2_o21ai_1 _6438_ (.B1(_2036_),
    .Y(_2039_),
    .A1(_3454_),
    .A2(_2029_));
 sg13g2_or4_1 _6439_ (.A(_2028_),
    .B(_2032_),
    .C(_2033_),
    .D(_2038_),
    .X(_2040_));
 sg13g2_o21ai_1 _6440_ (.B1(net2390),
    .Y(_2041_),
    .A1(_2039_),
    .A2(_2040_));
 sg13g2_a21oi_1 _6441_ (.A1(net2376),
    .A2(_2026_),
    .Y(_2043_),
    .B1(_3375_));
 sg13g2_and3_1 _6442_ (.X(_2044_),
    .A(_3045_),
    .B(_1374_),
    .C(_1576_));
 sg13g2_nor4_1 _6443_ (.A(_1196_),
    .B(_1571_),
    .C(_1574_),
    .D(_1575_),
    .Y(_2045_));
 sg13g2_o21ai_1 _6444_ (.B1(_2045_),
    .Y(_2046_),
    .A1(net2336),
    .A2(_2044_));
 sg13g2_nor3_1 _6445_ (.A(net2579),
    .B(_3107_),
    .C(_1585_),
    .Y(_2047_));
 sg13g2_a21oi_1 _6446_ (.A1(_3086_),
    .A2(_0585_),
    .Y(_2048_),
    .B1(net2416));
 sg13g2_nor3_1 _6447_ (.A(net2461),
    .B(_3030_),
    .C(_3097_),
    .Y(_2049_));
 sg13g2_nor4_1 _6448_ (.A(net2483),
    .B(_2047_),
    .C(_2048_),
    .D(_2049_),
    .Y(_2050_));
 sg13g2_o21ai_1 _6449_ (.B1(_3061_),
    .Y(_2051_),
    .A1(_3030_),
    .A2(_3093_));
 sg13g2_o21ai_1 _6450_ (.B1(net2312),
    .Y(_2052_),
    .A1(_3026_),
    .A2(_3093_));
 sg13g2_nand2_1 _6451_ (.Y(_2054_),
    .A(net2483),
    .B(_1180_));
 sg13g2_nand4_1 _6452_ (.B(_2051_),
    .C(_2052_),
    .A(net2389),
    .Y(_2055_),
    .D(_2054_));
 sg13g2_o21ai_1 _6453_ (.B1(_2046_),
    .Y(_2056_),
    .A1(_2050_),
    .A2(_2055_));
 sg13g2_a21oi_1 _6454_ (.A1(net2527),
    .A2(_1153_),
    .Y(_2057_),
    .B1(net2488));
 sg13g2_o21ai_1 _6455_ (.B1(_2057_),
    .Y(_2058_),
    .A1(_0694_),
    .A2(_1914_));
 sg13g2_o21ai_1 _6456_ (.B1(net2309),
    .Y(_2059_),
    .A1(net2020),
    .A2(_0434_));
 sg13g2_a22oi_1 _6457_ (.Y(_2060_),
    .B1(_1563_),
    .B2(net2338),
    .A2(_0684_),
    .A1(net2306));
 sg13g2_and4_1 _6458_ (.A(_0682_),
    .B(_1166_),
    .C(_2059_),
    .D(_2060_),
    .X(_2061_));
 sg13g2_a22oi_1 _6459_ (.Y(_2062_),
    .B1(_2061_),
    .B2(_1165_),
    .A2(_2058_),
    .A1(_1160_));
 sg13g2_nor2_1 _6460_ (.A(_3264_),
    .B(net1983),
    .Y(_2063_));
 sg13g2_a21oi_1 _6461_ (.A1(_3296_),
    .A2(_2063_),
    .Y(_2065_),
    .B1(net1979));
 sg13g2_o21ai_1 _6462_ (.B1(_2065_),
    .Y(_2066_),
    .A1(net1985),
    .A2(_2062_));
 sg13g2_a221oi_1 _6463_ (.B2(_3431_),
    .C1(_2066_),
    .B1(_2056_),
    .A1(_2041_),
    .Y(_2067_),
    .A2(_2043_));
 sg13g2_nor2_1 _6464_ (.A(_3308_),
    .B(_2067_),
    .Y(_2068_));
 sg13g2_a221oi_1 _6465_ (.B2(_2068_),
    .C1(_3506_),
    .B1(_2018_),
    .A1(_1937_),
    .Y(_2069_),
    .A2(_1938_));
 sg13g2_a21oi_1 _6466_ (.A1(_1783_),
    .A2(_1784_),
    .Y(_2070_),
    .B1(_2069_));
 sg13g2_nand3b_1 _6467_ (.B(net2016),
    .C(net2600),
    .Y(_2071_),
    .A_N(_3335_));
 sg13g2_o21ai_1 _6468_ (.B1(_2071_),
    .Y(_2072_),
    .A1(net2600),
    .A2(_1203_));
 sg13g2_a21oi_1 _6469_ (.A1(_1053_),
    .A2(_2072_),
    .Y(_2073_),
    .B1(net2327));
 sg13g2_nand3_1 _6470_ (.B(_1053_),
    .C(_1599_),
    .A(net1996),
    .Y(_2074_));
 sg13g2_o21ai_1 _6471_ (.B1(net2321),
    .Y(_2076_),
    .A1(_1597_),
    .A2(_2074_));
 sg13g2_nand3_1 _6472_ (.B(_2614_),
    .C(_0311_),
    .A(net2182),
    .Y(_2077_));
 sg13g2_nand4_1 _6473_ (.B(_0807_),
    .C(_1633_),
    .A(net2557),
    .Y(_2078_),
    .D(_2077_));
 sg13g2_nand3_1 _6474_ (.B(_1053_),
    .C(_1202_),
    .A(net2536),
    .Y(_2079_));
 sg13g2_a21oi_1 _6475_ (.A1(net2414),
    .A2(net2058),
    .Y(_2080_),
    .B1(net2498));
 sg13g2_nand3_1 _6476_ (.B(_2079_),
    .C(_2080_),
    .A(_2078_),
    .Y(_2081_));
 sg13g2_nand3_1 _6477_ (.B(_2076_),
    .C(_2081_),
    .A(_3300_),
    .Y(_2082_));
 sg13g2_nand3_1 _6478_ (.B(_3393_),
    .C(net1986),
    .A(_3183_),
    .Y(_2083_));
 sg13g2_nand3_1 _6479_ (.B(net1986),
    .C(_1594_),
    .A(net2321),
    .Y(_2084_));
 sg13g2_o21ai_1 _6480_ (.B1(_2084_),
    .Y(_2085_),
    .A1(net2321),
    .A2(_2083_));
 sg13g2_a21oi_1 _6481_ (.A1(net1984),
    .A2(_2085_),
    .Y(_2087_),
    .B1(_0559_));
 sg13g2_o21ai_1 _6482_ (.B1(_2087_),
    .Y(_2088_),
    .A1(_2073_),
    .A2(_2082_));
 sg13g2_o21ai_1 _6483_ (.B1(net2448),
    .Y(_2089_),
    .A1(_0824_),
    .A2(_0838_));
 sg13g2_nand4_1 _6484_ (.B(net2030),
    .C(net1988),
    .A(net2598),
    .Y(_2090_),
    .D(_1594_));
 sg13g2_nand3_1 _6485_ (.B(_1605_),
    .C(_2090_),
    .A(net2555),
    .Y(_2091_));
 sg13g2_a21oi_1 _6486_ (.A1(net2481),
    .A2(_2083_),
    .Y(_2092_),
    .B1(net2516));
 sg13g2_a22oi_1 _6487_ (.Y(_2093_),
    .B1(_2091_),
    .B2(_2092_),
    .A2(_2089_),
    .A1(_1601_));
 sg13g2_o21ai_1 _6488_ (.B1(net2536),
    .Y(_2094_),
    .A1(_0546_),
    .A2(_1643_));
 sg13g2_a221oi_1 _6489_ (.B2(net2554),
    .C1(net2516),
    .B1(_1627_),
    .A1(net2415),
    .Y(_2095_),
    .A2(_0751_));
 sg13g2_nand2b_1 _6490_ (.Y(_2096_),
    .B(_1617_),
    .A_N(_0902_));
 sg13g2_nand3_1 _6491_ (.B(_0494_),
    .C(_1287_),
    .A(net2016),
    .Y(_2098_));
 sg13g2_a22oi_1 _6492_ (.Y(_2099_),
    .B1(_2098_),
    .B2(net2448),
    .A2(_2096_),
    .A1(net2427));
 sg13g2_a22oi_1 _6493_ (.Y(_2100_),
    .B1(_2099_),
    .B2(_1619_),
    .A2(_2095_),
    .A1(_2094_));
 sg13g2_nor2_1 _6494_ (.A(net2297),
    .B(_2100_),
    .Y(_2101_));
 sg13g2_o21ai_1 _6495_ (.B1(net2399),
    .Y(_2102_),
    .A1(_1596_),
    .A2(_2093_));
 sg13g2_or2_1 _6496_ (.X(_2103_),
    .B(_2102_),
    .A(_2101_));
 sg13g2_o21ai_1 _6497_ (.B1(net2580),
    .Y(_2104_),
    .A1(_3034_),
    .A2(net2210));
 sg13g2_nand2_1 _6498_ (.Y(_2105_),
    .A(net2236),
    .B(net2216));
 sg13g2_nor4_1 _6499_ (.A(net2579),
    .B(net2138),
    .C(_3145_),
    .D(_2105_),
    .Y(_2106_));
 sg13g2_nor4_1 _6500_ (.A(net2579),
    .B(net2092),
    .C(net2244),
    .D(_2912_),
    .Y(_2107_));
 sg13g2_nor3_1 _6501_ (.A(net2525),
    .B(_2106_),
    .C(_2107_),
    .Y(_2109_));
 sg13g2_o21ai_1 _6502_ (.B1(_2109_),
    .Y(_2110_),
    .A1(_0464_),
    .A2(_2104_));
 sg13g2_nand2_1 _6503_ (.Y(_2111_),
    .A(_1702_),
    .B(_2110_));
 sg13g2_a21oi_1 _6504_ (.A1(_3103_),
    .A2(_3398_),
    .Y(_2112_),
    .B1(net2097));
 sg13g2_o21ai_1 _6505_ (.B1(net2409),
    .Y(_2113_),
    .A1(_1695_),
    .A2(_2112_));
 sg13g2_a21oi_1 _6506_ (.A1(net2423),
    .A2(_2328_),
    .Y(_2114_),
    .B1(net2505));
 sg13g2_nor3_1 _6507_ (.A(net2229),
    .B(_3091_),
    .C(_1430_),
    .Y(_2115_));
 sg13g2_o21ai_1 _6508_ (.B1(net2541),
    .Y(_2116_),
    .A1(_1692_),
    .A2(_2115_));
 sg13g2_nor2_2 _6509_ (.A(net2229),
    .B(_3629_),
    .Y(_2117_));
 sg13g2_o21ai_1 _6510_ (.B1(net2472),
    .Y(_2118_),
    .A1(_0450_),
    .A2(_2117_));
 sg13g2_nand4_1 _6511_ (.B(_2114_),
    .C(_2116_),
    .A(_2113_),
    .Y(_2120_),
    .D(_2118_));
 sg13g2_a21o_1 _6512_ (.A2(_2120_),
    .A1(_2111_),
    .B1(net2390),
    .X(_2121_));
 sg13g2_nand4_1 _6513_ (.B(net2049),
    .C(_0909_),
    .A(net2541),
    .Y(_2122_),
    .D(net1991));
 sg13g2_a22oi_1 _6514_ (.Y(_2123_),
    .B1(_2122_),
    .B2(net2420),
    .A2(_1670_),
    .A1(net2584));
 sg13g2_a21oi_1 _6515_ (.A1(net2562),
    .A2(_1670_),
    .Y(_2124_),
    .B1(net2541));
 sg13g2_nor3_1 _6516_ (.A(net2504),
    .B(_2123_),
    .C(_2124_),
    .Y(_2125_));
 sg13g2_a221oi_1 _6517_ (.B2(_1674_),
    .C1(net2523),
    .B1(_3028_),
    .A1(net2146),
    .Y(_2126_),
    .A2(_3023_));
 sg13g2_a22oi_1 _6518_ (.Y(_2127_),
    .B1(_3253_),
    .B2(net2047),
    .A2(_2778_),
    .A1(net2562));
 sg13g2_a21oi_1 _6519_ (.A1(net2145),
    .A2(_3513_),
    .Y(_2128_),
    .B1(net2541));
 sg13g2_o21ai_1 _6520_ (.B1(_2128_),
    .Y(_2129_),
    .A1(net2235),
    .A2(_3183_));
 sg13g2_o21ai_1 _6521_ (.B1(net2504),
    .Y(_2131_),
    .A1(_2127_),
    .A2(_2129_));
 sg13g2_nand3_1 _6522_ (.B(_0887_),
    .C(_1039_),
    .A(net2047),
    .Y(_2132_));
 sg13g2_a21oi_1 _6523_ (.A1(net2312),
    .A2(_2132_),
    .Y(_2133_),
    .B1(net2377));
 sg13g2_o21ai_1 _6524_ (.B1(_2133_),
    .Y(_2134_),
    .A1(_2126_),
    .A2(_2131_));
 sg13g2_o21ai_1 _6525_ (.B1(_2121_),
    .Y(_2135_),
    .A1(_2125_),
    .A2(_2134_));
 sg13g2_nor2_1 _6526_ (.A(net2571),
    .B(_1287_),
    .Y(_2136_));
 sg13g2_a21oi_1 _6527_ (.A1(_3124_),
    .A2(_1144_),
    .Y(_2137_),
    .B1(net2113));
 sg13g2_o21ai_1 _6528_ (.B1(net2310),
    .Y(_2138_),
    .A1(_0740_),
    .A2(_2137_));
 sg13g2_o21ai_1 _6529_ (.B1(net2168),
    .Y(_2139_),
    .A1(net2085),
    .A2(net2054));
 sg13g2_o21ai_1 _6530_ (.B1(_1227_),
    .Y(_2140_),
    .A1(net2595),
    .A2(_2139_));
 sg13g2_o21ai_1 _6531_ (.B1(net2323),
    .Y(_2142_),
    .A1(_2136_),
    .A2(_2140_));
 sg13g2_nand4_1 _6532_ (.B(net2018),
    .C(_0242_),
    .A(_3132_),
    .Y(_2143_),
    .D(_2139_));
 sg13g2_nand2_1 _6533_ (.Y(_2144_),
    .A(_3453_),
    .B(_2143_));
 sg13g2_o21ai_1 _6534_ (.B1(_3125_),
    .Y(_2145_),
    .A1(_2383_),
    .A2(_3163_));
 sg13g2_a21oi_1 _6535_ (.A1(net2112),
    .A2(_3078_),
    .Y(_2146_),
    .B1(net2466));
 sg13g2_nor2_1 _6536_ (.A(net2476),
    .B(_1421_),
    .Y(_2147_));
 sg13g2_a221oi_1 _6537_ (.B2(_2146_),
    .C1(_2147_),
    .B1(_2145_),
    .A1(_3358_),
    .Y(_2148_),
    .A2(_1136_));
 sg13g2_nand3_1 _6538_ (.B(_2142_),
    .C(_2144_),
    .A(_2138_),
    .Y(_2149_));
 sg13g2_o21ai_1 _6539_ (.B1(net2342),
    .Y(_2150_),
    .A1(_3131_),
    .A2(_1204_));
 sg13g2_a21oi_1 _6540_ (.A1(_2148_),
    .A2(_2150_),
    .Y(_2151_),
    .B1(net2493));
 sg13g2_o21ai_1 _6541_ (.B1(net2382),
    .Y(_2153_),
    .A1(_2149_),
    .A2(_2151_));
 sg13g2_o21ai_1 _6542_ (.B1(net2197),
    .Y(_2154_),
    .A1(_3092_),
    .A2(_0618_));
 sg13g2_nor2_1 _6543_ (.A(_3607_),
    .B(_2154_),
    .Y(_2155_));
 sg13g2_nor2_1 _6544_ (.A(_3432_),
    .B(_2155_),
    .Y(_2156_));
 sg13g2_o21ai_1 _6545_ (.B1(net2410),
    .Y(_2157_),
    .A1(_2438_),
    .A2(net2009));
 sg13g2_o21ai_1 _6546_ (.B1(net1997),
    .Y(_2158_),
    .A1(net2248),
    .A2(_2724_));
 sg13g2_a22oi_1 _6547_ (.Y(_2159_),
    .B1(_2158_),
    .B2(net2425),
    .A2(_1024_),
    .A1(_0398_));
 sg13g2_o21ai_1 _6548_ (.B1(net2443),
    .Y(_2160_),
    .A1(_0450_),
    .A2(_2117_));
 sg13g2_nand4_1 _6549_ (.B(_2157_),
    .C(_2159_),
    .A(_1652_),
    .Y(_2161_),
    .D(_2160_));
 sg13g2_o21ai_1 _6550_ (.B1(net2548),
    .Y(_2162_),
    .A1(_3392_),
    .A2(net2009));
 sg13g2_o21ai_1 _6551_ (.B1(net2411),
    .Y(_2164_),
    .A1(_3392_),
    .A2(_3574_));
 sg13g2_nand2_1 _6552_ (.Y(_2165_),
    .A(net2444),
    .B(_1533_));
 sg13g2_nand4_1 _6553_ (.B(_2162_),
    .C(_2164_),
    .A(_1665_),
    .Y(_2166_),
    .D(_2165_));
 sg13g2_nand3_1 _6554_ (.B(_2161_),
    .C(_2166_),
    .A(net2395),
    .Y(_2167_));
 sg13g2_and3_1 _6555_ (.X(_2168_),
    .A(_2153_),
    .B(_2156_),
    .C(_2167_));
 sg13g2_a221oi_1 _6556_ (.B2(net1982),
    .C1(_2168_),
    .B1(_2135_),
    .A1(_2088_),
    .Y(_2169_),
    .A2(_2103_));
 sg13g2_nand2_2 _6557_ (.Y(_2170_),
    .A(_0429_),
    .B(_0596_));
 sg13g2_o21ai_1 _6558_ (.B1(net2546),
    .Y(_2171_),
    .A1(_1380_),
    .A2(_2170_));
 sg13g2_nor2_1 _6559_ (.A(net2490),
    .B(_1754_),
    .Y(_2172_));
 sg13g2_nor3_1 _6560_ (.A(net2317),
    .B(_3256_),
    .C(_0229_),
    .Y(_2173_));
 sg13g2_o21ai_1 _6561_ (.B1(net2380),
    .Y(_2175_),
    .A1(net2326),
    .A2(_1154_));
 sg13g2_a221oi_1 _6562_ (.B2(_1384_),
    .C1(_2175_),
    .B1(_2173_),
    .A1(_2171_),
    .Y(_2176_),
    .A2(_2172_));
 sg13g2_nand2b_1 _6563_ (.Y(_2177_),
    .B(_1751_),
    .A_N(_2176_));
 sg13g2_nand3_1 _6564_ (.B(_1855_),
    .C(_0656_),
    .A(net2528),
    .Y(_2178_));
 sg13g2_nand3_1 _6565_ (.B(net2236),
    .C(net2217),
    .A(net2474),
    .Y(_2179_));
 sg13g2_a22oi_1 _6566_ (.Y(_2180_),
    .B1(_0451_),
    .B2(net2442),
    .A2(net2212),
    .A1(net2344));
 sg13g2_a21o_1 _6567_ (.A2(_2180_),
    .A1(_2179_),
    .B1(net2104),
    .X(_2181_));
 sg13g2_nand2b_1 _6568_ (.Y(_2182_),
    .B(net2106),
    .A_N(_0288_));
 sg13g2_nand2_1 _6569_ (.Y(_2183_),
    .A(_0808_),
    .B(_2182_));
 sg13g2_o21ai_1 _6570_ (.B1(net2524),
    .Y(_2184_),
    .A1(_3365_),
    .A2(_1739_));
 sg13g2_a21oi_1 _6571_ (.A1(net2083),
    .A2(_3528_),
    .Y(_2186_),
    .B1(net2238));
 sg13g2_a21oi_1 _6572_ (.A1(net2145),
    .A2(_2186_),
    .Y(_2187_),
    .B1(_3365_));
 sg13g2_a221oi_1 _6573_ (.B2(_3354_),
    .C1(net2429),
    .B1(_0257_),
    .A1(_3125_),
    .Y(_2188_),
    .A2(_0155_));
 sg13g2_o21ai_1 _6574_ (.B1(_2184_),
    .Y(_2189_),
    .A1(net2417),
    .A2(_2187_));
 sg13g2_or2_1 _6575_ (.X(_2190_),
    .B(_2188_),
    .A(_3606_));
 sg13g2_o21ai_1 _6576_ (.B1(net2202),
    .Y(_2191_),
    .A1(_2189_),
    .A2(_2190_));
 sg13g2_mux2_1 _6577_ (.A0(_3154_),
    .A1(_0169_),
    .S(net2106),
    .X(_2192_));
 sg13g2_o21ai_1 _6578_ (.B1(net2589),
    .Y(_2193_),
    .A1(_3514_),
    .A2(_2192_));
 sg13g2_nor4_1 _6579_ (.A(net2528),
    .B(_3514_),
    .C(_3594_),
    .D(_0434_),
    .Y(_2194_));
 sg13g2_a221oi_1 _6580_ (.B2(_2194_),
    .C1(net2194),
    .B1(_2193_),
    .A1(_1742_),
    .Y(_2195_),
    .A2(_2183_));
 sg13g2_nor2_1 _6581_ (.A(net1981),
    .B(_2195_),
    .Y(_2197_));
 sg13g2_a21oi_1 _6582_ (.A1(net2152),
    .A2(_0157_),
    .Y(_2198_),
    .B1(net2403));
 sg13g2_o21ai_1 _6583_ (.B1(net2474),
    .Y(_2199_),
    .A1(_3514_),
    .A2(_2192_));
 sg13g2_a21oi_1 _6584_ (.A1(_0808_),
    .A2(_2198_),
    .Y(_2200_),
    .B1(net2490));
 sg13g2_nand3_1 _6585_ (.B(_0808_),
    .C(_2182_),
    .A(net2545),
    .Y(_2201_));
 sg13g2_nand3_1 _6586_ (.B(_2200_),
    .C(_2201_),
    .A(_2199_),
    .Y(_2202_));
 sg13g2_a221oi_1 _6587_ (.B2(net2424),
    .C1(net2510),
    .B1(_1730_),
    .A1(net2442),
    .Y(_2203_),
    .A2(_0434_));
 sg13g2_nand4_1 _6588_ (.B(_2178_),
    .C(_2181_),
    .A(_3595_),
    .Y(_2204_),
    .D(_2203_));
 sg13g2_nand3_1 _6589_ (.B(_2202_),
    .C(_2204_),
    .A(net2380),
    .Y(_2205_));
 sg13g2_nand3_1 _6590_ (.B(_2197_),
    .C(_2205_),
    .A(_2191_),
    .Y(_2206_));
 sg13g2_a21oi_1 _6591_ (.A1(_3053_),
    .A2(_1761_),
    .Y(_2208_),
    .B1(net2402));
 sg13g2_o21ai_1 _6592_ (.B1(net2195),
    .Y(_2209_),
    .A1(_1768_),
    .A2(_2208_));
 sg13g2_nand2_1 _6593_ (.Y(_2210_),
    .A(net2475),
    .B(_1821_));
 sg13g2_nor2_1 _6594_ (.A(_3293_),
    .B(_3574_),
    .Y(_2211_));
 sg13g2_or3_1 _6595_ (.A(net2544),
    .B(_3293_),
    .C(_3574_),
    .X(_2212_));
 sg13g2_nand4_1 _6596_ (.B(_1901_),
    .C(_2210_),
    .A(_1771_),
    .Y(_2213_),
    .D(_2212_));
 sg13g2_a21oi_1 _6597_ (.A1(net2024),
    .A2(_0227_),
    .Y(_2214_),
    .B1(net2402));
 sg13g2_nand2_1 _6598_ (.Y(_2215_),
    .A(net2473),
    .B(_1764_));
 sg13g2_nand2_1 _6599_ (.Y(_2216_),
    .A(net2462),
    .B(_3033_));
 sg13g2_nand2_1 _6600_ (.Y(_2217_),
    .A(net2473),
    .B(_0783_));
 sg13g2_nand4_1 _6601_ (.B(_0951_),
    .C(_2216_),
    .A(net2506),
    .Y(_2219_),
    .D(_2217_));
 sg13g2_nand3_1 _6602_ (.B(_2213_),
    .C(_2219_),
    .A(net2379),
    .Y(_2220_));
 sg13g2_a221oi_1 _6603_ (.B2(net2473),
    .C1(_2214_),
    .B1(_1764_),
    .A1(net2547),
    .Y(_2221_),
    .A2(_1333_));
 sg13g2_nand2b_1 _6604_ (.Y(_2222_),
    .B(net2203),
    .A_N(_2221_));
 sg13g2_nand4_1 _6605_ (.B(_2209_),
    .C(_2220_),
    .A(net1984),
    .Y(_2223_),
    .D(_2222_));
 sg13g2_nand3_1 _6606_ (.B(_2206_),
    .C(_2223_),
    .A(_2177_),
    .Y(_2224_));
 sg13g2_a21oi_1 _6607_ (.A1(net1978),
    .A2(_2224_),
    .Y(_2225_),
    .B1(net1976));
 sg13g2_o21ai_1 _6608_ (.B1(_2225_),
    .Y(_2226_),
    .A1(net1978),
    .A2(_2169_));
 sg13g2_o21ai_1 _6609_ (.B1(net2551),
    .Y(_2227_),
    .A1(_0832_),
    .A2(_1402_));
 sg13g2_nand3_1 _6610_ (.B(net2005),
    .C(_0730_),
    .A(_3566_),
    .Y(_2228_));
 sg13g2_nand2_1 _6611_ (.Y(_2230_),
    .A(net2478),
    .B(_2228_));
 sg13g2_a21oi_1 _6612_ (.A1(net2018),
    .A2(net1991),
    .Y(_2231_),
    .B1(net2434));
 sg13g2_nor2_1 _6613_ (.A(net2494),
    .B(_2231_),
    .Y(_2232_));
 sg13g2_a21oi_1 _6614_ (.A1(net2084),
    .A2(_3020_),
    .Y(_2233_),
    .B1(net2124));
 sg13g2_o21ai_1 _6615_ (.B1(net2413),
    .Y(_2234_),
    .A1(_0740_),
    .A2(_2233_));
 sg13g2_nand4_1 _6616_ (.B(_2230_),
    .C(_2232_),
    .A(_2227_),
    .Y(_2235_),
    .D(_2234_));
 sg13g2_nand3_1 _6617_ (.B(_0098_),
    .C(_1421_),
    .A(net2011),
    .Y(_2236_));
 sg13g2_a21oi_1 _6618_ (.A1(net2011),
    .A2(_2034_),
    .Y(_2237_),
    .B1(net2465));
 sg13g2_o21ai_1 _6619_ (.B1(net2070),
    .Y(_2238_),
    .A1(net2229),
    .A2(_2826_));
 sg13g2_a21oi_1 _6620_ (.A1(_3566_),
    .A2(_0744_),
    .Y(_2239_),
    .B1(net2529));
 sg13g2_a22oi_1 _6621_ (.Y(_2241_),
    .B1(_2238_),
    .B2(_3606_),
    .A2(_2236_),
    .A1(net2412));
 sg13g2_nor3_1 _6622_ (.A(net2512),
    .B(_2237_),
    .C(_2239_),
    .Y(_2242_));
 sg13g2_nand2_1 _6623_ (.Y(_2243_),
    .A(_2241_),
    .B(_2242_));
 sg13g2_a21o_2 _6624_ (.A2(_2243_),
    .A1(_2235_),
    .B1(net2396),
    .X(_2244_));
 sg13g2_a21oi_1 _6625_ (.A1(_3546_),
    .A2(_1434_),
    .Y(_2245_),
    .B1(net2438));
 sg13g2_or4_1 _6626_ (.A(_1441_),
    .B(_1442_),
    .C(_1444_),
    .D(_2245_),
    .X(_2246_));
 sg13g2_nand4_1 _6627_ (.B(net2018),
    .C(net1994),
    .A(_3156_),
    .Y(_2247_),
    .D(_1432_));
 sg13g2_o21ai_1 _6628_ (.B1(net2309),
    .Y(_2248_),
    .A1(_0638_),
    .A2(_1439_));
 sg13g2_o21ai_1 _6629_ (.B1(net2307),
    .Y(_2249_),
    .A1(_0732_),
    .A2(_1435_));
 sg13g2_nand3_1 _6630_ (.B(_2248_),
    .C(_2249_),
    .A(net2396),
    .Y(_2250_));
 sg13g2_a221oi_1 _6631_ (.B2(net2323),
    .C1(_2250_),
    .B1(_2247_),
    .A1(net2512),
    .Y(_2252_),
    .A2(_2246_));
 sg13g2_nor2_1 _6632_ (.A(net2039),
    .B(_2252_),
    .Y(_2253_));
 sg13g2_a21o_1 _6633_ (.A2(_1472_),
    .A1(net2598),
    .B1(_1494_),
    .X(_2254_));
 sg13g2_nand3_1 _6634_ (.B(net1989),
    .C(_1471_),
    .A(_0094_),
    .Y(_2255_));
 sg13g2_a221oi_1 _6635_ (.B2(_0561_),
    .C1(net2399),
    .B1(_2255_),
    .A1(net2309),
    .Y(_2256_),
    .A2(_1472_));
 sg13g2_nand3_1 _6636_ (.B(net1990),
    .C(net1986),
    .A(net2576),
    .Y(_2257_));
 sg13g2_and2_1 _6637_ (.A(net2335),
    .B(_2257_),
    .X(_2258_));
 sg13g2_a22oi_1 _6638_ (.Y(_2259_),
    .B1(_2258_),
    .B2(_1606_),
    .A2(_2254_),
    .A1(net2340));
 sg13g2_a21o_1 _6639_ (.A2(net1986),
    .A1(net1989),
    .B1(net2315),
    .X(_2260_));
 sg13g2_a221oi_1 _6640_ (.B2(_1488_),
    .C1(net2036),
    .B1(_2260_),
    .A1(_2256_),
    .Y(_2261_),
    .A2(_2259_));
 sg13g2_a21o_1 _6641_ (.A2(_2253_),
    .A1(_2244_),
    .B1(_2261_),
    .X(_2263_));
 sg13g2_nand2_1 _6642_ (.Y(_2264_),
    .A(net2598),
    .B(net1986));
 sg13g2_nand3_1 _6643_ (.B(_3322_),
    .C(net1988),
    .A(net2576),
    .Y(_2265_));
 sg13g2_a22oi_1 _6644_ (.Y(_2266_),
    .B1(_2264_),
    .B2(_2265_),
    .A2(_1473_),
    .A1(_0298_));
 sg13g2_nor2_1 _6645_ (.A(net2555),
    .B(_2266_),
    .Y(_2267_));
 sg13g2_a21oi_1 _6646_ (.A1(net2598),
    .A2(_1472_),
    .Y(_2268_),
    .B1(_2255_));
 sg13g2_nor2_1 _6647_ (.A(net2535),
    .B(_2268_),
    .Y(_2269_));
 sg13g2_o21ai_1 _6648_ (.B1(net2205),
    .Y(_2270_),
    .A1(_2267_),
    .A2(_2269_));
 sg13g2_a21oi_1 _6649_ (.A1(net2015),
    .A2(net2004),
    .Y(_2271_),
    .B1(net2599));
 sg13g2_nor2_1 _6650_ (.A(_1455_),
    .B(_2271_),
    .Y(_2272_));
 sg13g2_a21oi_1 _6651_ (.A1(_1458_),
    .A2(_2272_),
    .Y(_2274_),
    .B1(net2192));
 sg13g2_nand2b_1 _6652_ (.Y(_2275_),
    .B(_2274_),
    .A_N(_1454_));
 sg13g2_a21oi_1 _6653_ (.A1(net2599),
    .A2(_0301_),
    .Y(_2276_),
    .B1(_2271_));
 sg13g2_a21oi_1 _6654_ (.A1(_1053_),
    .A2(_2276_),
    .Y(_2277_),
    .B1(net2327));
 sg13g2_nand3_1 _6655_ (.B(net2015),
    .C(net1993),
    .A(_3349_),
    .Y(_2278_));
 sg13g2_a221oi_1 _6656_ (.B2(net2414),
    .C1(_0296_),
    .B1(_0774_),
    .A1(_3026_),
    .Y(_2279_),
    .A2(net2052));
 sg13g2_a22oi_1 _6657_ (.Y(_2280_),
    .B1(_2278_),
    .B2(net2311),
    .A2(_1463_),
    .A1(net2321));
 sg13g2_o21ai_1 _6658_ (.B1(_2280_),
    .Y(_2281_),
    .A1(net2498),
    .A2(_2279_));
 sg13g2_o21ai_1 _6659_ (.B1(net2384),
    .Y(_2282_),
    .A1(_2277_),
    .A2(_2281_));
 sg13g2_nand3_1 _6660_ (.B(_2275_),
    .C(_2282_),
    .A(_2270_),
    .Y(_2283_));
 sg13g2_nand3_1 _6661_ (.B(net1986),
    .C(_1594_),
    .A(net2576),
    .Y(_2285_));
 sg13g2_nand3_1 _6662_ (.B(net1989),
    .C(net1986),
    .A(net2598),
    .Y(_2286_));
 sg13g2_a21oi_1 _6663_ (.A1(_2285_),
    .A2(_2286_),
    .Y(_2287_),
    .B1(net2331));
 sg13g2_nor3_1 _6664_ (.A(net2517),
    .B(_1478_),
    .C(_1501_),
    .Y(_2288_));
 sg13g2_nand4_1 _6665_ (.B(_3183_),
    .C(_3388_),
    .A(net2598),
    .Y(_2289_),
    .D(net1986));
 sg13g2_a21oi_1 _6666_ (.A1(_2257_),
    .A2(_2289_),
    .Y(_2290_),
    .B1(net2337));
 sg13g2_nor4_1 _6667_ (.A(net2384),
    .B(_2287_),
    .C(_2288_),
    .D(_2290_),
    .Y(_2291_));
 sg13g2_o21ai_1 _6668_ (.B1(net1982),
    .Y(_2292_),
    .A1(_1510_),
    .A2(_2291_));
 sg13g2_nand2_1 _6669_ (.Y(_2293_),
    .A(net1980),
    .B(_2292_));
 sg13g2_a221oi_1 _6670_ (.B2(_3300_),
    .C1(_2293_),
    .B1(_2283_),
    .A1(net2296),
    .Y(_2294_),
    .A2(_2263_));
 sg13g2_nand4_1 _6671_ (.B(net2042),
    .C(_3075_),
    .A(net2521),
    .Y(_2296_),
    .D(_0720_));
 sg13g2_a21oi_1 _6672_ (.A1(net2461),
    .A2(_2296_),
    .Y(_2297_),
    .B1(_1543_));
 sg13g2_nor3_1 _6673_ (.A(net2429),
    .B(_2328_),
    .C(_3191_),
    .Y(_2298_));
 sg13g2_nor3_1 _6674_ (.A(net2416),
    .B(net2034),
    .C(_3191_),
    .Y(_2299_));
 sg13g2_nor4_2 _6675_ (.A(net2502),
    .B(_2297_),
    .C(_2298_),
    .Y(_2300_),
    .D(_2299_));
 sg13g2_nand3_1 _6676_ (.B(_3192_),
    .C(_1258_),
    .A(_2339_),
    .Y(_2301_));
 sg13g2_o21ai_1 _6677_ (.B1(_3586_),
    .Y(_2302_),
    .A1(_3576_),
    .A2(net2002));
 sg13g2_nor2_1 _6678_ (.A(_2328_),
    .B(_2302_),
    .Y(_2303_));
 sg13g2_o21ai_1 _6679_ (.B1(_3195_),
    .Y(_2304_),
    .A1(_3605_),
    .A2(_0376_));
 sg13g2_a22oi_1 _6680_ (.Y(_2305_),
    .B1(_2304_),
    .B2(net2305),
    .A2(_2301_),
    .A1(net2339));
 sg13g2_o21ai_1 _6681_ (.B1(_2305_),
    .Y(_2307_),
    .A1(_0266_),
    .A2(_2303_));
 sg13g2_o21ai_1 _6682_ (.B1(net2377),
    .Y(_2308_),
    .A1(_2300_),
    .A2(_2307_));
 sg13g2_nor3_1 _6683_ (.A(net2029),
    .B(_0177_),
    .C(_1527_),
    .Y(_2309_));
 sg13g2_a21oi_1 _6684_ (.A1(net2026),
    .A2(_2309_),
    .Y(_2310_),
    .B1(net2464));
 sg13g2_a21o_1 _6685_ (.A2(_1539_),
    .A1(_1537_),
    .B1(net2430),
    .X(_2311_));
 sg13g2_nor2_1 _6686_ (.A(_1533_),
    .B(_1538_),
    .Y(_2312_));
 sg13g2_o21ai_1 _6687_ (.B1(_2311_),
    .Y(_2313_),
    .A1(net2341),
    .A2(_2312_));
 sg13g2_o21ai_1 _6688_ (.B1(net2202),
    .Y(_2314_),
    .A1(_2310_),
    .A2(_2313_));
 sg13g2_nand2_1 _6689_ (.Y(_2315_),
    .A(_3150_),
    .B(_0789_));
 sg13g2_nand3_1 _6690_ (.B(_0399_),
    .C(_0789_),
    .A(_3150_),
    .Y(_2316_));
 sg13g2_nand2_1 _6691_ (.Y(_2318_),
    .A(net2522),
    .B(_2316_));
 sg13g2_a21oi_2 _6692_ (.B1(_3473_),
    .Y(_2319_),
    .A2(_3131_),
    .A1(net2364));
 sg13g2_a21oi_1 _6693_ (.A1(_3130_),
    .A2(_3155_),
    .Y(_2320_),
    .B1(net2435));
 sg13g2_a21o_1 _6694_ (.A2(_0913_),
    .A1(net2079),
    .B1(net2110),
    .X(_2321_));
 sg13g2_a21oi_1 _6695_ (.A1(_3168_),
    .A2(_2321_),
    .Y(_2322_),
    .B1(net2419));
 sg13g2_a221oi_1 _6696_ (.B2(_2320_),
    .C1(_2322_),
    .B1(_2319_),
    .A1(net2476),
    .Y(_2323_),
    .A2(_0641_));
 sg13g2_a21o_1 _6697_ (.A2(_2323_),
    .A1(_2318_),
    .B1(net2194),
    .X(_2324_));
 sg13g2_nand4_1 _6698_ (.B(_2308_),
    .C(_2314_),
    .A(net1982),
    .Y(_2325_),
    .D(_2324_));
 sg13g2_a221oi_1 _6699_ (.B2(_3255_),
    .C1(net2491),
    .B1(_1559_),
    .A1(net2432),
    .Y(_2326_),
    .A2(_1153_));
 sg13g2_nor4_1 _6700_ (.A(net2392),
    .B(_1556_),
    .C(_1557_),
    .D(_2326_),
    .Y(_2327_));
 sg13g2_or2_1 _6701_ (.X(_2329_),
    .B(_2327_),
    .A(_1165_));
 sg13g2_nor2_1 _6702_ (.A(net2022),
    .B(_0684_),
    .Y(_2330_));
 sg13g2_o21ai_1 _6703_ (.B1(_3289_),
    .Y(_2331_),
    .A1(_3253_),
    .A2(_0166_));
 sg13g2_nor2_1 _6704_ (.A(_2330_),
    .B(_2331_),
    .Y(_2332_));
 sg13g2_nor3_1 _6705_ (.A(net1985),
    .B(_1565_),
    .C(_2332_),
    .Y(_2333_));
 sg13g2_a21oi_1 _6706_ (.A1(_2863_),
    .A2(_3031_),
    .Y(_2334_),
    .B1(net2579));
 sg13g2_o21ai_1 _6707_ (.B1(net2520),
    .Y(_2335_),
    .A1(_1583_),
    .A2(_2334_));
 sg13g2_nand3b_1 _6708_ (.B(_2335_),
    .C(net2202),
    .Y(_2336_),
    .A_N(_1585_));
 sg13g2_nand2b_1 _6709_ (.Y(_2337_),
    .B(_1179_),
    .A_N(_3026_));
 sg13g2_nand2_1 _6710_ (.Y(_2338_),
    .A(net2409),
    .B(_2337_));
 sg13g2_nor3_1 _6711_ (.A(net2461),
    .B(_3293_),
    .C(_3574_),
    .Y(_2340_));
 sg13g2_nor3_1 _6712_ (.A(net2194),
    .B(_1180_),
    .C(_2340_),
    .Y(_2341_));
 sg13g2_a22oi_1 _6713_ (.Y(_2342_),
    .B1(_3618_),
    .B2(net2312),
    .A2(_3238_),
    .A1(net2319));
 sg13g2_nand2_1 _6714_ (.Y(_2343_),
    .A(net2315),
    .B(_3420_));
 sg13g2_a21oi_1 _6715_ (.A1(net2148),
    .A2(net2318),
    .Y(_2344_),
    .B1(_3419_));
 sg13g2_o21ai_1 _6716_ (.B1(_2344_),
    .Y(_2345_),
    .A1(_3056_),
    .A2(_1373_));
 sg13g2_o21ai_1 _6717_ (.B1(_0426_),
    .Y(_2346_),
    .A1(net2045),
    .A2(_1189_));
 sg13g2_o21ai_1 _6718_ (.B1(_3045_),
    .Y(_2347_),
    .A1(net2585),
    .A2(_1820_));
 sg13g2_o21ai_1 _6719_ (.B1(net2334),
    .Y(_2348_),
    .A1(_3084_),
    .A2(_2347_));
 sg13g2_and4_1 _6720_ (.A(net2376),
    .B(_2342_),
    .C(_2345_),
    .D(_2346_),
    .X(_2349_));
 sg13g2_a22oi_1 _6721_ (.Y(_2351_),
    .B1(_2348_),
    .B2(_2349_),
    .A2(_2341_),
    .A1(_2338_));
 sg13g2_a21oi_2 _6722_ (.B1(net1981),
    .Y(_2352_),
    .A2(_2351_),
    .A1(_2336_));
 sg13g2_a221oi_1 _6723_ (.B2(_2333_),
    .C1(_2352_),
    .B1(_2329_),
    .A1(net1984),
    .Y(_2353_),
    .A2(_1520_));
 sg13g2_a21oi_1 _6724_ (.A1(_2325_),
    .A2(_2353_),
    .Y(_2354_),
    .B1(net1979));
 sg13g2_or3_1 _6725_ (.A(_3308_),
    .B(_2294_),
    .C(_2354_),
    .X(_2355_));
 sg13g2_a21o_1 _6726_ (.A2(_2355_),
    .A1(_2226_),
    .B1(_3506_),
    .X(_2356_));
 sg13g2_a21oi_1 _6727_ (.A1(_1202_),
    .A2(_1221_),
    .Y(_2357_),
    .B1(net2418));
 sg13g2_o21ai_1 _6728_ (.B1(_0847_),
    .Y(_2358_),
    .A1(net2600),
    .A2(_0555_));
 sg13g2_nor2_1 _6729_ (.A(net2341),
    .B(_0555_),
    .Y(_2359_));
 sg13g2_nor2_1 _6730_ (.A(_3299_),
    .B(_0738_),
    .Y(_2360_));
 sg13g2_o21ai_1 _6731_ (.B1(net2536),
    .Y(_2362_),
    .A1(_3436_),
    .A2(_2358_));
 sg13g2_nor3_1 _6732_ (.A(net2498),
    .B(_1634_),
    .C(_2357_),
    .Y(_2363_));
 sg13g2_a21o_1 _6733_ (.A2(_0849_),
    .A1(_3435_),
    .B1(net2536),
    .X(_2364_));
 sg13g2_o21ai_1 _6734_ (.B1(net2494),
    .Y(_2365_),
    .A1(net2468),
    .A2(net2001));
 sg13g2_nor3_1 _6735_ (.A(_2359_),
    .B(_2360_),
    .C(_2365_),
    .Y(_2366_));
 sg13g2_a221oi_1 _6736_ (.B2(_2366_),
    .C1(net2399),
    .B1(_2364_),
    .A1(_2362_),
    .Y(_2367_),
    .A2(_2363_));
 sg13g2_nand3_1 _6737_ (.B(net1996),
    .C(_2034_),
    .A(net2030),
    .Y(_2368_));
 sg13g2_a21oi_1 _6738_ (.A1(_0141_),
    .A2(_0529_),
    .Y(_2369_),
    .B1(net2435));
 sg13g2_a221oi_1 _6739_ (.B2(net2426),
    .C1(_2369_),
    .B1(_2368_),
    .A1(net2530),
    .Y(_2370_),
    .A2(_0787_));
 sg13g2_o21ai_1 _6740_ (.B1(net2303),
    .Y(_2371_),
    .A1(net2193),
    .A2(_2370_));
 sg13g2_nand2_2 _6741_ (.Y(_2373_),
    .A(net2575),
    .B(net2356));
 sg13g2_nand3_1 _6742_ (.B(_1612_),
    .C(_2373_),
    .A(_0529_),
    .Y(_2374_));
 sg13g2_o21ai_1 _6743_ (.B1(net2016),
    .Y(_2375_),
    .A1(net2248),
    .A2(_2724_));
 sg13g2_o21ai_1 _6744_ (.B1(net2426),
    .Y(_2376_),
    .A1(_0902_),
    .A2(_2375_));
 sg13g2_a21oi_1 _6745_ (.A1(net2355),
    .A2(_3161_),
    .Y(_2377_),
    .B1(net2265));
 sg13g2_o21ai_1 _6746_ (.B1(_1287_),
    .Y(_2378_),
    .A1(net2001),
    .A2(_2377_));
 sg13g2_a22oi_1 _6747_ (.Y(_2379_),
    .B1(_2378_),
    .B2(net2445),
    .A2(_2374_),
    .A1(net2530));
 sg13g2_a21oi_1 _6748_ (.A1(_2376_),
    .A2(_2379_),
    .Y(_2380_),
    .B1(net2200));
 sg13g2_or3_2 _6749_ (.A(_2367_),
    .B(_2371_),
    .C(_2380_),
    .X(_2381_));
 sg13g2_nor2_1 _6750_ (.A(_0298_),
    .B(_1226_),
    .Y(_2382_));
 sg13g2_o21ai_1 _6751_ (.B1(net2057),
    .Y(_2384_),
    .A1(_3090_),
    .A2(_0428_));
 sg13g2_a22oi_1 _6752_ (.Y(_2385_),
    .B1(_2384_),
    .B2(_1453_),
    .A2(_2382_),
    .A1(net2555));
 sg13g2_o21ai_1 _6753_ (.B1(net2206),
    .Y(_2386_),
    .A1(_1597_),
    .A2(_2385_));
 sg13g2_a21oi_1 _6754_ (.A1(_2647_),
    .A2(net2211),
    .Y(_2387_),
    .B1(net1987));
 sg13g2_a221oi_1 _6755_ (.B2(_2387_),
    .C1(net2398),
    .B1(_3393_),
    .A1(net2497),
    .Y(_2388_),
    .A2(net2437));
 sg13g2_nor3_1 _6756_ (.A(net2177),
    .B(net2212),
    .C(net2060),
    .Y(_2389_));
 sg13g2_nor2_1 _6757_ (.A(net1987),
    .B(_2389_),
    .Y(_2390_));
 sg13g2_a21oi_1 _6758_ (.A1(net2192),
    .A2(_0560_),
    .Y(_2391_),
    .B1(_2390_));
 sg13g2_nor3_1 _6759_ (.A(net2303),
    .B(_2388_),
    .C(_2391_),
    .Y(_2392_));
 sg13g2_a21oi_2 _6760_ (.B1(net2037),
    .Y(_2393_),
    .A2(_2392_),
    .A1(_2386_));
 sg13g2_o21ai_1 _6761_ (.B1(_1227_),
    .Y(_2395_),
    .A1(net2595),
    .A2(net2230));
 sg13g2_o21ai_1 _6762_ (.B1(net2529),
    .Y(_2396_),
    .A1(_0739_),
    .A2(_2395_));
 sg13g2_nor3_1 _6763_ (.A(net2163),
    .B(net2067),
    .C(_0328_),
    .Y(_2397_));
 sg13g2_nor3_1 _6764_ (.A(net2116),
    .B(net2065),
    .C(_1715_),
    .Y(_2398_));
 sg13g2_or3_1 _6765_ (.A(net2419),
    .B(_2397_),
    .C(_2398_),
    .X(_2399_));
 sg13g2_nor3_1 _6766_ (.A(net2164),
    .B(_3076_),
    .C(_1430_),
    .Y(_2400_));
 sg13g2_o21ai_1 _6767_ (.B1(net2443),
    .Y(_2401_),
    .A1(_2137_),
    .A2(_2400_));
 sg13g2_nand4_1 _6768_ (.B(_2396_),
    .C(_2399_),
    .A(net2493),
    .Y(_2402_),
    .D(_2401_));
 sg13g2_nand3_1 _6769_ (.B(net2374),
    .C(_3077_),
    .A(net2593),
    .Y(_2403_));
 sg13g2_nand3_1 _6770_ (.B(_3343_),
    .C(_2403_),
    .A(net2113),
    .Y(_2404_));
 sg13g2_nand3_1 _6771_ (.B(_2816_),
    .C(net2023),
    .A(net2227),
    .Y(_2406_));
 sg13g2_a21oi_1 _6772_ (.A1(_2145_),
    .A2(_2404_),
    .Y(_2407_),
    .B1(net2337));
 sg13g2_nand3b_1 _6773_ (.B(_0308_),
    .C(_0880_),
    .Y(_2408_),
    .A_N(_3570_));
 sg13g2_nand3_1 _6774_ (.B(net2219),
    .C(_3397_),
    .A(net2118),
    .Y(_2409_));
 sg13g2_and3_1 _6775_ (.X(_2410_),
    .A(net2335),
    .B(net2007),
    .C(_2409_));
 sg13g2_a22oi_1 _6776_ (.Y(_2411_),
    .B1(_2408_),
    .B2(_2410_),
    .A2(_2407_),
    .A1(_2406_));
 sg13g2_a21o_1 _6777_ (.A2(_2411_),
    .A1(_2402_),
    .B1(net2395),
    .X(_2412_));
 sg13g2_nor3_1 _6778_ (.A(net2375),
    .B(_3153_),
    .C(_3253_),
    .Y(_2413_));
 sg13g2_nand2_1 _6779_ (.Y(_2414_),
    .A(net2584),
    .B(_0130_));
 sg13g2_nor4_1 _6780_ (.A(net2522),
    .B(_0450_),
    .C(_0473_),
    .D(_2413_),
    .Y(_2415_));
 sg13g2_nor3_1 _6781_ (.A(net2403),
    .B(net2063),
    .C(_0165_),
    .Y(_2417_));
 sg13g2_a22oi_1 _6782_ (.Y(_2418_),
    .B1(_2417_),
    .B2(_0229_),
    .A2(_2415_),
    .A1(_2414_));
 sg13g2_nor4_1 _6783_ (.A(net2570),
    .B(_3594_),
    .C(_1538_),
    .D(_1653_),
    .Y(_2419_));
 sg13g2_nor2_1 _6784_ (.A(_3028_),
    .B(_0398_),
    .Y(_2420_));
 sg13g2_o21ai_1 _6785_ (.B1(net2531),
    .Y(_2421_),
    .A1(_2419_),
    .A2(_2420_));
 sg13g2_a21oi_1 _6786_ (.A1(_2418_),
    .A2(_2421_),
    .Y(_2422_),
    .B1(net2200));
 sg13g2_nand2b_1 _6787_ (.Y(_2423_),
    .B(_2409_),
    .A_N(_0920_));
 sg13g2_nand2_1 _6788_ (.Y(_2424_),
    .A(net2410),
    .B(_2423_));
 sg13g2_a21oi_2 _6789_ (.B1(net2465),
    .Y(_2425_),
    .A2(_2409_),
    .A1(net2007));
 sg13g2_a221oi_1 _6790_ (.B2(net2343),
    .C1(net2193),
    .B1(_3392_),
    .A1(net2476),
    .Y(_2426_),
    .A2(net2028));
 sg13g2_nor2b_1 _6791_ (.A(_2425_),
    .B_N(_2426_),
    .Y(_2428_));
 sg13g2_o21ai_1 _6792_ (.B1(net2443),
    .Y(_2429_),
    .A1(_3541_),
    .A2(_1538_));
 sg13g2_o21ai_1 _6793_ (.B1(net2425),
    .Y(_2430_),
    .A1(_0622_),
    .A2(_1662_));
 sg13g2_and4_1 _6794_ (.A(_2424_),
    .B(_2428_),
    .C(_2429_),
    .D(_2430_),
    .X(_2431_));
 sg13g2_nor3_1 _6795_ (.A(net1981),
    .B(_2422_),
    .C(_2431_),
    .Y(_2432_));
 sg13g2_nand3_1 _6796_ (.B(net2047),
    .C(_2734_),
    .A(net2560),
    .Y(_2433_));
 sg13g2_a21oi_1 _6797_ (.A1(_2104_),
    .A2(_2433_),
    .Y(_2434_),
    .B1(_3074_));
 sg13g2_nor2_1 _6798_ (.A(net2330),
    .B(_2434_),
    .Y(_2435_));
 sg13g2_a22oi_1 _6799_ (.Y(_2436_),
    .B1(_2117_),
    .B2(net2320),
    .A2(_2112_),
    .A1(net2312));
 sg13g2_nand2_1 _6800_ (.Y(_2437_),
    .A(net2051),
    .B(_1694_));
 sg13g2_nand2_1 _6801_ (.Y(_2439_),
    .A(_2328_),
    .B(_3061_));
 sg13g2_a22oi_1 _6802_ (.Y(_2440_),
    .B1(_1115_),
    .B2(net2309),
    .A2(_0890_),
    .A1(_0426_));
 sg13g2_a22oi_1 _6803_ (.Y(_2441_),
    .B1(_2437_),
    .B2(net2306),
    .A2(_1700_),
    .A1(net2338));
 sg13g2_nand4_1 _6804_ (.B(_2439_),
    .C(_2440_),
    .A(_2436_),
    .Y(_2442_),
    .D(_2441_));
 sg13g2_o21ai_1 _6805_ (.B1(net2376),
    .Y(_2443_),
    .A1(_2435_),
    .A2(_2442_));
 sg13g2_a21oi_1 _6806_ (.A1(net2240),
    .A2(_2383_),
    .Y(_2444_),
    .B1(net2140));
 sg13g2_nor3_2 _6807_ (.A(net2353),
    .B(net2034),
    .C(_2444_),
    .Y(_2445_));
 sg13g2_nand3_1 _6808_ (.B(_0978_),
    .C(net1991),
    .A(net2049),
    .Y(_2446_));
 sg13g2_a22oi_1 _6809_ (.Y(_2447_),
    .B1(_2446_),
    .B2(net2591),
    .A2(_2122_),
    .A1(net2420));
 sg13g2_a21oi_1 _6810_ (.A1(_2124_),
    .A2(_2445_),
    .Y(_2448_),
    .B1(_2447_));
 sg13g2_a221oi_1 _6811_ (.B2(_3028_),
    .C1(net2520),
    .B1(_1674_),
    .A1(net2560),
    .Y(_2450_),
    .A2(_3044_));
 sg13g2_nor2_1 _6812_ (.A(net2402),
    .B(_1674_),
    .Y(_2451_));
 sg13g2_nor3_1 _6813_ (.A(net2461),
    .B(_2394_),
    .C(_1675_),
    .Y(_2452_));
 sg13g2_nor4_1 _6814_ (.A(net2199),
    .B(_2450_),
    .C(_2451_),
    .D(_2452_),
    .Y(_2453_));
 sg13g2_a21oi_1 _6815_ (.A1(net2196),
    .A2(_2448_),
    .Y(_2454_),
    .B1(_2453_));
 sg13g2_a21oi_2 _6816_ (.B1(_3375_),
    .Y(_2455_),
    .A2(_2454_),
    .A1(_2443_));
 sg13g2_a221oi_1 _6817_ (.B2(_2432_),
    .C1(_2455_),
    .B1(_2412_),
    .A1(_2381_),
    .Y(_2456_),
    .A2(_2393_));
 sg13g2_a22oi_1 _6818_ (.Y(_2457_),
    .B1(_2170_),
    .B2(net2566),
    .A2(_1154_),
    .A1(net2475));
 sg13g2_a21oi_1 _6819_ (.A1(_2171_),
    .A2(_2457_),
    .Y(_2458_),
    .B1(net2491));
 sg13g2_o21ai_1 _6820_ (.B1(net2589),
    .Y(_2459_),
    .A1(_3269_),
    .A2(_0229_));
 sg13g2_a21oi_1 _6821_ (.A1(_1156_),
    .A2(_2459_),
    .Y(_2461_),
    .B1(net2326));
 sg13g2_o21ai_1 _6822_ (.B1(net2565),
    .Y(_2462_),
    .A1(_3269_),
    .A2(_0229_));
 sg13g2_a21oi_1 _6823_ (.A1(_1384_),
    .A2(_2462_),
    .Y(_2463_),
    .B1(net2313));
 sg13g2_nor4_1 _6824_ (.A(net2394),
    .B(_2458_),
    .C(_2461_),
    .D(_2463_),
    .Y(_2464_));
 sg13g2_a21oi_1 _6825_ (.A1(net2566),
    .A2(net2021),
    .Y(_2465_),
    .B1(_3271_));
 sg13g2_nor3_1 _6826_ (.A(net2510),
    .B(_0153_),
    .C(_2465_),
    .Y(_2466_));
 sg13g2_nor3_1 _6827_ (.A(net2380),
    .B(_1750_),
    .C(_2466_),
    .Y(_2467_));
 sg13g2_o21ai_1 _6828_ (.B1(_3300_),
    .Y(_2468_),
    .A1(_2464_),
    .A2(_2467_));
 sg13g2_a221oi_1 _6829_ (.B2(net2069),
    .C1(_2075_),
    .B1(_1882_),
    .A1(net2584),
    .Y(_2469_),
    .A2(_1715_));
 sg13g2_nand2b_1 _6830_ (.Y(_2470_),
    .B(_1032_),
    .A_N(_2469_));
 sg13g2_a22oi_1 _6831_ (.Y(_2472_),
    .B1(_0273_),
    .B2(_2826_),
    .A2(_0257_),
    .A1(net2464));
 sg13g2_a221oi_1 _6832_ (.B2(net2105),
    .C1(_1363_),
    .B1(_2472_),
    .A1(net2463),
    .Y(_2473_),
    .A2(_0473_));
 sg13g2_a21o_1 _6833_ (.A2(_2473_),
    .A1(_2470_),
    .B1(net2490),
    .X(_2474_));
 sg13g2_o21ai_1 _6834_ (.B1(_3150_),
    .Y(_2475_),
    .A1(_0157_),
    .A2(_1336_));
 sg13g2_o21ai_1 _6835_ (.B1(_3349_),
    .Y(_2476_),
    .A1(net2597),
    .A2(_3127_));
 sg13g2_o21ai_1 _6836_ (.B1(net2320),
    .Y(_2477_),
    .A1(_2475_),
    .A2(_2476_));
 sg13g2_nor3_1 _6837_ (.A(net2258),
    .B(net2214),
    .C(net2212),
    .Y(_2478_));
 sg13g2_and2_1 _6838_ (.A(net2104),
    .B(_2478_),
    .X(_2479_));
 sg13g2_o21ai_1 _6839_ (.B1(net2104),
    .Y(_2480_),
    .A1(_3145_),
    .A2(_2478_));
 sg13g2_o21ai_1 _6840_ (.B1(net2152),
    .Y(_2481_),
    .A1(_3154_),
    .A2(_1715_));
 sg13g2_a21o_1 _6841_ (.A2(_2481_),
    .A1(_2480_),
    .B1(net2326),
    .X(_2483_));
 sg13g2_nand4_1 _6842_ (.B(_2474_),
    .C(_2477_),
    .A(net2393),
    .Y(_2484_),
    .D(_2483_));
 sg13g2_nand3_1 _6843_ (.B(net2092),
    .C(_3221_),
    .A(net2579),
    .Y(_2485_));
 sg13g2_a21oi_1 _6844_ (.A1(_2559_),
    .A2(net2217),
    .Y(_2486_),
    .B1(_2075_));
 sg13g2_o21ai_1 _6845_ (.B1(_2485_),
    .Y(_2487_),
    .A1(_3025_),
    .A2(_2486_));
 sg13g2_nand3_1 _6846_ (.B(net2453),
    .C(net2277),
    .A(net2586),
    .Y(_2488_));
 sg13g2_nand4_1 _6847_ (.B(net2079),
    .C(_3528_),
    .A(net2148),
    .Y(_2489_),
    .D(_2488_));
 sg13g2_a221oi_1 _6848_ (.B2(_3221_),
    .C1(net2148),
    .B1(net2080),
    .A1(net2451),
    .Y(_2490_),
    .A2(net2360));
 sg13g2_nor2_1 _6849_ (.A(net2313),
    .B(_2490_),
    .Y(_2491_));
 sg13g2_nor3_2 _6850_ (.A(net2178),
    .B(net2060),
    .C(_0168_),
    .Y(_2492_));
 sg13g2_nand3_1 _6851_ (.B(net2056),
    .C(_0169_),
    .A(net2126),
    .Y(_2494_));
 sg13g2_nand4_1 _6852_ (.B(_3586_),
    .C(_0664_),
    .A(net2027),
    .Y(_2495_),
    .D(_2494_));
 sg13g2_o21ai_1 _6853_ (.B1(net2333),
    .Y(_2496_),
    .A1(_2475_),
    .A2(_2479_));
 sg13g2_nand4_1 _6854_ (.B(_0664_),
    .C(_2373_),
    .A(net2027),
    .Y(_2497_),
    .D(_2480_));
 sg13g2_a22oi_1 _6855_ (.Y(_2498_),
    .B1(_2497_),
    .B2(net2340),
    .A2(_2495_),
    .A1(net2310));
 sg13g2_a22oi_1 _6856_ (.Y(_2499_),
    .B1(_2489_),
    .B2(_2491_),
    .A2(_2487_),
    .A1(net2328));
 sg13g2_nand4_1 _6857_ (.B(_2496_),
    .C(_2498_),
    .A(net2380),
    .Y(_2500_),
    .D(_2499_));
 sg13g2_a21oi_1 _6858_ (.A1(_2484_),
    .A2(_2500_),
    .Y(_2501_),
    .B1(net1981));
 sg13g2_nand2_1 _6859_ (.Y(_2502_),
    .A(_0784_),
    .B(_0951_));
 sg13g2_nor2_2 _6860_ (.A(_2853_),
    .B(_3607_),
    .Y(_2503_));
 sg13g2_a22oi_1 _6861_ (.Y(_2505_),
    .B1(_2503_),
    .B2(net2506),
    .A2(_2502_),
    .A1(net2339));
 sg13g2_nand3_1 _6862_ (.B(net2101),
    .C(_3542_),
    .A(net2473),
    .Y(_2506_));
 sg13g2_o21ai_1 _6863_ (.B1(_2506_),
    .Y(_2507_),
    .A1(net2563),
    .A2(_3045_));
 sg13g2_o21ai_1 _6864_ (.B1(_1322_),
    .Y(_2508_),
    .A1(net2586),
    .A2(_1336_));
 sg13g2_a22oi_1 _6865_ (.Y(_2509_),
    .B1(_2508_),
    .B2(net2332),
    .A2(_2211_),
    .A1(_3061_));
 sg13g2_a22oi_1 _6866_ (.Y(_2510_),
    .B1(_2507_),
    .B2(net2489),
    .A2(_1330_),
    .A1(net2328));
 sg13g2_nand3_1 _6867_ (.B(_2509_),
    .C(_2510_),
    .A(_2505_),
    .Y(_2511_));
 sg13g2_a21oi_1 _6868_ (.A1(net2024),
    .A2(_0227_),
    .Y(_2512_),
    .B1(net2567));
 sg13g2_o21ai_1 _6869_ (.B1(net2547),
    .Y(_2513_),
    .A1(_1334_),
    .A2(_2512_));
 sg13g2_nand3b_1 _6870_ (.B(_2215_),
    .C(_2513_),
    .Y(_2514_),
    .A_N(_2214_));
 sg13g2_a221oi_1 _6871_ (.B2(net2563),
    .C1(_1762_),
    .B1(_3054_),
    .A1(net2101),
    .Y(_2516_),
    .A2(net2080));
 sg13g2_a21oi_1 _6872_ (.A1(_3289_),
    .A2(_1764_),
    .Y(_2517_),
    .B1(net1983));
 sg13g2_o21ai_1 _6873_ (.B1(_2517_),
    .Y(_2518_),
    .A1(_3460_),
    .A2(_2516_));
 sg13g2_a221oi_1 _6874_ (.B2(net2203),
    .C1(_2518_),
    .B1(_2514_),
    .A1(net2378),
    .Y(_2519_),
    .A2(_2511_));
 sg13g2_nor3_1 _6875_ (.A(net1977),
    .B(_2501_),
    .C(_2519_),
    .Y(_2520_));
 sg13g2_a21oi_1 _6876_ (.A1(_2468_),
    .A2(_2520_),
    .Y(_2521_),
    .B1(net1976));
 sg13g2_o21ai_1 _6877_ (.B1(_2521_),
    .Y(_2522_),
    .A1(net1978),
    .A2(_2456_));
 sg13g2_o21ai_1 _6878_ (.B1(_1482_),
    .Y(_2523_),
    .A1(_0429_),
    .A2(_1484_));
 sg13g2_o21ai_1 _6879_ (.B1(net2324),
    .Y(_2524_),
    .A1(net1987),
    .A2(_2492_));
 sg13g2_a21oi_1 _6880_ (.A1(_1065_),
    .A2(_1482_),
    .Y(_2525_),
    .B1(_2343_));
 sg13g2_a221oi_1 _6881_ (.B2(_3419_),
    .C1(_2525_),
    .B1(_2523_),
    .A1(net2082),
    .Y(_2527_),
    .A2(net2307));
 sg13g2_a21o_1 _6882_ (.A2(_2527_),
    .A1(_2524_),
    .B1(net2383),
    .X(_2528_));
 sg13g2_a21oi_2 _6883_ (.B1(net2127),
    .Y(_2529_),
    .A2(_3102_),
    .A1(_2064_));
 sg13g2_nor2_1 _6884_ (.A(net2308),
    .B(_2529_),
    .Y(_2530_));
 sg13g2_o21ai_1 _6885_ (.B1(_3102_),
    .Y(_2531_),
    .A1(net2083),
    .A2(net2239));
 sg13g2_a221oi_1 _6886_ (.B2(_1032_),
    .C1(net2497),
    .B1(_2531_),
    .A1(net2553),
    .Y(_2532_),
    .A2(net1987));
 sg13g2_a21oi_1 _6887_ (.A1(net2480),
    .A2(_2529_),
    .Y(_2533_),
    .B1(_2492_));
 sg13g2_o21ai_1 _6888_ (.B1(_2533_),
    .Y(_2534_),
    .A1(_2530_),
    .A2(_2532_));
 sg13g2_and3_1 _6889_ (.X(_2535_),
    .A(_0094_),
    .B(_0418_),
    .C(_2494_));
 sg13g2_a21oi_1 _6890_ (.A1(_0561_),
    .A2(_2535_),
    .Y(_2536_),
    .B1(net2397));
 sg13g2_a21oi_1 _6891_ (.A1(_2534_),
    .A2(_2536_),
    .Y(_2538_),
    .B1(net2303));
 sg13g2_o21ai_1 _6892_ (.B1(net2533),
    .Y(_2539_),
    .A1(net1987),
    .A2(_2492_));
 sg13g2_o21ai_1 _6893_ (.B1(net2553),
    .Y(_2540_),
    .A1(net1987),
    .A2(_2389_));
 sg13g2_nand3_1 _6894_ (.B(_2539_),
    .C(_2540_),
    .A(_2000_),
    .Y(_2541_));
 sg13g2_or3_1 _6895_ (.A(_3131_),
    .B(_0434_),
    .C(_1450_),
    .X(_2542_));
 sg13g2_nand4_1 _6896_ (.B(net1998),
    .C(_0640_),
    .A(_3395_),
    .Y(_2543_),
    .D(_1451_));
 sg13g2_a22oi_1 _6897_ (.Y(_2544_),
    .B1(_2543_),
    .B2(net2480),
    .A2(_2542_),
    .A1(net2342));
 sg13g2_nand2b_1 _6898_ (.Y(_2545_),
    .B(_0124_),
    .A_N(_2544_));
 sg13g2_and2_1 _6899_ (.A(_1507_),
    .B(_2523_),
    .X(_2546_));
 sg13g2_or3_1 _6900_ (.A(_3131_),
    .B(_0434_),
    .C(net1987),
    .X(_2547_));
 sg13g2_a21o_1 _6901_ (.A2(_2547_),
    .A1(_0122_),
    .B1(net2296),
    .X(_2549_));
 sg13g2_a221oi_1 _6902_ (.B2(net2386),
    .C1(_2549_),
    .B1(_2546_),
    .A1(net2205),
    .Y(_2550_),
    .A2(_2541_));
 sg13g2_a221oi_1 _6903_ (.B2(_2550_),
    .C1(net2036),
    .B1(_2545_),
    .A1(_2528_),
    .Y(_2551_),
    .A2(_2538_));
 sg13g2_nor2_1 _6904_ (.A(net2594),
    .B(net2067),
    .Y(_2552_));
 sg13g2_o21ai_1 _6905_ (.B1(_0101_),
    .Y(_2553_),
    .A1(_1956_),
    .A2(_2552_));
 sg13g2_a21oi_1 _6906_ (.A1(_1227_),
    .A2(_1401_),
    .Y(_2554_),
    .B1(net2529));
 sg13g2_a221oi_1 _6907_ (.B2(_3297_),
    .C1(_2554_),
    .B1(_2553_),
    .A1(net2529),
    .Y(_2555_),
    .A2(_3567_));
 sg13g2_a21oi_1 _6908_ (.A1(_3566_),
    .A2(_0743_),
    .Y(_2556_),
    .B1(net2434));
 sg13g2_a221oi_1 _6909_ (.B2(_3343_),
    .C1(net2418),
    .B1(_1616_),
    .A1(net2061),
    .Y(_2557_),
    .A2(_0216_));
 sg13g2_mux4_1 _6910_ (.S0(net2113),
    .A0(_3007_),
    .A1(net2215),
    .A2(_3163_),
    .A3(_3421_),
    .S1(net2284),
    .X(_2558_));
 sg13g2_nor2_1 _6911_ (.A(net2405),
    .B(_2558_),
    .Y(_2560_));
 sg13g2_nor3_1 _6912_ (.A(_2425_),
    .B(_2556_),
    .C(_2560_),
    .Y(_2561_));
 sg13g2_nor3_1 _6913_ (.A(net2512),
    .B(_2237_),
    .C(_2557_),
    .Y(_2562_));
 sg13g2_o21ai_1 _6914_ (.B1(net2514),
    .Y(_2563_),
    .A1(net2466),
    .A2(_0639_));
 sg13g2_o21ai_1 _6915_ (.B1(net2343),
    .Y(_2564_),
    .A1(_0513_),
    .A2(_0638_));
 sg13g2_nor3_1 _6916_ (.A(net2465),
    .B(_3231_),
    .C(net2001),
    .Y(_2565_));
 sg13g2_nor3_1 _6917_ (.A(_2245_),
    .B(_2563_),
    .C(_2565_),
    .Y(_2566_));
 sg13g2_nand2_1 _6918_ (.Y(_2567_),
    .A(_3156_),
    .B(net2016));
 sg13g2_o21ai_1 _6919_ (.B1(net2494),
    .Y(_2568_),
    .A1(net2435),
    .A2(_3528_));
 sg13g2_a22oi_1 _6920_ (.Y(_2569_),
    .B1(_2567_),
    .B2(net2412),
    .A2(_0754_),
    .A1(net2550));
 sg13g2_nor3_1 _6921_ (.A(net2551),
    .B(_3380_),
    .C(_1432_),
    .Y(_2571_));
 sg13g2_nor3_1 _6922_ (.A(_0732_),
    .B(_2568_),
    .C(_2571_),
    .Y(_2572_));
 sg13g2_a221oi_1 _6923_ (.B2(_2562_),
    .C1(net2396),
    .B1(_2561_),
    .A1(_2232_),
    .Y(_2573_),
    .A2(_2555_));
 sg13g2_a221oi_1 _6924_ (.B2(_2572_),
    .C1(net2382),
    .B1(_2569_),
    .A1(_2564_),
    .Y(_2574_),
    .A2(_2566_));
 sg13g2_o21ai_1 _6925_ (.B1(net1984),
    .Y(_2575_),
    .A1(_2573_),
    .A2(_2574_));
 sg13g2_nand3_1 _6926_ (.B(net2004),
    .C(_1053_),
    .A(net2019),
    .Y(_2576_));
 sg13g2_o21ai_1 _6927_ (.B1(net2329),
    .Y(_2577_),
    .A1(_0325_),
    .A2(_2576_));
 sg13g2_a22oi_1 _6928_ (.Y(_2578_),
    .B1(_2278_),
    .B2(net2321),
    .A2(_0838_),
    .A1(net2311));
 sg13g2_a21oi_1 _6929_ (.A1(net2019),
    .A2(net2003),
    .Y(_2579_),
    .B1(net2342));
 sg13g2_nand2_1 _6930_ (.Y(_2580_),
    .A(net2342),
    .B(net2227));
 sg13g2_o21ai_1 _6931_ (.B1(_1451_),
    .Y(_2582_),
    .A1(net1989),
    .A2(_2580_));
 sg13g2_o21ai_1 _6932_ (.B1(net2517),
    .Y(_2583_),
    .A1(_2579_),
    .A2(_2582_));
 sg13g2_nand4_1 _6933_ (.B(_2577_),
    .C(_2578_),
    .A(net2386),
    .Y(_2584_),
    .D(_2583_));
 sg13g2_nand3_1 _6934_ (.B(net1998),
    .C(_1451_),
    .A(net2019),
    .Y(_2585_));
 sg13g2_o21ai_1 _6935_ (.B1(net2324),
    .Y(_2586_),
    .A1(_0333_),
    .A2(_2585_));
 sg13g2_a21oi_1 _6936_ (.A1(net2213),
    .A2(net2013),
    .Y(_2587_),
    .B1(_0514_));
 sg13g2_o21ai_1 _6937_ (.B1(net2398),
    .Y(_2588_),
    .A1(_1456_),
    .A2(_2343_));
 sg13g2_a221oi_1 _6938_ (.B2(net2340),
    .C1(_2588_),
    .B1(_2587_),
    .A1(_1551_),
    .Y(_2589_),
    .A2(_2529_));
 sg13g2_o21ai_1 _6939_ (.B1(net2329),
    .Y(_2590_),
    .A1(_0324_),
    .A2(_1066_));
 sg13g2_nand2b_1 _6940_ (.Y(_2591_),
    .B(net2335),
    .A_N(_2535_));
 sg13g2_nand4_1 _6941_ (.B(_2589_),
    .C(_2590_),
    .A(_2586_),
    .Y(_2593_),
    .D(_2591_));
 sg13g2_nand3_1 _6942_ (.B(_2584_),
    .C(_2593_),
    .A(_3300_),
    .Y(_2594_));
 sg13g2_nand3b_1 _6943_ (.B(_2575_),
    .C(_2594_),
    .Y(_2595_),
    .A_N(_2551_));
 sg13g2_a221oi_1 _6944_ (.B2(net2142),
    .C1(_3149_),
    .B1(_0398_),
    .A1(_2647_),
    .Y(_2596_),
    .A2(_3326_));
 sg13g2_nand2b_1 _6945_ (.Y(_2597_),
    .B(net2408),
    .A_N(_2596_));
 sg13g2_a221oi_1 _6946_ (.B2(_3153_),
    .C1(_3091_),
    .B1(net2062),
    .A1(_2570_),
    .Y(_2598_),
    .A2(_2948_));
 sg13g2_a21oi_1 _6947_ (.A1(_2816_),
    .A2(net2055),
    .Y(_2599_),
    .B1(net2063));
 sg13g2_o21ai_1 _6948_ (.B1(_2321_),
    .Y(_2600_),
    .A1(_3253_),
    .A2(_2599_));
 sg13g2_o21ai_1 _6949_ (.B1(net2542),
    .Y(_2601_),
    .A1(_2598_),
    .A2(_2600_));
 sg13g2_o21ai_1 _6950_ (.B1(net2472),
    .Y(_2602_),
    .A1(_0641_),
    .A2(_2315_));
 sg13g2_nand4_1 _6951_ (.B(_2597_),
    .C(_2601_),
    .A(net2485),
    .Y(_2604_),
    .D(_2602_));
 sg13g2_a21oi_1 _6952_ (.A1(net2112),
    .A2(net2072),
    .Y(_2605_),
    .B1(net2593));
 sg13g2_nand4_1 _6953_ (.B(_0720_),
    .C(_2034_),
    .A(net2027),
    .Y(_2606_),
    .D(_2605_));
 sg13g2_nand3_1 _6954_ (.B(_1019_),
    .C(_1531_),
    .A(net2026),
    .Y(_2607_));
 sg13g2_nand3_1 _6955_ (.B(_2606_),
    .C(_2607_),
    .A(net2548),
    .Y(_2608_));
 sg13g2_o21ai_1 _6956_ (.B1(net2410),
    .Y(_2609_),
    .A1(_1533_),
    .A2(_1538_));
 sg13g2_a21oi_1 _6957_ (.A1(_3130_),
    .A2(_0687_),
    .Y(_2610_),
    .B1(net2466));
 sg13g2_a21oi_1 _6958_ (.A1(_2319_),
    .A2(_2610_),
    .Y(_2611_),
    .B1(net2493));
 sg13g2_nand3_1 _6959_ (.B(_2609_),
    .C(_2611_),
    .A(_2608_),
    .Y(_2612_));
 sg13g2_a21oi_1 _6960_ (.A1(_2604_),
    .A2(_2612_),
    .Y(_2613_),
    .B1(net2377));
 sg13g2_o21ai_1 _6961_ (.B1(net2033),
    .Y(_2615_),
    .A1(_2787_),
    .A2(_1424_));
 sg13g2_nor2_1 _6962_ (.A(net2034),
    .B(_0375_),
    .Y(_2616_));
 sg13g2_a21oi_1 _6963_ (.A1(_2615_),
    .A2(_2616_),
    .Y(_2617_),
    .B1(net2314));
 sg13g2_nor2_1 _6964_ (.A(net2561),
    .B(_0288_),
    .Y(_2618_));
 sg13g2_o21ai_1 _6965_ (.B1(net2334),
    .Y(_2619_),
    .A1(_2315_),
    .A2(_2618_));
 sg13g2_o21ai_1 _6966_ (.B1(net2559),
    .Y(_2620_),
    .A1(net2090),
    .A2(_2251_));
 sg13g2_a21oi_1 _6967_ (.A1(net2521),
    .A2(_3191_),
    .Y(_2621_),
    .B1(_2328_));
 sg13g2_o21ai_1 _6968_ (.B1(_2619_),
    .Y(_2622_),
    .A1(net2483),
    .A2(_2621_));
 sg13g2_nand2_1 _6969_ (.Y(_2623_),
    .A(_0880_),
    .B(_2620_));
 sg13g2_a21oi_1 _6970_ (.A1(_3192_),
    .A2(_2623_),
    .Y(_2624_),
    .B1(net2325));
 sg13g2_nor4_1 _6971_ (.A(net2388),
    .B(_2617_),
    .C(_2622_),
    .D(_2624_),
    .Y(_2626_));
 sg13g2_o21ai_1 _6972_ (.B1(net1982),
    .Y(_2627_),
    .A1(_2613_),
    .A2(_2626_));
 sg13g2_o21ai_1 _6973_ (.B1(net2333),
    .Y(_2628_),
    .A1(_3269_),
    .A2(_0229_));
 sg13g2_o21ai_1 _6974_ (.B1(_2628_),
    .Y(_2629_),
    .A1(net2336),
    .A2(_1153_));
 sg13g2_a21o_1 _6975_ (.A2(_2170_),
    .A1(net2491),
    .B1(_2629_),
    .X(_2630_));
 sg13g2_o21ai_1 _6976_ (.B1(net2381),
    .Y(_2631_),
    .A1(_1158_),
    .A2(_2630_));
 sg13g2_nand2_1 _6977_ (.Y(_2632_),
    .A(net2432),
    .B(_1563_));
 sg13g2_o21ai_1 _6978_ (.B1(net2565),
    .Y(_2633_),
    .A1(net2020),
    .A2(_1616_));
 sg13g2_a21oi_1 _6979_ (.A1(_2632_),
    .A2(_2633_),
    .Y(_2634_),
    .B1(net2201));
 sg13g2_a21oi_1 _6980_ (.A1(_0685_),
    .A2(_1384_),
    .Y(_2635_),
    .B1(_3460_));
 sg13g2_nor4_1 _6981_ (.A(net1985),
    .B(_2332_),
    .C(_2634_),
    .D(_2635_),
    .Y(_2637_));
 sg13g2_nor2_1 _6982_ (.A(net2199),
    .B(_3271_),
    .Y(_2638_));
 sg13g2_a221oi_1 _6983_ (.B2(_2063_),
    .C1(net1979),
    .B1(_2638_),
    .A1(_2631_),
    .Y(_2639_),
    .A2(_2637_));
 sg13g2_nor3_1 _6984_ (.A(net2563),
    .B(_0230_),
    .C(_0736_),
    .Y(_2640_));
 sg13g2_o21ai_1 _6985_ (.B1(net2520),
    .Y(_2641_),
    .A1(_2334_),
    .A2(_2640_));
 sg13g2_a221oi_1 _6986_ (.B2(_1585_),
    .C1(_3089_),
    .B1(_1122_),
    .A1(net2471),
    .Y(_2642_),
    .A2(_3030_));
 sg13g2_a21o_1 _6987_ (.A2(_2642_),
    .A1(_2641_),
    .B1(net2199),
    .X(_2643_));
 sg13g2_and2_1 _6988_ (.A(net2338),
    .B(_1192_),
    .X(_2644_));
 sg13g2_nor2_1 _6989_ (.A(net2330),
    .B(_2347_),
    .Y(_2645_));
 sg13g2_o21ai_1 _6990_ (.B1(_0773_),
    .Y(_2646_),
    .A1(_2644_),
    .A2(_2645_));
 sg13g2_a21oi_1 _6991_ (.A1(net2544),
    .A2(_3056_),
    .Y(_2648_),
    .B1(net2506));
 sg13g2_nand2_1 _6992_ (.Y(_2649_),
    .A(_0271_),
    .B(_2648_));
 sg13g2_o21ai_1 _6993_ (.B1(net2379),
    .Y(_2650_),
    .A1(_3229_),
    .A2(_2649_));
 sg13g2_nand2b_1 _6994_ (.Y(_2651_),
    .B(_2646_),
    .A_N(_2650_));
 sg13g2_nand4_1 _6995_ (.B(_3032_),
    .C(_0206_),
    .A(net2539),
    .Y(_2652_),
    .D(_1179_));
 sg13g2_o21ai_1 _6996_ (.B1(_0522_),
    .Y(_2653_),
    .A1(_3293_),
    .A2(_1038_));
 sg13g2_nand3_1 _6997_ (.B(_2652_),
    .C(_2653_),
    .A(net2196),
    .Y(_2654_));
 sg13g2_nand4_1 _6998_ (.B(_2643_),
    .C(_2651_),
    .A(_3431_),
    .Y(_2655_),
    .D(_2654_));
 sg13g2_nand3_1 _6999_ (.B(_2639_),
    .C(_2655_),
    .A(_2627_),
    .Y(_2656_));
 sg13g2_a21oi_1 _7000_ (.A1(net1980),
    .A2(_2595_),
    .Y(_2657_),
    .B1(_3308_));
 sg13g2_a21oi_1 _7001_ (.A1(_2656_),
    .A2(_2657_),
    .Y(_2659_),
    .B1(_3505_));
 sg13g2_a21oi_1 _7002_ (.A1(_2522_),
    .A2(_2659_),
    .Y(_2660_),
    .B1(_1085_));
 sg13g2_a221oi_1 _7003_ (.B2(_2660_),
    .C1(_0616_),
    .B1(_2356_),
    .A1(_1085_),
    .Y(_2661_),
    .A2(_2070_));
 sg13g2_nand2_1 _7004_ (.Y(_2662_),
    .A(\logo_top[8] ),
    .B(_0790_));
 sg13g2_xnor2_1 _7005_ (.Y(_2663_),
    .A(\logo_top[8] ),
    .B(\pix_y[8] ));
 sg13g2_a21oi_2 _7006_ (.B1(_3307_),
    .Y(_2664_),
    .A2(\pix_y[7] ),
    .A1(_0680_));
 sg13g2_nand2_1 _7007_ (.Y(_2665_),
    .A(\logo_left[8] ),
    .B(_0779_));
 sg13g2_xnor2_1 _7008_ (.Y(_2666_),
    .A(\logo_left[8] ),
    .B(\pix_x[8] ));
 sg13g2_nand3_1 _7009_ (.B(_1624_),
    .C(_2666_),
    .A(_1382_),
    .Y(_2667_));
 sg13g2_xnor2_1 _7010_ (.Y(_2668_),
    .A(\logo_left[9] ),
    .B(\pix_x[9] ));
 sg13g2_xnor2_1 _7011_ (.Y(_2670_),
    .A(_2665_),
    .B(_2668_));
 sg13g2_xnor2_1 _7012_ (.Y(_2671_),
    .A(\logo_top[9] ),
    .B(\pix_y[9] ));
 sg13g2_xnor2_1 _7013_ (.Y(_2672_),
    .A(_2662_),
    .B(_2671_));
 sg13g2_a21oi_1 _7014_ (.A1(_1382_),
    .A2(_1624_),
    .Y(_2673_),
    .B1(_2666_));
 sg13g2_a21oi_1 _7015_ (.A1(_2663_),
    .A2(_2664_),
    .Y(_2674_),
    .B1(_2673_));
 sg13g2_and4_1 _7016_ (.A(_2667_),
    .B(_2670_),
    .C(_2672_),
    .D(_2674_),
    .X(_2675_));
 sg13g2_o21ai_1 _7017_ (.B1(_2675_),
    .Y(_2676_),
    .A1(_2663_),
    .A2(_2664_));
 sg13g2_a221oi_1 _7018_ (.B2(_0933_),
    .C1(_2661_),
    .B1(_2676_),
    .A1(_0614_),
    .Y(_2677_),
    .A2(_1400_));
 sg13g2_nand2_1 _7019_ (.Y(_2678_),
    .A(net2606),
    .B(\frame_counter[5] ));
 sg13g2_xnor2_1 _7020_ (.Y(_2679_),
    .A(net2606),
    .B(\frame_counter[5] ));
 sg13g2_nand2_1 _7021_ (.Y(_2681_),
    .A(net2607),
    .B(\frame_counter[4] ));
 sg13g2_or2_1 _7022_ (.X(_2682_),
    .B(\frame_counter[2] ),
    .A(net2611));
 sg13g2_nor2_1 _7023_ (.A(\pix_y[1] ),
    .B(\frame_counter[1] ),
    .Y(_2683_));
 sg13g2_nand2_1 _7024_ (.Y(_2684_),
    .A(\frame_counter[0] ),
    .B(net2613));
 sg13g2_a22oi_1 _7025_ (.Y(_2685_),
    .B1(\frame_counter[1] ),
    .B2(\pix_y[1] ),
    .A2(\frame_counter[2] ),
    .A1(net2611));
 sg13g2_o21ai_1 _7026_ (.B1(_2685_),
    .Y(_2686_),
    .A1(_2683_),
    .A2(_2684_));
 sg13g2_a22oi_1 _7027_ (.Y(_2687_),
    .B1(_2682_),
    .B2(_2686_),
    .A2(\frame_counter[3] ),
    .A1(net2609));
 sg13g2_or2_1 _7028_ (.X(_2688_),
    .B(\frame_counter[4] ),
    .A(net2607));
 sg13g2_o21ai_1 _7029_ (.B1(_2688_),
    .Y(_2689_),
    .A1(net2609),
    .A2(\frame_counter[3] ));
 sg13g2_o21ai_1 _7030_ (.B1(_2681_),
    .Y(_2690_),
    .A1(_2687_),
    .A2(_2689_));
 sg13g2_nand2b_1 _7031_ (.Y(_2692_),
    .B(_2690_),
    .A_N(_2679_));
 sg13g2_xnor2_1 _7032_ (.Y(_2693_),
    .A(_2679_),
    .B(_2690_));
 sg13g2_nand2_1 _7033_ (.Y(_2694_),
    .A(net2621),
    .B(\frame_counter[5] ));
 sg13g2_xor2_1 _7034_ (.B(\frame_counter[5] ),
    .A(net2621),
    .X(_2695_));
 sg13g2_or2_1 _7035_ (.X(_2696_),
    .B(\frame_counter[4] ),
    .A(\pix_x[4] ));
 sg13g2_nor2_1 _7036_ (.A(\pix_x[1] ),
    .B(\frame_counter[1] ),
    .Y(_2697_));
 sg13g2_nand2_1 _7037_ (.Y(_2698_),
    .A(\frame_counter[0] ),
    .B(\pix_x[0] ));
 sg13g2_a22oi_1 _7038_ (.Y(_2699_),
    .B1(\frame_counter[1] ),
    .B2(\pix_x[1] ),
    .A2(\frame_counter[2] ),
    .A1(\pix_x[2] ));
 sg13g2_o21ai_1 _7039_ (.B1(_2699_),
    .Y(_2700_),
    .A1(_2697_),
    .A2(_2698_));
 sg13g2_nor2_1 _7040_ (.A(\pix_x[3] ),
    .B(\frame_counter[3] ),
    .Y(_2701_));
 sg13g2_o21ai_1 _7041_ (.B1(_2700_),
    .Y(_2703_),
    .A1(\pix_x[2] ),
    .A2(\frame_counter[2] ));
 sg13g2_a22oi_1 _7042_ (.Y(_2704_),
    .B1(\frame_counter[3] ),
    .B2(\pix_x[3] ),
    .A2(\frame_counter[4] ),
    .A1(\pix_x[4] ));
 sg13g2_o21ai_1 _7043_ (.B1(_2704_),
    .Y(_2705_),
    .A1(_2701_),
    .A2(_2703_));
 sg13g2_nand3_1 _7044_ (.B(_2696_),
    .C(_2705_),
    .A(_2695_),
    .Y(_2706_));
 sg13g2_a21o_1 _7045_ (.A2(_2705_),
    .A1(_2696_),
    .B1(_2695_),
    .X(_2707_));
 sg13g2_and2_1 _7046_ (.A(_2706_),
    .B(_2707_),
    .X(_2708_));
 sg13g2_xnor2_1 _7047_ (.Y(_2709_),
    .A(net2604),
    .B(net2620));
 sg13g2_xnor2_1 _7048_ (.Y(_2710_),
    .A(_2708_),
    .B(_2709_));
 sg13g2_xnor2_1 _7049_ (.Y(_2711_),
    .A(_2693_),
    .B(_2710_));
 sg13g2_xnor2_1 _7050_ (.Y(_2712_),
    .A(net2620),
    .B(\frame_counter[6] ));
 sg13g2_a21oi_1 _7051_ (.A1(_2694_),
    .A2(_2706_),
    .Y(_2714_),
    .B1(_2712_));
 sg13g2_nand3_1 _7052_ (.B(_2706_),
    .C(_2712_),
    .A(_2694_),
    .Y(_2715_));
 sg13g2_nor2b_1 _7053_ (.A(_2714_),
    .B_N(_2715_),
    .Y(_2716_));
 sg13g2_xnor2_1 _7054_ (.Y(_2717_),
    .A(\pix_y[7] ),
    .B(_2716_));
 sg13g2_xnor2_1 _7055_ (.Y(_2718_),
    .A(_2711_),
    .B(_2717_));
 sg13g2_nor2_1 _7056_ (.A(_2677_),
    .B(_2718_),
    .Y(_2719_));
 sg13g2_nand4_1 _7057_ (.B(\pix_y[7] ),
    .C(net2603),
    .A(\pix_y[8] ),
    .Y(_2720_),
    .D(net2605));
 sg13g2_nor2_1 _7058_ (.A(\pix_y[9] ),
    .B(net2622),
    .Y(_2721_));
 sg13g2_o21ai_1 _7059_ (.B1(\pix_x[9] ),
    .Y(_2722_),
    .A1(\pix_x[8] ),
    .A2(net2619));
 sg13g2_nand3_1 _7060_ (.B(_2721_),
    .C(_2722_),
    .A(_2720_),
    .Y(_2723_));
 sg13g2_nor2_1 _7061_ (.A(net141),
    .B(_0944_),
    .Y(_2725_));
 sg13g2_nor3_1 _7062_ (.A(net186),
    .B(\color_index[0] ),
    .C(_0944_),
    .Y(_2726_));
 sg13g2_and2_1 _7063_ (.A(_2677_),
    .B(_2726_),
    .X(_2727_));
 sg13g2_nor3_1 _7064_ (.A(_2719_),
    .B(_2723_),
    .C(_2727_),
    .Y(_0015_));
 sg13g2_xnor2_1 _7065_ (.Y(_2728_),
    .A(\pix_y[8] ),
    .B(\frame_counter[7] ));
 sg13g2_xnor2_1 _7066_ (.Y(_2729_),
    .A(net2619),
    .B(_2728_));
 sg13g2_a21oi_1 _7067_ (.A1(net2620),
    .A2(\frame_counter[6] ),
    .Y(_2730_),
    .B1(_2714_));
 sg13g2_xnor2_1 _7068_ (.Y(_2731_),
    .A(_2729_),
    .B(_2730_));
 sg13g2_xnor2_1 _7069_ (.Y(_2732_),
    .A(_2711_),
    .B(_2731_));
 sg13g2_nand2_1 _7070_ (.Y(_2733_),
    .A(net141),
    .B(\color_index[0] ));
 sg13g2_xor2_1 _7071_ (.B(\color_index[0] ),
    .A(\color_index[2] ),
    .X(_2735_));
 sg13g2_nor3_1 _7072_ (.A(net185),
    .B(_0944_),
    .C(_2735_),
    .Y(_2736_));
 sg13g2_mux2_1 _7073_ (.A0(_2732_),
    .A1(_2736_),
    .S(_2677_),
    .X(_2737_));
 sg13g2_nor2_1 _7074_ (.A(_2723_),
    .B(_2737_),
    .Y(_0016_));
 sg13g2_and3_1 _7075_ (.X(_2738_),
    .A(\pix_x[0] ),
    .B(net187),
    .C(net132));
 sg13g2_and2_1 _7076_ (.A(net161),
    .B(_2738_),
    .X(_2739_));
 sg13g2_and2_2 _7077_ (.A(\pix_x[4] ),
    .B(_2739_),
    .X(_2740_));
 sg13g2_nor4_2 _7078_ (.A(net182),
    .B(net2620),
    .C(net2621),
    .Y(_2741_),
    .D(_2722_));
 sg13g2_nand2_2 _7079_ (.Y(_2742_),
    .A(_2740_),
    .B(_2741_));
 sg13g2_a21oi_2 _7080_ (.B1(net2622),
    .Y(_2743_),
    .A2(_2741_),
    .A1(_2740_));
 sg13g2_nand2_1 _7081_ (.Y(_2745_),
    .A(net2626),
    .B(_2742_));
 sg13g2_and2_1 _7082_ (.A(net93),
    .B(_2743_),
    .X(_0017_));
 sg13g2_xnor2_1 _7083_ (.Y(_2746_),
    .A(\pix_x[0] ),
    .B(net145));
 sg13g2_nor2_1 _7084_ (.A(net2304),
    .B(net146),
    .Y(_0018_));
 sg13g2_a21oi_1 _7085_ (.A1(\pix_x[0] ),
    .A2(\pix_x[1] ),
    .Y(_2747_),
    .B1(net132));
 sg13g2_nor3_1 _7086_ (.A(_0878_),
    .B(_2738_),
    .C(net133),
    .Y(_0019_));
 sg13g2_o21ai_1 _7087_ (.B1(net2628),
    .Y(_2748_),
    .A1(net161),
    .A2(_2738_));
 sg13g2_nor2_1 _7088_ (.A(_2739_),
    .B(net162),
    .Y(_0020_));
 sg13g2_o21ai_1 _7089_ (.B1(net2629),
    .Y(_2749_),
    .A1(net172),
    .A2(_2739_));
 sg13g2_nor2_1 _7090_ (.A(_2740_),
    .B(_2749_),
    .Y(_0021_));
 sg13g2_o21ai_1 _7091_ (.B1(_2743_),
    .Y(_2751_),
    .A1(net2621),
    .A2(_2740_));
 sg13g2_a21oi_1 _7092_ (.A1(net2621),
    .A2(_2740_),
    .Y(_0022_),
    .B1(_2751_));
 sg13g2_a21oi_1 _7093_ (.A1(net2621),
    .A2(_2740_),
    .Y(_2752_),
    .B1(net2620));
 sg13g2_nor2b_2 _7094_ (.A(_1009_),
    .B_N(_2739_),
    .Y(_2753_));
 sg13g2_nor3_1 _7095_ (.A(net2304),
    .B(_2752_),
    .C(_2753_),
    .Y(_0023_));
 sg13g2_xnor2_1 _7096_ (.Y(_2754_),
    .A(net2619),
    .B(_2753_));
 sg13g2_nor2_1 _7097_ (.A(_2745_),
    .B(_2754_),
    .Y(_0024_));
 sg13g2_nand3_1 _7098_ (.B(net2619),
    .C(_2753_),
    .A(\pix_x[8] ),
    .Y(_2755_));
 sg13g2_a21o_1 _7099_ (.A2(_2753_),
    .A1(net159),
    .B1(\pix_x[8] ),
    .X(_2756_));
 sg13g2_and3_1 _7100_ (.X(_0025_),
    .A(_2743_),
    .B(_2755_),
    .C(net160));
 sg13g2_xor2_1 _7101_ (.B(_2755_),
    .A(net134),
    .X(_2758_));
 sg13g2_nor2_1 _7102_ (.A(net2304),
    .B(net135),
    .Y(_0026_));
 sg13g2_nand2b_1 _7103_ (.Y(_2759_),
    .B(net2613),
    .A_N(\prev_y[0] ));
 sg13g2_nand2b_1 _7104_ (.Y(_2760_),
    .B(net2607),
    .A_N(\prev_y[4] ));
 sg13g2_nand2b_1 _7105_ (.Y(_2761_),
    .B(net2610),
    .A_N(\prev_y[2] ));
 sg13g2_a22oi_1 _7106_ (.Y(_2762_),
    .B1(\prev_y[8] ),
    .B2(_0790_),
    .A2(\prev_y[0] ),
    .A1(_0867_));
 sg13g2_xor2_1 _7107_ (.B(\prev_y[9] ),
    .A(\pix_y[9] ),
    .X(_2763_));
 sg13g2_xor2_1 _7108_ (.B(\prev_y[3] ),
    .A(net2608),
    .X(_2764_));
 sg13g2_o21ai_1 _7109_ (.B1(_2759_),
    .Y(_2765_),
    .A1(_0812_),
    .A2(\prev_y[7] ));
 sg13g2_xor2_1 _7110_ (.B(\prev_y[5] ),
    .A(net2605),
    .X(_2766_));
 sg13g2_nor4_2 _7111_ (.A(_2763_),
    .B(_2764_),
    .C(_2765_),
    .Y(_2768_),
    .D(_2766_));
 sg13g2_a22oi_1 _7112_ (.Y(_2769_),
    .B1(_0911_),
    .B2(\pix_y[8] ),
    .A2(\prev_y[1] ),
    .A1(_0856_));
 sg13g2_a22oi_1 _7113_ (.Y(_2770_),
    .B1(\prev_y[6] ),
    .B2(_0823_),
    .A2(\prev_y[4] ),
    .A1(_0834_));
 sg13g2_nand4_1 _7114_ (.B(_2761_),
    .C(_2762_),
    .A(_2760_),
    .Y(_2771_),
    .D(_2770_));
 sg13g2_a221oi_1 _7115_ (.B2(_0812_),
    .C1(_2771_),
    .B1(\prev_y[7] ),
    .A1(_0845_),
    .Y(_2772_),
    .A2(\prev_y[2] ));
 sg13g2_a22oi_1 _7116_ (.Y(_2773_),
    .B1(_0900_),
    .B2(net2603),
    .A2(_0889_),
    .A1(net2612));
 sg13g2_and3_1 _7117_ (.X(_2774_),
    .A(_2769_),
    .B(_2772_),
    .C(_2773_));
 sg13g2_nor3_1 _7118_ (.A(net2604),
    .B(net2605),
    .C(net2607),
    .Y(_2775_));
 sg13g2_nor3_1 _7119_ (.A(\pix_y[8] ),
    .B(net2612),
    .C(net2613),
    .Y(_2776_));
 sg13g2_nand3_1 _7120_ (.B(_2775_),
    .C(_2776_),
    .A(_0812_),
    .Y(_2777_));
 sg13g2_or4_1 _7121_ (.A(\pix_y[9] ),
    .B(net2611),
    .C(net2608),
    .D(_2777_),
    .X(_2779_));
 sg13g2_a21oi_2 _7122_ (.B1(_2779_),
    .Y(_2780_),
    .A2(_2774_),
    .A1(_2768_));
 sg13g2_o21ai_1 _7123_ (.B1(net2627),
    .Y(_2781_),
    .A1(\logo_left[0] ),
    .A2(net2190));
 sg13g2_a21oi_1 _7124_ (.A1(_0768_),
    .A2(net2190),
    .Y(_0027_),
    .B1(_2781_));
 sg13g2_nor2b_1 _7125_ (.A(net2617),
    .B_N(\logo_left[1] ),
    .Y(_2782_));
 sg13g2_nand2b_1 _7126_ (.Y(_2783_),
    .B(net2617),
    .A_N(\logo_left[1] ));
 sg13g2_nand2b_1 _7127_ (.Y(_2784_),
    .B(_2783_),
    .A_N(_2782_));
 sg13g2_xnor2_1 _7128_ (.Y(_2785_),
    .A(net106),
    .B(_2784_));
 sg13g2_o21ai_1 _7129_ (.B1(net2627),
    .Y(_2786_),
    .A1(net130),
    .A2(net2191));
 sg13g2_a21oi_1 _7130_ (.A1(net2191),
    .A2(_2785_),
    .Y(_0028_),
    .B1(_2786_));
 sg13g2_xor2_1 _7131_ (.B(\logo_left[2] ),
    .A(net2617),
    .X(_2788_));
 sg13g2_o21ai_1 _7132_ (.B1(_2783_),
    .Y(_2789_),
    .A1(\logo_left[0] ),
    .A2(_2782_));
 sg13g2_nor2_1 _7133_ (.A(_2788_),
    .B(_2789_),
    .Y(_2790_));
 sg13g2_xnor2_1 _7134_ (.Y(_2791_),
    .A(_2788_),
    .B(_2789_));
 sg13g2_o21ai_1 _7135_ (.B1(net2627),
    .Y(_2792_),
    .A1(net170),
    .A2(net2190));
 sg13g2_a21oi_1 _7136_ (.A1(net2190),
    .A2(_2791_),
    .Y(_0029_),
    .B1(_2792_));
 sg13g2_a21oi_1 _7137_ (.A1(_0669_),
    .A2(\logo_left[2] ),
    .Y(_2793_),
    .B1(_2790_));
 sg13g2_nand2_1 _7138_ (.Y(_2794_),
    .A(_0669_),
    .B(\logo_left[3] ));
 sg13g2_nor2_1 _7139_ (.A(_0669_),
    .B(net2618),
    .Y(_2795_));
 sg13g2_xor2_1 _7140_ (.B(net2618),
    .A(net2617),
    .X(_2796_));
 sg13g2_xnor2_1 _7141_ (.Y(_2798_),
    .A(_2793_),
    .B(_2796_));
 sg13g2_o21ai_1 _7142_ (.B1(net2627),
    .Y(_2799_),
    .A1(net2618),
    .A2(net2189));
 sg13g2_a21oi_1 _7143_ (.A1(net2189),
    .A2(_2798_),
    .Y(_0030_),
    .B1(_2799_));
 sg13g2_nand2_1 _7144_ (.Y(_2800_),
    .A(_0669_),
    .B(\logo_left[4] ));
 sg13g2_xor2_1 _7145_ (.B(\logo_left[4] ),
    .A(net2616),
    .X(_2801_));
 sg13g2_a21oi_1 _7146_ (.A1(_2793_),
    .A2(_2794_),
    .Y(_2802_),
    .B1(_2795_));
 sg13g2_nand2b_1 _7147_ (.Y(_2803_),
    .B(_2802_),
    .A_N(_2801_));
 sg13g2_xor2_1 _7148_ (.B(_2802_),
    .A(_2801_),
    .X(_2804_));
 sg13g2_o21ai_1 _7149_ (.B1(net2627),
    .Y(_2805_),
    .A1(net168),
    .A2(net2189));
 sg13g2_a21oi_1 _7150_ (.A1(net2189),
    .A2(_2804_),
    .Y(_0031_),
    .B1(_2805_));
 sg13g2_xor2_1 _7151_ (.B(\logo_left[5] ),
    .A(net2616),
    .X(_2807_));
 sg13g2_nand2_1 _7152_ (.Y(_2808_),
    .A(_2800_),
    .B(_2803_));
 sg13g2_o21ai_1 _7153_ (.B1(net2189),
    .Y(_2809_),
    .A1(_2807_),
    .A2(_2808_));
 sg13g2_a21oi_1 _7154_ (.A1(_2807_),
    .A2(_2808_),
    .Y(_2810_),
    .B1(_2809_));
 sg13g2_nand2_2 _7155_ (.Y(_2811_),
    .A(net2628),
    .B(net2190));
 sg13g2_o21ai_1 _7156_ (.B1(net2627),
    .Y(_2812_),
    .A1(net176),
    .A2(net2189));
 sg13g2_nor2_1 _7157_ (.A(_2810_),
    .B(_2812_),
    .Y(_0032_));
 sg13g2_o21ai_1 _7158_ (.B1(_2811_),
    .Y(_2813_),
    .A1(\logo_left[6] ),
    .A2(net2622));
 sg13g2_nor2b_1 _7159_ (.A(net2616),
    .B_N(\logo_left[6] ),
    .Y(_2814_));
 sg13g2_xnor2_1 _7160_ (.Y(_2815_),
    .A(net2616),
    .B(\logo_left[6] ));
 sg13g2_inv_1 _7161_ (.Y(_2817_),
    .A(_2815_));
 sg13g2_o21ai_1 _7162_ (.B1(_2800_),
    .Y(_2818_),
    .A1(net2616),
    .A2(_0757_));
 sg13g2_or2_1 _7163_ (.X(_2819_),
    .B(_2807_),
    .A(_2803_));
 sg13g2_nand2b_1 _7164_ (.Y(_2820_),
    .B(_2819_),
    .A_N(_2818_));
 sg13g2_and2_1 _7165_ (.A(_2815_),
    .B(_2820_),
    .X(_2821_));
 sg13g2_o21ai_1 _7166_ (.B1(net2189),
    .Y(_2822_),
    .A1(_2815_),
    .A2(_2820_));
 sg13g2_o21ai_1 _7167_ (.B1(_2813_),
    .Y(_0033_),
    .A1(_2821_),
    .A2(_2822_));
 sg13g2_o21ai_1 _7168_ (.B1(_2811_),
    .Y(_2823_),
    .A1(\logo_left[7] ),
    .A2(_0878_));
 sg13g2_nor2b_1 _7169_ (.A(net2616),
    .B_N(\logo_left[7] ),
    .Y(_2824_));
 sg13g2_xor2_1 _7170_ (.B(\logo_left[7] ),
    .A(net2616),
    .X(_2825_));
 sg13g2_a21oi_1 _7171_ (.A1(_2815_),
    .A2(_2820_),
    .Y(_2827_),
    .B1(_2814_));
 sg13g2_and2_1 _7172_ (.A(_2825_),
    .B(_2827_),
    .X(_2828_));
 sg13g2_o21ai_1 _7173_ (.B1(net2189),
    .Y(_2829_),
    .A1(_2825_),
    .A2(_2827_));
 sg13g2_o21ai_1 _7174_ (.B1(_2823_),
    .Y(_0034_),
    .A1(_2828_),
    .A2(_2829_));
 sg13g2_nor3_1 _7175_ (.A(_2817_),
    .B(_2819_),
    .C(_2825_),
    .Y(_2830_));
 sg13g2_nor4_2 _7176_ (.A(_2814_),
    .B(_2818_),
    .C(_2824_),
    .Y(_2831_),
    .D(_2830_));
 sg13g2_nand2_1 _7177_ (.Y(_2832_),
    .A(dir_x),
    .B(_2831_));
 sg13g2_o21ai_1 _7178_ (.B1(net2191),
    .Y(_2833_),
    .A1(net2616),
    .A2(_2831_));
 sg13g2_nor2b_1 _7179_ (.A(_2833_),
    .B_N(_2832_),
    .Y(_2834_));
 sg13g2_o21ai_1 _7180_ (.B1(net2628),
    .Y(_2835_),
    .A1(net147),
    .A2(_2834_));
 sg13g2_a21oi_1 _7181_ (.A1(net147),
    .A2(_2834_),
    .Y(_0035_),
    .B1(_2835_));
 sg13g2_nor2_1 _7182_ (.A(\logo_left[8] ),
    .B(_2831_),
    .Y(_2837_));
 sg13g2_a21oi_1 _7183_ (.A1(_0669_),
    .A2(\logo_left[8] ),
    .Y(_2838_),
    .B1(_2837_));
 sg13g2_and3_1 _7184_ (.X(_2839_),
    .A(net2191),
    .B(_2832_),
    .C(_2838_));
 sg13g2_o21ai_1 _7185_ (.B1(net2627),
    .Y(_2840_),
    .A1(net156),
    .A2(_2839_));
 sg13g2_a21oi_1 _7186_ (.A1(net156),
    .A2(_2839_),
    .Y(_0036_),
    .B1(_2840_));
 sg13g2_o21ai_1 _7187_ (.B1(net2625),
    .Y(_2841_),
    .A1(\logo_top[0] ),
    .A2(net2187));
 sg13g2_a21oi_1 _7188_ (.A1(_0746_),
    .A2(net2187),
    .Y(_0037_),
    .B1(_2841_));
 sg13g2_xnor2_1 _7189_ (.Y(_2842_),
    .A(net2615),
    .B(\logo_top[1] ));
 sg13g2_xnor2_1 _7190_ (.Y(_2843_),
    .A(_0746_),
    .B(_2842_));
 sg13g2_o21ai_1 _7191_ (.B1(net2625),
    .Y(_2845_),
    .A1(net131),
    .A2(net2187));
 sg13g2_a21oi_1 _7192_ (.A1(net2187),
    .A2(_2843_),
    .Y(_0038_),
    .B1(_2845_));
 sg13g2_xor2_1 _7193_ (.B(\logo_top[2] ),
    .A(net2615),
    .X(_2846_));
 sg13g2_a21o_1 _7194_ (.A2(\logo_top[1] ),
    .A1(net2602),
    .B1(\logo_top[0] ),
    .X(_2847_));
 sg13g2_o21ai_1 _7195_ (.B1(_2847_),
    .Y(_2848_),
    .A1(net2602),
    .A2(\logo_top[1] ));
 sg13g2_nor2_1 _7196_ (.A(_2846_),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_xnor2_1 _7197_ (.Y(_2850_),
    .A(_2846_),
    .B(_2848_));
 sg13g2_o21ai_1 _7198_ (.B1(net1),
    .Y(_2851_),
    .A1(net165),
    .A2(net2187));
 sg13g2_a21oi_1 _7199_ (.A1(net2187),
    .A2(_2850_),
    .Y(_0039_),
    .B1(_2851_));
 sg13g2_a21oi_1 _7200_ (.A1(net2602),
    .A2(\logo_top[2] ),
    .Y(_2852_),
    .B1(_2849_));
 sg13g2_nand2_1 _7201_ (.Y(_2854_),
    .A(net2602),
    .B(\logo_top[3] ));
 sg13g2_nor2_1 _7202_ (.A(net2602),
    .B(\logo_top[3] ),
    .Y(_2855_));
 sg13g2_xor2_1 _7203_ (.B(\logo_top[3] ),
    .A(net2615),
    .X(_2856_));
 sg13g2_xnor2_1 _7204_ (.Y(_2857_),
    .A(_2852_),
    .B(_2856_));
 sg13g2_o21ai_1 _7205_ (.B1(net2626),
    .Y(_2858_),
    .A1(net175),
    .A2(net2187));
 sg13g2_a21oi_1 _7206_ (.A1(net2187),
    .A2(_2857_),
    .Y(_0040_),
    .B1(_2858_));
 sg13g2_o21ai_1 _7207_ (.B1(_2811_),
    .Y(_2859_),
    .A1(net177),
    .A2(net2622));
 sg13g2_nand2_1 _7208_ (.Y(_2860_),
    .A(_0658_),
    .B(\logo_top[4] ));
 sg13g2_xnor2_1 _7209_ (.Y(_2861_),
    .A(net2614),
    .B(\logo_top[4] ));
 sg13g2_a21oi_1 _7210_ (.A1(_2852_),
    .A2(_2854_),
    .Y(_2862_),
    .B1(_2855_));
 sg13g2_nor2_1 _7211_ (.A(_2861_),
    .B(_2862_),
    .Y(_2864_));
 sg13g2_nand2_1 _7212_ (.Y(_2865_),
    .A(_2861_),
    .B(_2862_));
 sg13g2_nand2_1 _7213_ (.Y(_2866_),
    .A(_2780_),
    .B(_2865_));
 sg13g2_o21ai_1 _7214_ (.B1(_2859_),
    .Y(_0041_),
    .A1(_2864_),
    .A2(_2866_));
 sg13g2_xor2_1 _7215_ (.B(\logo_top[5] ),
    .A(net2615),
    .X(_2867_));
 sg13g2_nand3_1 _7216_ (.B(_2865_),
    .C(_2867_),
    .A(_2860_),
    .Y(_2868_));
 sg13g2_a21oi_1 _7217_ (.A1(_2860_),
    .A2(_2865_),
    .Y(_2869_),
    .B1(_2867_));
 sg13g2_nand2_1 _7218_ (.Y(_2870_),
    .A(net2188),
    .B(_2868_));
 sg13g2_o21ai_1 _7219_ (.B1(_2811_),
    .Y(_2871_),
    .A1(net174),
    .A2(net2622));
 sg13g2_o21ai_1 _7220_ (.B1(_2871_),
    .Y(_0042_),
    .A1(_2869_),
    .A2(_2870_));
 sg13g2_nor2_1 _7221_ (.A(net2615),
    .B(_0691_),
    .Y(_2873_));
 sg13g2_xor2_1 _7222_ (.B(\logo_top[6] ),
    .A(net2614),
    .X(_2874_));
 sg13g2_nor2_1 _7223_ (.A(_2865_),
    .B(_2867_),
    .Y(_2875_));
 sg13g2_a21oi_1 _7224_ (.A1(_0702_),
    .A2(_0713_),
    .Y(_2876_),
    .B1(net2614));
 sg13g2_nor2_1 _7225_ (.A(_2875_),
    .B(_2876_),
    .Y(_2877_));
 sg13g2_nand2_1 _7226_ (.Y(_2878_),
    .A(_2874_),
    .B(_2877_));
 sg13g2_nor2_1 _7227_ (.A(_2874_),
    .B(_2877_),
    .Y(_2879_));
 sg13g2_nand2_1 _7228_ (.Y(_2880_),
    .A(net2188),
    .B(_2878_));
 sg13g2_o21ai_1 _7229_ (.B1(_2811_),
    .Y(_2881_),
    .A1(net171),
    .A2(net2622));
 sg13g2_o21ai_1 _7230_ (.B1(_2881_),
    .Y(_0043_),
    .A1(_2879_),
    .A2(_2880_));
 sg13g2_o21ai_1 _7231_ (.B1(net2629),
    .Y(_2883_),
    .A1(net166),
    .A2(net2188));
 sg13g2_xnor2_1 _7232_ (.Y(_2884_),
    .A(net2614),
    .B(\logo_top[7] ));
 sg13g2_nor2_1 _7233_ (.A(_2873_),
    .B(_2879_),
    .Y(_2885_));
 sg13g2_o21ai_1 _7234_ (.B1(net2188),
    .Y(_2886_),
    .A1(_2884_),
    .A2(_2885_));
 sg13g2_a21oi_1 _7235_ (.A1(_2884_),
    .A2(_2885_),
    .Y(_2887_),
    .B1(_2886_));
 sg13g2_nor2_1 _7236_ (.A(_2883_),
    .B(_2887_),
    .Y(_0044_));
 sg13g2_nor2b_1 _7237_ (.A(_2874_),
    .B_N(_2884_),
    .Y(_2888_));
 sg13g2_or2_1 _7238_ (.X(_2889_),
    .B(_2876_),
    .A(_2873_));
 sg13g2_a221oi_1 _7239_ (.B2(_2888_),
    .C1(_2889_),
    .B1(_2875_),
    .A1(_0658_),
    .Y(_2890_),
    .A2(\logo_top[7] ));
 sg13g2_o21ai_1 _7240_ (.B1(net2188),
    .Y(_2891_),
    .A1(net2614),
    .A2(_2890_));
 sg13g2_a21oi_1 _7241_ (.A1(net2614),
    .A2(_2890_),
    .Y(_2893_),
    .B1(_2891_));
 sg13g2_o21ai_1 _7242_ (.B1(net2626),
    .Y(_2894_),
    .A1(net153),
    .A2(_2893_));
 sg13g2_nand2_1 _7243_ (.Y(_2895_),
    .A(net2602),
    .B(\logo_top[8] ));
 sg13g2_a21oi_1 _7244_ (.A1(net153),
    .A2(_2893_),
    .Y(_0045_),
    .B1(_2894_));
 sg13g2_nor2_1 _7245_ (.A(\logo_top[8] ),
    .B(_2890_),
    .Y(_2896_));
 sg13g2_a21oi_1 _7246_ (.A1(net2614),
    .A2(_2890_),
    .Y(_2897_),
    .B1(_2896_));
 sg13g2_and3_1 _7247_ (.X(_2898_),
    .A(net2188),
    .B(_2895_),
    .C(_2897_));
 sg13g2_o21ai_1 _7248_ (.B1(net2626),
    .Y(_2899_),
    .A1(net127),
    .A2(_2898_));
 sg13g2_a21oi_1 _7249_ (.A1(net127),
    .A2(_2898_),
    .Y(_0046_),
    .B1(_2899_));
 sg13g2_nand3_1 _7250_ (.B(\logo_left[1] ),
    .C(\logo_left[0] ),
    .A(\logo_left[2] ),
    .Y(_2900_));
 sg13g2_nand4_1 _7251_ (.B(\logo_left[5] ),
    .C(\logo_left[4] ),
    .A(\logo_left[6] ),
    .Y(_2902_),
    .D(net2618));
 sg13g2_nor2_1 _7252_ (.A(_2900_),
    .B(_2902_),
    .Y(_2903_));
 sg13g2_nor2_1 _7253_ (.A(\logo_left[8] ),
    .B(_0004_),
    .Y(_2904_));
 sg13g2_and4_1 _7254_ (.A(\logo_left[9] ),
    .B(\logo_left[7] ),
    .C(_2903_),
    .D(_2904_),
    .X(_2905_));
 sg13g2_nor2b_1 _7255_ (.A(\logo_left[9] ),
    .B_N(_0004_),
    .Y(_2906_));
 sg13g2_nor3_1 _7256_ (.A(\logo_left[9] ),
    .B(\logo_left[7] ),
    .C(_2903_),
    .Y(_2907_));
 sg13g2_nor4_1 _7257_ (.A(_0669_),
    .B(_2905_),
    .C(_2906_),
    .D(_2907_),
    .Y(_2908_));
 sg13g2_nor4_1 _7258_ (.A(net2617),
    .B(\logo_left[9] ),
    .C(\logo_left[7] ),
    .D(\logo_left[6] ),
    .Y(_2909_));
 sg13g2_or2_1 _7259_ (.X(_2910_),
    .B(\logo_left[2] ),
    .A(net2618));
 sg13g2_nand4_1 _7260_ (.B(_0003_),
    .C(_0004_),
    .A(\logo_left[0] ),
    .Y(_2911_),
    .D(_2909_));
 sg13g2_nor4_1 _7261_ (.A(\logo_left[5] ),
    .B(\logo_left[1] ),
    .C(_2910_),
    .D(_2911_),
    .Y(_2913_));
 sg13g2_o21ai_1 _7262_ (.B1(net2190),
    .Y(_2914_),
    .A1(_2908_),
    .A2(_2913_));
 sg13g2_nor2_1 _7263_ (.A(_0669_),
    .B(net102),
    .Y(_2915_));
 sg13g2_a21oi_1 _7264_ (.A1(net2617),
    .A2(_2914_),
    .Y(_2916_),
    .B1(_0878_));
 sg13g2_o21ai_1 _7265_ (.B1(_2916_),
    .Y(_0047_),
    .A1(_2914_),
    .A2(_2915_));
 sg13g2_nor4_1 _7266_ (.A(net2614),
    .B(\logo_top[7] ),
    .C(\logo_top[6] ),
    .D(\logo_top[3] ),
    .Y(_2917_));
 sg13g2_nand4_1 _7267_ (.B(_0006_),
    .C(_0007_),
    .A(_0724_),
    .Y(_2918_),
    .D(_2917_));
 sg13g2_nand2b_1 _7268_ (.Y(_2919_),
    .B(_2918_),
    .A_N(\logo_top[1] ));
 sg13g2_nor3_1 _7269_ (.A(\logo_top[9] ),
    .B(\logo_top[5] ),
    .C(_0735_),
    .Y(_2920_));
 sg13g2_nand3_1 _7270_ (.B(\logo_top[3] ),
    .C(\logo_top[2] ),
    .A(\logo_top[4] ),
    .Y(_2921_));
 sg13g2_or4_1 _7271_ (.A(_0658_),
    .B(\logo_top[8] ),
    .C(_0680_),
    .D(_0691_),
    .X(_2923_));
 sg13g2_o21ai_1 _7272_ (.B1(\logo_top[1] ),
    .Y(_2924_),
    .A1(_2921_),
    .A2(_2923_));
 sg13g2_nand4_1 _7273_ (.B(_2919_),
    .C(_2920_),
    .A(net2188),
    .Y(_2925_),
    .D(_2924_));
 sg13g2_and2_1 _7274_ (.A(net2602),
    .B(_2925_),
    .X(_2926_));
 sg13g2_nor3_1 _7275_ (.A(net2602),
    .B(net116),
    .C(_2925_),
    .Y(_2927_));
 sg13g2_nor3_1 _7276_ (.A(net2622),
    .B(_2926_),
    .C(_2927_),
    .Y(_0048_));
 sg13g2_nand2_2 _7277_ (.Y(_2928_),
    .A(_2914_),
    .B(_2925_));
 sg13g2_o21ai_1 _7278_ (.B1(net2626),
    .Y(_2929_),
    .A1(\color_index[0] ),
    .A2(_2928_));
 sg13g2_a21oi_1 _7279_ (.A1(_0647_),
    .A2(_2928_),
    .Y(_0049_),
    .B1(_2929_));
 sg13g2_and2_1 _7280_ (.A(\color_index[0] ),
    .B(_2928_),
    .X(_2930_));
 sg13g2_nand2_1 _7281_ (.Y(_2932_),
    .A(net143),
    .B(_2930_));
 sg13g2_o21ai_1 _7282_ (.B1(net2626),
    .Y(_2933_),
    .A1(net143),
    .A2(_2930_));
 sg13g2_nor2b_1 _7283_ (.A(net144),
    .B_N(_2932_),
    .Y(_0050_));
 sg13g2_o21ai_1 _7284_ (.B1(net2626),
    .Y(_2934_),
    .A1(_0636_),
    .A2(_2932_));
 sg13g2_a21oi_1 _7285_ (.A1(_0636_),
    .A2(_2932_),
    .Y(_0051_),
    .B1(_2934_));
 sg13g2_mux2_1 _7286_ (.A0(net125),
    .A1(net2613),
    .S(net2623),
    .X(_0052_));
 sg13g2_nand2_1 _7287_ (.Y(_2935_),
    .A(net2612),
    .B(net2623));
 sg13g2_o21ai_1 _7288_ (.B1(_2935_),
    .Y(_0053_),
    .A1(net2624),
    .A2(_0889_));
 sg13g2_mux2_1 _7289_ (.A0(net121),
    .A1(net2610),
    .S(net2623),
    .X(_0054_));
 sg13g2_mux2_1 _7290_ (.A0(net115),
    .A1(net2608),
    .S(net2625),
    .X(_0055_));
 sg13g2_nor2_1 _7291_ (.A(net2623),
    .B(net113),
    .Y(_2937_));
 sg13g2_a21oi_1 _7292_ (.A1(_0834_),
    .A2(net2623),
    .Y(_0056_),
    .B1(_2937_));
 sg13g2_mux2_1 _7293_ (.A0(net119),
    .A1(net2605),
    .S(net2625),
    .X(_0057_));
 sg13g2_nor2_1 _7294_ (.A(net2623),
    .B(net108),
    .Y(_2938_));
 sg13g2_a21oi_1 _7295_ (.A1(_0823_),
    .A2(net2623),
    .Y(_0058_),
    .B1(_2938_));
 sg13g2_nor2_1 _7296_ (.A(net2624),
    .B(net122),
    .Y(_2939_));
 sg13g2_a21oi_1 _7297_ (.A1(_0812_),
    .A2(net2624),
    .Y(_0059_),
    .B1(_2939_));
 sg13g2_nor2_1 _7298_ (.A(net2624),
    .B(net118),
    .Y(_2940_));
 sg13g2_a21oi_1 _7299_ (.A1(_0790_),
    .A2(net2623),
    .Y(_0060_),
    .B1(_2940_));
 sg13g2_a21oi_1 _7300_ (.A1(net2622),
    .A2(_0922_),
    .Y(_0061_),
    .B1(_2721_));
 sg13g2_nor2_1 _7301_ (.A(net111),
    .B(_2811_),
    .Y(_2942_));
 sg13g2_nor3_2 _7302_ (.A(\frame_divider[0] ),
    .B(net111),
    .C(_2811_),
    .Y(_2943_));
 sg13g2_mux2_1 _7303_ (.A0(\frame_counter[0] ),
    .A1(net100),
    .S(_2943_),
    .X(_0062_));
 sg13g2_nand3_1 _7304_ (.B(\frame_counter[1] ),
    .C(_2943_),
    .A(net179),
    .Y(_2944_));
 sg13g2_a21o_1 _7305_ (.A2(_2943_),
    .A1(net179),
    .B1(\frame_counter[1] ),
    .X(_2945_));
 sg13g2_and2_1 _7306_ (.A(_2944_),
    .B(net180),
    .X(_0063_));
 sg13g2_nand4_1 _7307_ (.B(\frame_counter[2] ),
    .C(\frame_counter[1] ),
    .A(\frame_counter[0] ),
    .Y(_2946_),
    .D(_2943_));
 sg13g2_xnor2_1 _7308_ (.Y(_0064_),
    .A(net151),
    .B(_2944_));
 sg13g2_nor2_1 _7309_ (.A(_0955_),
    .B(_2946_),
    .Y(_2947_));
 sg13g2_xnor2_1 _7310_ (.Y(_0065_),
    .A(net149),
    .B(_2946_));
 sg13g2_and2_1 _7311_ (.A(\frame_counter[4] ),
    .B(_2947_),
    .X(_2949_));
 sg13g2_xor2_1 _7312_ (.B(_2947_),
    .A(net139),
    .X(_0066_));
 sg13g2_xor2_1 _7313_ (.B(_2949_),
    .A(net154),
    .X(_0067_));
 sg13g2_nand3_1 _7314_ (.B(net178),
    .C(_2949_),
    .A(net154),
    .Y(_2950_));
 sg13g2_a21o_1 _7315_ (.A2(_2949_),
    .A1(net154),
    .B1(net178),
    .X(_2951_));
 sg13g2_and2_1 _7316_ (.A(_2950_),
    .B(_2951_),
    .X(_0068_));
 sg13g2_xnor2_1 _7317_ (.Y(_0069_),
    .A(net128),
    .B(_2950_));
 sg13g2_mux2_1 _7318_ (.A0(net98),
    .A1(\frame_divider[0] ),
    .S(_2811_),
    .X(_0070_));
 sg13g2_nand3_1 _7319_ (.B(net2627),
    .C(net2190),
    .A(\frame_divider[0] ),
    .Y(_2952_));
 sg13g2_a22oi_1 _7320_ (.Y(_2953_),
    .B1(_2952_),
    .B2(net111),
    .A2(_2942_),
    .A1(\frame_divider[0] ));
 sg13g2_inv_1 _7321_ (.Y(_0071_),
    .A(net112));
 sg13g2_and2_1 _7322_ (.A(net183),
    .B(_2725_),
    .X(_2955_));
 sg13g2_a21oi_1 _7323_ (.A1(_2677_),
    .A2(_2955_),
    .Y(_0072_),
    .B1(_2723_));
 sg13g2_xnor2_1 _7324_ (.Y(_2956_),
    .A(net2604),
    .B(\frame_counter[6] ));
 sg13g2_a21oi_1 _7325_ (.A1(_2678_),
    .A2(_2692_),
    .Y(_2957_),
    .B1(_2956_));
 sg13g2_nand3_1 _7326_ (.B(_2692_),
    .C(_2956_),
    .A(_2678_),
    .Y(_2958_));
 sg13g2_nor2b_1 _7327_ (.A(_2957_),
    .B_N(_2958_),
    .Y(_2959_));
 sg13g2_xnor2_1 _7328_ (.Y(_2960_),
    .A(net2619),
    .B(_2959_));
 sg13g2_xnor2_1 _7329_ (.Y(_2961_),
    .A(_2718_),
    .B(_2960_));
 sg13g2_nor2_1 _7330_ (.A(_2677_),
    .B(_2961_),
    .Y(_2962_));
 sg13g2_and4_1 _7331_ (.A(net143),
    .B(net3),
    .C(_2677_),
    .D(_2733_),
    .X(_2964_));
 sg13g2_nor3_1 _7332_ (.A(_2723_),
    .B(_2962_),
    .C(_2964_),
    .Y(_0073_));
 sg13g2_xor2_1 _7333_ (.B(_2960_),
    .A(_2711_),
    .X(_2965_));
 sg13g2_nand2_1 _7334_ (.Y(_2966_),
    .A(_0636_),
    .B(\color_index[1] ));
 sg13g2_nand3b_1 _7335_ (.B(net3),
    .C(_2966_),
    .Y(_2967_),
    .A_N(\color_index[0] ));
 sg13g2_nand2_1 _7336_ (.Y(_2968_),
    .A(net143),
    .B(_2955_));
 sg13g2_nand2_1 _7337_ (.Y(_2969_),
    .A(_2967_),
    .B(_2968_));
 sg13g2_mux2_1 _7338_ (.A0(_2965_),
    .A1(_2969_),
    .S(_2677_),
    .X(_2970_));
 sg13g2_nor2_1 _7339_ (.A(_2723_),
    .B(_2970_),
    .Y(_0074_));
 sg13g2_and3_1 _7340_ (.X(_2971_),
    .A(net3),
    .B(_2735_),
    .C(_2966_));
 sg13g2_a21oi_1 _7341_ (.A1(net2604),
    .A2(\frame_counter[6] ),
    .Y(_2973_),
    .B1(_2957_));
 sg13g2_xnor2_1 _7342_ (.Y(_2974_),
    .A(\pix_x[8] ),
    .B(\pix_y[7] ));
 sg13g2_xnor2_1 _7343_ (.Y(_2975_),
    .A(\frame_counter[7] ),
    .B(_2974_));
 sg13g2_xnor2_1 _7344_ (.Y(_2976_),
    .A(_2973_),
    .B(_2975_));
 sg13g2_xnor2_1 _7345_ (.Y(_2977_),
    .A(_2711_),
    .B(_2976_));
 sg13g2_mux2_1 _7346_ (.A0(_2977_),
    .A1(_2971_),
    .S(_2677_),
    .X(_2978_));
 sg13g2_nor2_1 _7347_ (.A(_2723_),
    .B(_2978_),
    .Y(_0075_));
 sg13g2_nand3_1 _7348_ (.B(net2610),
    .C(net2609),
    .A(\pix_y[9] ),
    .Y(_2979_));
 sg13g2_o21ai_1 _7349_ (.B1(net2625),
    .Y(_2980_),
    .A1(_2777_),
    .A2(_2979_));
 sg13g2_inv_1 _7350_ (.Y(_2981_),
    .A(_2980_));
 sg13g2_nor2_2 _7351_ (.A(_2742_),
    .B(_2980_),
    .Y(_2983_));
 sg13g2_a22oi_1 _7352_ (.Y(_2984_),
    .B1(_2983_),
    .B2(net94),
    .A2(_2743_),
    .A1(net2613));
 sg13g2_inv_1 _7353_ (.Y(_0076_),
    .A(net95));
 sg13g2_and2_1 _7354_ (.A(net2612),
    .B(net2613),
    .X(_2985_));
 sg13g2_xor2_1 _7355_ (.B(net2613),
    .A(net2612),
    .X(_2986_));
 sg13g2_a22oi_1 _7356_ (.Y(_2987_),
    .B1(_2983_),
    .B2(_2986_),
    .A2(_2743_),
    .A1(net2612));
 sg13g2_inv_1 _7357_ (.Y(_0077_),
    .A(_2987_));
 sg13g2_and2_1 _7358_ (.A(net2610),
    .B(_2985_),
    .X(_2988_));
 sg13g2_nor2_1 _7359_ (.A(_2980_),
    .B(_2988_),
    .Y(_2989_));
 sg13g2_nor2_1 _7360_ (.A(_2743_),
    .B(_2989_),
    .Y(_2990_));
 sg13g2_a21oi_1 _7361_ (.A1(net2304),
    .A2(_2985_),
    .Y(_2992_),
    .B1(net2610));
 sg13g2_nor2_1 _7362_ (.A(_2990_),
    .B(_2992_),
    .Y(_0078_));
 sg13g2_o21ai_1 _7363_ (.B1(net2608),
    .Y(_2993_),
    .A1(_2743_),
    .A2(_2989_));
 sg13g2_nand2_1 _7364_ (.Y(_2994_),
    .A(_2983_),
    .B(_2988_));
 sg13g2_o21ai_1 _7365_ (.B1(_2993_),
    .Y(_0079_),
    .A1(net2608),
    .A2(_2994_));
 sg13g2_and3_1 _7366_ (.X(_2995_),
    .A(net2607),
    .B(net2608),
    .C(_2988_));
 sg13g2_o21ai_1 _7367_ (.B1(net2304),
    .Y(_2996_),
    .A1(_2980_),
    .A2(_2995_));
 sg13g2_nand4_1 _7368_ (.B(net2608),
    .C(net2304),
    .A(net2610),
    .Y(_2997_),
    .D(_2985_));
 sg13g2_nand2_1 _7369_ (.Y(_2998_),
    .A(_0834_),
    .B(_2997_));
 sg13g2_and2_1 _7370_ (.A(_2996_),
    .B(_2998_),
    .X(_0080_));
 sg13g2_nand2_1 _7371_ (.Y(_3000_),
    .A(net2605),
    .B(_2996_));
 sg13g2_nand2_1 _7372_ (.Y(_3001_),
    .A(_2983_),
    .B(_2995_));
 sg13g2_o21ai_1 _7373_ (.B1(_3000_),
    .Y(_0081_),
    .A1(net2605),
    .A2(_3001_));
 sg13g2_and2_1 _7374_ (.A(net2605),
    .B(_2995_),
    .X(_3002_));
 sg13g2_a21oi_1 _7375_ (.A1(net2603),
    .A2(_3002_),
    .Y(_3003_),
    .B1(_2980_));
 sg13g2_nor2_1 _7376_ (.A(_2743_),
    .B(_3003_),
    .Y(_3004_));
 sg13g2_a21oi_1 _7377_ (.A1(net2304),
    .A2(_3002_),
    .Y(_3005_),
    .B1(net2603));
 sg13g2_nor2_1 _7378_ (.A(_3004_),
    .B(_3005_),
    .Y(_0082_));
 sg13g2_nand4_1 _7379_ (.B(net2603),
    .C(_2983_),
    .A(_0812_),
    .Y(_3006_),
    .D(_3002_));
 sg13g2_o21ai_1 _7380_ (.B1(_3006_),
    .Y(_0083_),
    .A1(_0812_),
    .A2(_3004_));
 sg13g2_a21oi_1 _7381_ (.A1(_2720_),
    .A2(_2981_),
    .Y(_3008_),
    .B1(_2996_));
 sg13g2_nand4_1 _7382_ (.B(net2603),
    .C(net2304),
    .A(net173),
    .Y(_3009_),
    .D(_3002_));
 sg13g2_a21oi_1 _7383_ (.A1(_0790_),
    .A2(_3009_),
    .Y(_0084_),
    .B1(_3008_));
 sg13g2_or3_1 _7384_ (.A(_0966_),
    .B(_2980_),
    .C(_3009_),
    .X(_3010_));
 sg13g2_o21ai_1 _7385_ (.B1(_3010_),
    .Y(_0085_),
    .A1(_0801_),
    .A2(_3008_));
 sg13g2_dfrbp_1 _7386_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(_0015_),
    .Q_N(_3690_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7387_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net74),
    .D(_0016_),
    .Q_N(_3689_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7388_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net73),
    .D(_0017_),
    .Q_N(_0014_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _7389_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net72),
    .D(_0018_),
    .Q_N(_3688_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _7390_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net71),
    .D(_0019_),
    .Q_N(_3687_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _7391_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net70),
    .D(_0020_),
    .Q_N(_3686_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _7392_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net69),
    .D(_0021_),
    .Q_N(_3685_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _7393_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net68),
    .D(_0022_),
    .Q_N(_3684_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _7394_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net67),
    .D(_0023_),
    .Q_N(_3683_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _7395_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net66),
    .D(_0024_),
    .Q_N(_3682_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _7396_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net65),
    .D(_0025_),
    .Q_N(_3681_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _7397_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net64),
    .D(_0026_),
    .Q_N(_3680_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _7398_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net63),
    .D(net107),
    .Q_N(_0013_),
    .Q(\logo_left[0] ));
 sg13g2_dfrbp_1 _7399_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net61),
    .D(_0028_),
    .Q_N(_3679_),
    .Q(\logo_left[1] ));
 sg13g2_dfrbp_1 _7400_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net59),
    .D(_0029_),
    .Q_N(_3678_),
    .Q(\logo_left[2] ));
 sg13g2_dfrbp_1 _7401_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net57),
    .D(_0030_),
    .Q_N(_3677_),
    .Q(\logo_left[3] ));
 sg13g2_dfrbp_1 _7402_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net55),
    .D(net169),
    .Q_N(_0003_),
    .Q(\logo_left[4] ));
 sg13g2_dfrbp_1 _7403_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net53),
    .D(_0032_),
    .Q_N(_3676_),
    .Q(\logo_left[5] ));
 sg13g2_dfrbp_1 _7404_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net51),
    .D(_0033_),
    .Q_N(_3675_),
    .Q(\logo_left[6] ));
 sg13g2_dfrbp_1 _7405_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net49),
    .D(_0034_),
    .Q_N(_3674_),
    .Q(\logo_left[7] ));
 sg13g2_dfrbp_1 _7406_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net47),
    .D(net148),
    .Q_N(_0004_),
    .Q(\logo_left[8] ));
 sg13g2_dfrbp_1 _7407_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net45),
    .D(net157),
    .Q_N(_3673_),
    .Q(\logo_left[9] ));
 sg13g2_dfrbp_1 _7408_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net43),
    .D(net105),
    .Q_N(_0012_),
    .Q(\logo_top[0] ));
 sg13g2_dfrbp_1 _7409_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net41),
    .D(_0038_),
    .Q_N(_3672_),
    .Q(\logo_top[1] ));
 sg13g2_dfrbp_1 _7410_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net39),
    .D(_0039_),
    .Q_N(_3671_),
    .Q(\logo_top[2] ));
 sg13g2_dfrbp_1 _7411_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net37),
    .D(_0040_),
    .Q_N(_3670_),
    .Q(\logo_top[3] ));
 sg13g2_dfrbp_1 _7412_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net35),
    .D(_0041_),
    .Q_N(_0006_),
    .Q(\logo_top[4] ));
 sg13g2_dfrbp_1 _7413_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net33),
    .D(_0042_),
    .Q_N(_3669_),
    .Q(\logo_top[5] ));
 sg13g2_dfrbp_1 _7414_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net31),
    .D(_0043_),
    .Q_N(_3668_),
    .Q(\logo_top[6] ));
 sg13g2_dfrbp_1 _7415_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net29),
    .D(net167),
    .Q_N(_3667_),
    .Q(\logo_top[7] ));
 sg13g2_dfrbp_1 _7416_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net27),
    .D(_0045_),
    .Q_N(_0007_),
    .Q(\logo_top[8] ));
 sg13g2_dfrbp_1 _7417_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net25),
    .D(_0046_),
    .Q_N(_3666_),
    .Q(\logo_top[9] ));
 sg13g2_dfrbp_1 _7418_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net23),
    .D(net103),
    .Q_N(_0002_),
    .Q(dir_x));
 sg13g2_dfrbp_1 _7419_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net21),
    .D(net117),
    .Q_N(_0005_),
    .Q(dir_y));
 sg13g2_dfrbp_1 _7420_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net91),
    .D(net97),
    .Q_N(_0011_),
    .Q(\color_index[0] ));
 sg13g2_dfrbp_1 _7421_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net89),
    .D(_0050_),
    .Q_N(_3665_),
    .Q(\color_index[1] ));
 sg13g2_dfrbp_1 _7422_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net87),
    .D(net142),
    .Q_N(_3664_),
    .Q(\color_index[2] ));
 sg13g2_dfrbp_1 _7423_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net85),
    .D(net126),
    .Q_N(_3663_),
    .Q(\prev_y[0] ));
 sg13g2_dfrbp_1 _7424_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net84),
    .D(net124),
    .Q_N(_3662_),
    .Q(\prev_y[1] ));
 sg13g2_dfrbp_1 _7425_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net83),
    .D(_0054_),
    .Q_N(_3661_),
    .Q(\prev_y[2] ));
 sg13g2_dfrbp_1 _7426_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net82),
    .D(_0055_),
    .Q_N(_3660_),
    .Q(\prev_y[3] ));
 sg13g2_dfrbp_1 _7427_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(net114),
    .Q_N(_3659_),
    .Q(\prev_y[4] ));
 sg13g2_dfrbp_1 _7428_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net79),
    .D(net120),
    .Q_N(_3658_),
    .Q(\prev_y[5] ));
 sg13g2_dfrbp_1 _7429_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net78),
    .D(_0058_),
    .Q_N(_3657_),
    .Q(\prev_y[6] ));
 sg13g2_dfrbp_1 _7430_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net77),
    .D(_0059_),
    .Q_N(_3656_),
    .Q(\prev_y[7] ));
 sg13g2_dfrbp_1 _7431_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net76),
    .D(_0060_),
    .Q_N(_3655_),
    .Q(\prev_y[8] ));
 sg13g2_dfrbp_1 _7432_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net75),
    .D(net110),
    .Q_N(_3654_),
    .Q(\prev_y[9] ));
 sg13g2_dfrbp_1 _7433_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net62),
    .D(net101),
    .Q_N(_0010_),
    .Q(\frame_counter[0] ));
 sg13g2_dfrbp_1 _7434_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net60),
    .D(net181),
    .Q_N(_3653_),
    .Q(\frame_counter[1] ));
 sg13g2_dfrbp_1 _7435_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net58),
    .D(net152),
    .Q_N(_3652_),
    .Q(\frame_counter[2] ));
 sg13g2_dfrbp_1 _7436_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net56),
    .D(net150),
    .Q_N(_3651_),
    .Q(\frame_counter[3] ));
 sg13g2_dfrbp_1 _7437_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net54),
    .D(net140),
    .Q_N(_3650_),
    .Q(\frame_counter[4] ));
 sg13g2_dfrbp_1 _7438_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net52),
    .D(net155),
    .Q_N(_3649_),
    .Q(\frame_counter[5] ));
 sg13g2_dfrbp_1 _7439_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net50),
    .D(_0068_),
    .Q_N(_3648_),
    .Q(\frame_counter[6] ));
 sg13g2_dfrbp_1 _7440_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net48),
    .D(net129),
    .Q_N(_3647_),
    .Q(\frame_counter[7] ));
 sg13g2_dfrbp_1 _7441_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net46),
    .D(net99),
    .Q_N(_0009_),
    .Q(\frame_divider[0] ));
 sg13g2_dfrbp_1 _7442_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net44),
    .D(_0071_),
    .Q_N(_3646_),
    .Q(\frame_divider[1] ));
 sg13g2_dfrbp_1 _7443_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net42),
    .D(_0072_),
    .Q_N(_3645_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7444_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(_0073_),
    .Q_N(_3644_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7445_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net38),
    .D(_0074_),
    .Q_N(_3643_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7446_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net92),
    .D(_0075_),
    .Q_N(_3691_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7447_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net36),
    .D(net138),
    .Q_N(_3642_),
    .Q(hsync));
 sg13g2_dfrbp_1 _7448_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net34),
    .D(_0076_),
    .Q_N(_0008_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _7449_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net30),
    .D(_0077_),
    .Q_N(_3641_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _7450_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net26),
    .D(_0078_),
    .Q_N(_3640_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _7451_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net22),
    .D(_0079_),
    .Q_N(_3639_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _7452_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0080_),
    .Q_N(_3638_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _7453_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net86),
    .D(_0081_),
    .Q_N(_3637_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _7454_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net28),
    .D(_0082_),
    .Q_N(_3636_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _7455_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net20),
    .D(_0083_),
    .Q_N(_3635_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _7456_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net32),
    .D(_0084_),
    .Q_N(_3634_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _7457_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net24),
    .D(_0085_),
    .Q_N(_3692_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _7458_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net88),
    .D(_0001_),
    .Q_N(_3633_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_tiehi _7419__21 (.L_HI(net21));
 sg13g2_tiehi _7451__22 (.L_HI(net22));
 sg13g2_tiehi _7418__23 (.L_HI(net23));
 sg13g2_tiehi _7457__24 (.L_HI(net24));
 sg13g2_tiehi _7417__25 (.L_HI(net25));
 sg13g2_tiehi _7450__26 (.L_HI(net26));
 sg13g2_tiehi _7416__27 (.L_HI(net27));
 sg13g2_tiehi _7454__28 (.L_HI(net28));
 sg13g2_tiehi _7415__29 (.L_HI(net29));
 sg13g2_tiehi _7449__30 (.L_HI(net30));
 sg13g2_tiehi _7414__31 (.L_HI(net31));
 sg13g2_tiehi _7456__32 (.L_HI(net32));
 sg13g2_tiehi _7413__33 (.L_HI(net33));
 sg13g2_tiehi _7448__34 (.L_HI(net34));
 sg13g2_tiehi _7412__35 (.L_HI(net35));
 sg13g2_tiehi _7447__36 (.L_HI(net36));
 sg13g2_tiehi _7411__37 (.L_HI(net37));
 sg13g2_tiehi _7445__38 (.L_HI(net38));
 sg13g2_tiehi _7410__39 (.L_HI(net39));
 sg13g2_tiehi _7444__40 (.L_HI(net40));
 sg13g2_tiehi _7409__41 (.L_HI(net41));
 sg13g2_tiehi _7443__42 (.L_HI(net42));
 sg13g2_tiehi _7408__43 (.L_HI(net43));
 sg13g2_tiehi _7442__44 (.L_HI(net44));
 sg13g2_tiehi _7407__45 (.L_HI(net45));
 sg13g2_tiehi _7441__46 (.L_HI(net46));
 sg13g2_tiehi _7406__47 (.L_HI(net47));
 sg13g2_tiehi _7440__48 (.L_HI(net48));
 sg13g2_tiehi _7405__49 (.L_HI(net49));
 sg13g2_tiehi _7439__50 (.L_HI(net50));
 sg13g2_tiehi _7404__51 (.L_HI(net51));
 sg13g2_tiehi _7438__52 (.L_HI(net52));
 sg13g2_tiehi _7403__53 (.L_HI(net53));
 sg13g2_tiehi _7437__54 (.L_HI(net54));
 sg13g2_tiehi _7402__55 (.L_HI(net55));
 sg13g2_tiehi _7436__56 (.L_HI(net56));
 sg13g2_tiehi _7401__57 (.L_HI(net57));
 sg13g2_tiehi _7435__58 (.L_HI(net58));
 sg13g2_tiehi _7400__59 (.L_HI(net59));
 sg13g2_tiehi _7434__60 (.L_HI(net60));
 sg13g2_tiehi _7399__61 (.L_HI(net61));
 sg13g2_tiehi _7433__62 (.L_HI(net62));
 sg13g2_tiehi _7398__63 (.L_HI(net63));
 sg13g2_tiehi _7397__64 (.L_HI(net64));
 sg13g2_tiehi _7396__65 (.L_HI(net65));
 sg13g2_tiehi _7395__66 (.L_HI(net66));
 sg13g2_tiehi _7394__67 (.L_HI(net67));
 sg13g2_tiehi _7393__68 (.L_HI(net68));
 sg13g2_tiehi _7392__69 (.L_HI(net69));
 sg13g2_tiehi _7391__70 (.L_HI(net70));
 sg13g2_tiehi _7390__71 (.L_HI(net71));
 sg13g2_tiehi _7389__72 (.L_HI(net72));
 sg13g2_tiehi _7388__73 (.L_HI(net73));
 sg13g2_tiehi _7387__74 (.L_HI(net74));
 sg13g2_tiehi _7432__75 (.L_HI(net75));
 sg13g2_tiehi _7431__76 (.L_HI(net76));
 sg13g2_tiehi _7430__77 (.L_HI(net77));
 sg13g2_tiehi _7429__78 (.L_HI(net78));
 sg13g2_tiehi _7428__79 (.L_HI(net79));
 sg13g2_tiehi _7427__80 (.L_HI(net80));
 sg13g2_tiehi _7386__81 (.L_HI(net81));
 sg13g2_tiehi _7426__82 (.L_HI(net82));
 sg13g2_tiehi _7425__83 (.L_HI(net83));
 sg13g2_tiehi _7424__84 (.L_HI(net84));
 sg13g2_tiehi _7423__85 (.L_HI(net85));
 sg13g2_tiehi _7453__86 (.L_HI(net86));
 sg13g2_tiehi _7422__87 (.L_HI(net87));
 sg13g2_tiehi _7458__88 (.L_HI(net88));
 sg13g2_tiehi _7421__89 (.L_HI(net89));
 sg13g2_tiehi _7452__90 (.L_HI(net90));
 sg13g2_tiehi _7420__91 (.L_HI(net91));
 sg13g2_tiehi _7446__92 (.L_HI(net92));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_5 (.L_LO(net5));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_6 (.L_LO(net6));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_7 (.L_LO(net7));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_8 (.L_LO(net8));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_9 (.L_LO(net9));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_10 (.L_LO(net10));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_11 (.L_LO(net11));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_12 (.L_LO(net12));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_13 (.L_LO(net13));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_14 (.L_LO(net14));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_15 (.L_LO(net15));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_16 (.L_LO(net16));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_17 (.L_LO(net17));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_18 (.L_LO(net18));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_19 (.L_LO(net19));
 sg13g2_tiehi _7455__20 (.L_HI(net20));
 sg13g2_buf_2 _7548_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _7549_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout1976 (.A(_3309_),
    .X(net1976));
 sg13g2_buf_4 fanout1977 (.X(net1977),
    .A(_3214_));
 sg13g2_buf_2 fanout1978 (.A(net1979),
    .X(net1978));
 sg13g2_buf_4 fanout1979 (.X(net1979),
    .A(net1980));
 sg13g2_buf_4 fanout1980 (.X(net1980),
    .A(_3213_));
 sg13g2_buf_8 fanout1981 (.A(_3432_),
    .X(net1981));
 sg13g2_buf_8 fanout1982 (.A(_3374_),
    .X(net1982));
 sg13g2_buf_4 fanout1983 (.X(net1983),
    .A(_3311_));
 sg13g2_buf_8 fanout1984 (.A(_3310_),
    .X(net1984));
 sg13g2_buf_4 fanout1985 (.X(net1985),
    .A(_3301_));
 sg13g2_buf_2 fanout1986 (.A(_1479_),
    .X(net1986));
 sg13g2_buf_4 fanout1987 (.X(net1987),
    .A(_1478_));
 sg13g2_buf_2 fanout1988 (.A(_1471_),
    .X(net1988));
 sg13g2_buf_2 fanout1989 (.A(_1469_),
    .X(net1989));
 sg13g2_buf_1 fanout1990 (.A(_1469_),
    .X(net1990));
 sg13g2_buf_4 fanout1991 (.X(net1991),
    .A(_1288_));
 sg13g2_buf_4 fanout1992 (.X(net1992),
    .A(_1057_));
 sg13g2_buf_4 fanout1993 (.X(net1993),
    .A(_0750_));
 sg13g2_buf_2 fanout1994 (.A(_0731_),
    .X(net1994));
 sg13g2_buf_8 fanout1995 (.A(_0640_),
    .X(net1995));
 sg13g2_buf_4 fanout1996 (.X(net1996),
    .A(_0547_));
 sg13g2_buf_4 fanout1997 (.X(net1997),
    .A(_0474_));
 sg13g2_buf_4 fanout1998 (.X(net1998),
    .A(net1999));
 sg13g2_buf_2 fanout1999 (.A(_0323_),
    .X(net1999));
 sg13g2_buf_4 fanout2000 (.X(net2000),
    .A(_0321_));
 sg13g2_buf_4 fanout2001 (.X(net2001),
    .A(_0299_));
 sg13g2_buf_2 fanout2002 (.A(_0299_),
    .X(net2002));
 sg13g2_buf_4 fanout2003 (.X(net2003),
    .A(_0295_));
 sg13g2_buf_2 fanout2004 (.A(_0295_),
    .X(net2004));
 sg13g2_buf_2 fanout2005 (.A(net2006),
    .X(net2005));
 sg13g2_buf_1 fanout2006 (.A(net2007),
    .X(net2006));
 sg13g2_buf_2 fanout2007 (.A(net2008),
    .X(net2007));
 sg13g2_buf_4 fanout2008 (.X(net2008),
    .A(_0253_));
 sg13g2_buf_4 fanout2009 (.X(net2009),
    .A(_3578_));
 sg13g2_buf_2 fanout2010 (.A(_3456_),
    .X(net2010));
 sg13g2_buf_4 fanout2011 (.X(net2011),
    .A(net2012));
 sg13g2_buf_4 fanout2012 (.X(net2012),
    .A(_3442_));
 sg13g2_buf_4 fanout2013 (.X(net2013),
    .A(net2015));
 sg13g2_buf_2 fanout2014 (.A(net2015),
    .X(net2014));
 sg13g2_buf_2 fanout2015 (.A(net2016),
    .X(net2015));
 sg13g2_buf_4 fanout2016 (.X(net2016),
    .A(_3434_));
 sg13g2_buf_4 fanout2017 (.X(net2017),
    .A(_3395_));
 sg13g2_buf_4 fanout2018 (.X(net2018),
    .A(net2019));
 sg13g2_buf_4 fanout2019 (.X(net2019),
    .A(_3376_));
 sg13g2_buf_2 fanout2020 (.A(_3285_),
    .X(net2020));
 sg13g2_buf_2 fanout2021 (.A(_3263_),
    .X(net2021));
 sg13g2_buf_4 fanout2022 (.X(net2022),
    .A(_3252_));
 sg13g2_buf_4 fanout2023 (.X(net2023),
    .A(_3252_));
 sg13g2_buf_4 fanout2024 (.X(net2024),
    .A(_3247_));
 sg13g2_buf_4 fanout2025 (.X(net2025),
    .A(_3204_));
 sg13g2_buf_2 fanout2026 (.A(net2027),
    .X(net2026));
 sg13g2_buf_4 fanout2027 (.X(net2027),
    .A(_3202_));
 sg13g2_buf_4 fanout2028 (.X(net2028),
    .A(_3181_));
 sg13g2_buf_2 fanout2029 (.A(_3137_),
    .X(net2029));
 sg13g2_buf_4 fanout2030 (.X(net2030),
    .A(net2032));
 sg13g2_buf_2 fanout2031 (.A(net2032),
    .X(net2031));
 sg13g2_buf_4 fanout2032 (.X(net2032),
    .A(_3134_));
 sg13g2_buf_4 fanout2033 (.X(net2033),
    .A(_3090_));
 sg13g2_buf_4 fanout2034 (.X(net2034),
    .A(_3074_));
 sg13g2_buf_8 fanout2035 (.A(_3073_),
    .X(net2035));
 sg13g2_buf_4 fanout2036 (.X(net2036),
    .A(_3073_));
 sg13g2_buf_4 fanout2037 (.X(net2037),
    .A(net2038));
 sg13g2_buf_4 fanout2038 (.X(net2038),
    .A(net2039));
 sg13g2_buf_4 fanout2039 (.X(net2039),
    .A(_3072_));
 sg13g2_buf_8 fanout2040 (.A(net2041),
    .X(net2040));
 sg13g2_buf_8 fanout2041 (.A(_3024_),
    .X(net2041));
 sg13g2_buf_4 fanout2042 (.X(net2042),
    .A(_2806_));
 sg13g2_buf_2 fanout2043 (.A(_2806_),
    .X(net2043));
 sg13g2_buf_2 fanout2044 (.A(_2636_),
    .X(net2044));
 sg13g2_buf_4 fanout2045 (.X(net2045),
    .A(_2625_));
 sg13g2_buf_2 fanout2046 (.A(net2048),
    .X(net2046));
 sg13g2_buf_2 fanout2047 (.A(net2048),
    .X(net2047));
 sg13g2_buf_4 fanout2048 (.X(net2048),
    .A(net2049));
 sg13g2_buf_4 fanout2049 (.X(net2049),
    .A(_2405_));
 sg13g2_buf_2 fanout2050 (.A(_2097_),
    .X(net2050));
 sg13g2_buf_1 fanout2051 (.A(_2097_),
    .X(net2051));
 sg13g2_buf_4 fanout2052 (.X(net2052),
    .A(net2053));
 sg13g2_buf_4 fanout2053 (.X(net2053),
    .A(_0737_));
 sg13g2_buf_4 fanout2054 (.X(net2054),
    .A(_3342_));
 sg13g2_buf_4 fanout2055 (.X(net2055),
    .A(_3217_));
 sg13g2_buf_4 fanout2056 (.X(net2056),
    .A(_3178_));
 sg13g2_buf_2 fanout2057 (.A(_3178_),
    .X(net2057));
 sg13g2_buf_4 fanout2058 (.X(net2058),
    .A(net2059));
 sg13g2_buf_4 fanout2059 (.X(net2059),
    .A(net2060));
 sg13g2_buf_8 fanout2060 (.A(_3177_),
    .X(net2060));
 sg13g2_buf_4 fanout2061 (.X(net2061),
    .A(_3165_));
 sg13g2_buf_4 fanout2062 (.X(net2062),
    .A(_3148_));
 sg13g2_buf_4 fanout2063 (.X(net2063),
    .A(_3128_));
 sg13g2_buf_4 fanout2064 (.X(net2064),
    .A(_3128_));
 sg13g2_buf_4 fanout2065 (.X(net2065),
    .A(_3123_));
 sg13g2_buf_2 fanout2066 (.A(_3123_),
    .X(net2066));
 sg13g2_buf_4 fanout2067 (.X(net2067),
    .A(_3119_));
 sg13g2_buf_4 fanout2068 (.X(net2068),
    .A(_3117_));
 sg13g2_buf_4 fanout2069 (.X(net2069),
    .A(_3116_));
 sg13g2_buf_4 fanout2070 (.X(net2070),
    .A(_3100_));
 sg13g2_buf_2 fanout2071 (.A(_3100_),
    .X(net2071));
 sg13g2_buf_4 fanout2072 (.X(net2072),
    .A(_3099_));
 sg13g2_buf_4 fanout2073 (.X(net2073),
    .A(_3099_));
 sg13g2_buf_8 fanout2074 (.A(_3029_),
    .X(net2074));
 sg13g2_buf_8 fanout2075 (.A(_2901_),
    .X(net2075));
 sg13g2_buf_4 fanout2076 (.X(net2076),
    .A(_2427_));
 sg13g2_buf_4 fanout2077 (.X(net2077),
    .A(_2372_));
 sg13g2_buf_4 fanout2078 (.X(net2078),
    .A(_2317_));
 sg13g2_buf_4 fanout2079 (.X(net2079),
    .A(_2064_));
 sg13g2_buf_4 fanout2080 (.X(net2080),
    .A(_2020_));
 sg13g2_buf_4 fanout2081 (.X(net2081),
    .A(net2082));
 sg13g2_buf_8 fanout2082 (.A(_2009_),
    .X(net2082));
 sg13g2_buf_4 fanout2083 (.X(net2083),
    .A(net2084));
 sg13g2_buf_4 fanout2084 (.X(net2084),
    .A(_1932_));
 sg13g2_buf_4 fanout2085 (.X(net2085),
    .A(net2087));
 sg13g2_buf_2 fanout2086 (.A(net2087),
    .X(net2086));
 sg13g2_buf_8 fanout2087 (.A(_1921_),
    .X(net2087));
 sg13g2_buf_4 fanout2088 (.X(net2088),
    .A(_1800_));
 sg13g2_buf_4 fanout2089 (.X(net2089),
    .A(net2091));
 sg13g2_buf_2 fanout2090 (.A(net2091),
    .X(net2090));
 sg13g2_buf_2 fanout2091 (.A(net2094),
    .X(net2091));
 sg13g2_buf_2 fanout2092 (.A(net2094),
    .X(net2092));
 sg13g2_buf_4 fanout2093 (.X(net2093),
    .A(net2094));
 sg13g2_buf_2 fanout2094 (.A(net2100),
    .X(net2094));
 sg13g2_buf_2 fanout2095 (.A(net2096),
    .X(net2095));
 sg13g2_buf_4 fanout2096 (.X(net2096),
    .A(net2100));
 sg13g2_buf_2 fanout2097 (.A(net2099),
    .X(net2097));
 sg13g2_buf_1 fanout2098 (.A(net2099),
    .X(net2098));
 sg13g2_buf_4 fanout2099 (.X(net2099),
    .A(net2100));
 sg13g2_buf_2 fanout2100 (.A(net2132),
    .X(net2100));
 sg13g2_buf_2 fanout2101 (.A(net2102),
    .X(net2101));
 sg13g2_buf_4 fanout2102 (.X(net2102),
    .A(net2103));
 sg13g2_buf_4 fanout2103 (.X(net2103),
    .A(net2109));
 sg13g2_buf_4 fanout2104 (.X(net2104),
    .A(net2106));
 sg13g2_buf_4 fanout2105 (.X(net2105),
    .A(net2106));
 sg13g2_buf_4 fanout2106 (.X(net2106),
    .A(net2109));
 sg13g2_buf_4 fanout2107 (.X(net2107),
    .A(net2109));
 sg13g2_buf_2 fanout2108 (.A(net2109),
    .X(net2108));
 sg13g2_buf_2 fanout2109 (.A(net2132),
    .X(net2109));
 sg13g2_buf_2 fanout2110 (.A(net2114),
    .X(net2110));
 sg13g2_buf_1 fanout2111 (.A(net2114),
    .X(net2111));
 sg13g2_buf_2 fanout2112 (.A(net2114),
    .X(net2112));
 sg13g2_buf_4 fanout2113 (.X(net2113),
    .A(net2114));
 sg13g2_buf_1 fanout2114 (.A(net2125),
    .X(net2114));
 sg13g2_buf_4 fanout2115 (.X(net2115),
    .A(net2117));
 sg13g2_buf_4 fanout2116 (.X(net2116),
    .A(net2117));
 sg13g2_buf_2 fanout2117 (.A(net2125),
    .X(net2117));
 sg13g2_buf_4 fanout2118 (.X(net2118),
    .A(net2120));
 sg13g2_buf_2 fanout2119 (.A(net2120),
    .X(net2119));
 sg13g2_buf_4 fanout2120 (.X(net2120),
    .A(net2125));
 sg13g2_buf_2 fanout2121 (.A(net2122),
    .X(net2121));
 sg13g2_buf_2 fanout2122 (.A(net2125),
    .X(net2122));
 sg13g2_buf_4 fanout2123 (.X(net2123),
    .A(net2124));
 sg13g2_buf_4 fanout2124 (.X(net2124),
    .A(net2125));
 sg13g2_buf_4 fanout2125 (.X(net2125),
    .A(net2132));
 sg13g2_buf_2 fanout2126 (.A(net2127),
    .X(net2126));
 sg13g2_buf_4 fanout2127 (.X(net2127),
    .A(net2128));
 sg13g2_buf_4 fanout2128 (.X(net2128),
    .A(net2132));
 sg13g2_buf_2 fanout2129 (.A(net2131),
    .X(net2129));
 sg13g2_buf_2 fanout2130 (.A(net2131),
    .X(net2130));
 sg13g2_buf_2 fanout2131 (.A(net2132),
    .X(net2131));
 sg13g2_buf_4 fanout2132 (.X(net2132),
    .A(_1646_));
 sg13g2_buf_4 fanout2133 (.X(net2133),
    .A(net2134));
 sg13g2_buf_2 fanout2134 (.A(net2157),
    .X(net2134));
 sg13g2_buf_4 fanout2135 (.X(net2135),
    .A(net2136));
 sg13g2_buf_4 fanout2136 (.X(net2136),
    .A(net2139));
 sg13g2_buf_2 fanout2137 (.A(net2138),
    .X(net2137));
 sg13g2_buf_4 fanout2138 (.X(net2138),
    .A(net2139));
 sg13g2_buf_2 fanout2139 (.A(net2157),
    .X(net2139));
 sg13g2_buf_4 fanout2140 (.X(net2140),
    .A(net2147));
 sg13g2_buf_2 fanout2141 (.A(net2147),
    .X(net2141));
 sg13g2_buf_4 fanout2142 (.X(net2142),
    .A(net2144));
 sg13g2_buf_4 fanout2143 (.X(net2143),
    .A(net2144));
 sg13g2_buf_2 fanout2144 (.A(net2147),
    .X(net2144));
 sg13g2_buf_4 fanout2145 (.X(net2145),
    .A(net2146));
 sg13g2_buf_4 fanout2146 (.X(net2146),
    .A(net2147));
 sg13g2_buf_2 fanout2147 (.A(net2157),
    .X(net2147));
 sg13g2_buf_2 fanout2148 (.A(net2150),
    .X(net2148));
 sg13g2_buf_4 fanout2149 (.X(net2149),
    .A(net2151));
 sg13g2_buf_1 fanout2150 (.A(net2151),
    .X(net2150));
 sg13g2_buf_2 fanout2151 (.A(net2156),
    .X(net2151));
 sg13g2_buf_2 fanout2152 (.A(net2153),
    .X(net2152));
 sg13g2_buf_4 fanout2153 (.X(net2153),
    .A(net2155));
 sg13g2_buf_2 fanout2154 (.A(net2155),
    .X(net2154));
 sg13g2_buf_4 fanout2155 (.X(net2155),
    .A(net2156));
 sg13g2_buf_2 fanout2156 (.A(net2157),
    .X(net2156));
 sg13g2_buf_4 fanout2157 (.X(net2157),
    .A(_1635_));
 sg13g2_buf_4 fanout2158 (.X(net2158),
    .A(net2160));
 sg13g2_buf_2 fanout2159 (.A(net2160),
    .X(net2159));
 sg13g2_buf_2 fanout2160 (.A(net2165),
    .X(net2160));
 sg13g2_buf_2 fanout2161 (.A(net2165),
    .X(net2161));
 sg13g2_buf_2 fanout2162 (.A(net2165),
    .X(net2162));
 sg13g2_buf_2 fanout2163 (.A(net2164),
    .X(net2163));
 sg13g2_buf_2 fanout2164 (.A(net2165),
    .X(net2164));
 sg13g2_buf_1 fanout2165 (.A(net2172),
    .X(net2165));
 sg13g2_buf_4 fanout2166 (.X(net2166),
    .A(net2168));
 sg13g2_buf_1 fanout2167 (.A(net2168),
    .X(net2167));
 sg13g2_buf_2 fanout2168 (.A(net2172),
    .X(net2168));
 sg13g2_buf_4 fanout2169 (.X(net2169),
    .A(net2171));
 sg13g2_buf_4 fanout2170 (.X(net2170),
    .A(net2171));
 sg13g2_buf_4 fanout2171 (.X(net2171),
    .A(net2172));
 sg13g2_buf_4 fanout2172 (.X(net2172),
    .A(_1635_));
 sg13g2_buf_4 fanout2173 (.X(net2173),
    .A(net2176));
 sg13g2_buf_4 fanout2174 (.X(net2174),
    .A(net2176));
 sg13g2_buf_2 fanout2175 (.A(net2176),
    .X(net2175));
 sg13g2_buf_2 fanout2176 (.A(net2186),
    .X(net2176));
 sg13g2_buf_2 fanout2177 (.A(net2178),
    .X(net2177));
 sg13g2_buf_2 fanout2178 (.A(net2179),
    .X(net2178));
 sg13g2_buf_2 fanout2179 (.A(net2186),
    .X(net2179));
 sg13g2_buf_2 fanout2180 (.A(net2181),
    .X(net2180));
 sg13g2_buf_2 fanout2181 (.A(net2183),
    .X(net2181));
 sg13g2_buf_4 fanout2182 (.X(net2182),
    .A(net2183));
 sg13g2_buf_2 fanout2183 (.A(net2186),
    .X(net2183));
 sg13g2_buf_2 fanout2184 (.A(net2185),
    .X(net2184));
 sg13g2_buf_2 fanout2185 (.A(net2186),
    .X(net2185));
 sg13g2_buf_2 fanout2186 (.A(_1635_),
    .X(net2186));
 sg13g2_buf_2 fanout2187 (.A(net2188),
    .X(net2187));
 sg13g2_buf_2 fanout2188 (.A(_2780_),
    .X(net2188));
 sg13g2_buf_2 fanout2189 (.A(net2190),
    .X(net2189));
 sg13g2_buf_4 fanout2190 (.X(net2190),
    .A(net2191));
 sg13g2_buf_2 fanout2191 (.A(_2780_),
    .X(net2191));
 sg13g2_buf_4 fanout2192 (.X(net2192),
    .A(net2193));
 sg13g2_buf_4 fanout2193 (.X(net2193),
    .A(net2194));
 sg13g2_buf_8 fanout2194 (.A(_3282_),
    .X(net2194));
 sg13g2_buf_4 fanout2195 (.X(net2195),
    .A(net2196));
 sg13g2_buf_8 fanout2196 (.A(net2198),
    .X(net2196));
 sg13g2_buf_8 fanout2197 (.A(net2198),
    .X(net2197));
 sg13g2_buf_4 fanout2198 (.X(net2198),
    .A(_3281_));
 sg13g2_buf_8 fanout2199 (.A(net2201),
    .X(net2199));
 sg13g2_buf_8 fanout2200 (.A(net2201),
    .X(net2200));
 sg13g2_buf_8 fanout2201 (.A(_3216_),
    .X(net2201));
 sg13g2_buf_4 fanout2202 (.X(net2202),
    .A(net2204));
 sg13g2_buf_4 fanout2203 (.X(net2203),
    .A(net2204));
 sg13g2_buf_4 fanout2204 (.X(net2204),
    .A(_3215_));
 sg13g2_buf_4 fanout2205 (.X(net2205),
    .A(net2207));
 sg13g2_buf_2 fanout2206 (.A(net2207),
    .X(net2206));
 sg13g2_buf_8 fanout2207 (.A(_3215_),
    .X(net2207));
 sg13g2_buf_8 fanout2208 (.A(_3152_),
    .X(net2208));
 sg13g2_buf_4 fanout2209 (.X(net2209),
    .A(net2210));
 sg13g2_buf_4 fanout2210 (.X(net2210),
    .A(_3143_));
 sg13g2_buf_4 fanout2211 (.X(net2211),
    .A(_3127_));
 sg13g2_buf_4 fanout2212 (.X(net2212),
    .A(net2213));
 sg13g2_buf_4 fanout2213 (.X(net2213),
    .A(_3126_));
 sg13g2_buf_4 fanout2214 (.X(net2214),
    .A(_3121_));
 sg13g2_buf_4 fanout2215 (.X(net2215),
    .A(_3078_));
 sg13g2_buf_4 fanout2216 (.X(net2216),
    .A(_2972_));
 sg13g2_buf_8 fanout2217 (.A(_2963_),
    .X(net2217));
 sg13g2_buf_4 fanout2218 (.X(net2218),
    .A(_2963_));
 sg13g2_buf_4 fanout2219 (.X(net2219),
    .A(net2220));
 sg13g2_buf_4 fanout2220 (.X(net2220),
    .A(_2954_));
 sg13g2_buf_4 fanout2221 (.X(net2221),
    .A(_2844_));
 sg13g2_buf_8 fanout2222 (.A(_2767_),
    .X(net2222));
 sg13g2_buf_8 fanout2223 (.A(_2757_),
    .X(net2223));
 sg13g2_buf_8 fanout2224 (.A(_2658_),
    .X(net2224));
 sg13g2_buf_2 fanout2225 (.A(_2658_),
    .X(net2225));
 sg13g2_buf_4 fanout2226 (.X(net2226),
    .A(_2361_));
 sg13g2_buf_4 fanout2227 (.X(net2227),
    .A(_2361_));
 sg13g2_buf_8 fanout2228 (.A(net2229),
    .X(net2228));
 sg13g2_buf_8 fanout2229 (.A(_2350_),
    .X(net2229));
 sg13g2_buf_4 fanout2230 (.X(net2230),
    .A(net2231));
 sg13g2_buf_4 fanout2231 (.X(net2231),
    .A(_2295_));
 sg13g2_buf_8 fanout2232 (.A(_2284_),
    .X(net2232));
 sg13g2_buf_4 fanout2233 (.X(net2233),
    .A(_2284_));
 sg13g2_buf_8 fanout2234 (.A(_2207_),
    .X(net2234));
 sg13g2_buf_4 fanout2235 (.X(net2235),
    .A(_2196_));
 sg13g2_buf_4 fanout2236 (.X(net2236),
    .A(_2053_));
 sg13g2_buf_4 fanout2237 (.X(net2237),
    .A(_2053_));
 sg13g2_buf_4 fanout2238 (.X(net2238),
    .A(_2042_));
 sg13g2_buf_4 fanout2239 (.X(net2239),
    .A(_2042_));
 sg13g2_buf_4 fanout2240 (.X(net2240),
    .A(net2241));
 sg13g2_buf_4 fanout2241 (.X(net2241),
    .A(net2243));
 sg13g2_buf_8 fanout2242 (.A(net2243),
    .X(net2242));
 sg13g2_buf_2 fanout2243 (.A(_1910_),
    .X(net2243));
 sg13g2_buf_4 fanout2244 (.X(net2244),
    .A(_1899_));
 sg13g2_buf_8 fanout2245 (.A(_1844_),
    .X(net2245));
 sg13g2_buf_4 fanout2246 (.X(net2246),
    .A(net2247));
 sg13g2_buf_8 fanout2247 (.A(_1789_),
    .X(net2247));
 sg13g2_buf_4 fanout2248 (.X(net2248),
    .A(net2249));
 sg13g2_buf_8 fanout2249 (.A(_1778_),
    .X(net2249));
 sg13g2_buf_4 fanout2250 (.X(net2250),
    .A(net2255));
 sg13g2_buf_2 fanout2251 (.A(net2255),
    .X(net2251));
 sg13g2_buf_4 fanout2252 (.X(net2252),
    .A(net2255));
 sg13g2_buf_4 fanout2253 (.X(net2253),
    .A(net2255));
 sg13g2_buf_4 fanout2254 (.X(net2254),
    .A(net2255));
 sg13g2_buf_4 fanout2255 (.X(net2255),
    .A(net2272));
 sg13g2_buf_4 fanout2256 (.X(net2256),
    .A(net2257));
 sg13g2_buf_4 fanout2257 (.X(net2257),
    .A(net2272));
 sg13g2_buf_4 fanout2258 (.X(net2258),
    .A(net2260));
 sg13g2_buf_1 fanout2259 (.A(net2260),
    .X(net2259));
 sg13g2_buf_4 fanout2260 (.X(net2260),
    .A(net2272));
 sg13g2_buf_4 fanout2261 (.X(net2261),
    .A(net2262));
 sg13g2_buf_4 fanout2262 (.X(net2262),
    .A(net2267));
 sg13g2_buf_4 fanout2263 (.X(net2263),
    .A(net2264));
 sg13g2_buf_2 fanout2264 (.A(net2267),
    .X(net2264));
 sg13g2_buf_4 fanout2265 (.X(net2265),
    .A(net2267));
 sg13g2_buf_4 fanout2266 (.X(net2266),
    .A(net2267));
 sg13g2_buf_2 fanout2267 (.A(net2272),
    .X(net2267));
 sg13g2_buf_4 fanout2268 (.X(net2268),
    .A(net2271));
 sg13g2_buf_4 fanout2269 (.X(net2269),
    .A(net2270));
 sg13g2_buf_4 fanout2270 (.X(net2270),
    .A(net2271));
 sg13g2_buf_4 fanout2271 (.X(net2271),
    .A(net2272));
 sg13g2_buf_4 fanout2272 (.X(net2272),
    .A(_1745_));
 sg13g2_buf_2 fanout2273 (.A(net2274),
    .X(net2273));
 sg13g2_buf_4 fanout2274 (.X(net2274),
    .A(net2276));
 sg13g2_buf_4 fanout2275 (.X(net2275),
    .A(net2276));
 sg13g2_buf_4 fanout2276 (.X(net2276),
    .A(net2281));
 sg13g2_buf_4 fanout2277 (.X(net2277),
    .A(net2278));
 sg13g2_buf_4 fanout2278 (.X(net2278),
    .A(net2281));
 sg13g2_buf_4 fanout2279 (.X(net2279),
    .A(net2281));
 sg13g2_buf_2 fanout2280 (.A(net2281),
    .X(net2280));
 sg13g2_buf_4 fanout2281 (.X(net2281),
    .A(_1734_));
 sg13g2_buf_4 fanout2282 (.X(net2282),
    .A(net2283));
 sg13g2_buf_4 fanout2283 (.X(net2283),
    .A(net2288));
 sg13g2_buf_4 fanout2284 (.X(net2284),
    .A(net2287));
 sg13g2_buf_2 fanout2285 (.A(net2287),
    .X(net2285));
 sg13g2_buf_4 fanout2286 (.X(net2286),
    .A(net2287));
 sg13g2_buf_2 fanout2287 (.A(net2288),
    .X(net2287));
 sg13g2_buf_4 fanout2288 (.X(net2288),
    .A(net2293));
 sg13g2_buf_4 fanout2289 (.X(net2289),
    .A(net2290));
 sg13g2_buf_2 fanout2290 (.A(net2293),
    .X(net2290));
 sg13g2_buf_4 fanout2291 (.X(net2291),
    .A(net2293));
 sg13g2_buf_1 fanout2292 (.A(net2293),
    .X(net2292));
 sg13g2_buf_2 fanout2293 (.A(_1734_),
    .X(net2293));
 sg13g2_buf_4 fanout2294 (.X(net2294),
    .A(net2299));
 sg13g2_buf_4 fanout2295 (.X(net2295),
    .A(net2299));
 sg13g2_buf_4 fanout2296 (.X(net2296),
    .A(net2298));
 sg13g2_buf_2 fanout2297 (.A(net2298),
    .X(net2297));
 sg13g2_buf_4 fanout2298 (.X(net2298),
    .A(net2299));
 sg13g2_buf_4 fanout2299 (.X(net2299),
    .A(_1261_));
 sg13g2_buf_4 fanout2300 (.X(net2300),
    .A(net2301));
 sg13g2_buf_8 fanout2301 (.A(_1250_),
    .X(net2301));
 sg13g2_buf_4 fanout2302 (.X(net2302),
    .A(net2303));
 sg13g2_buf_4 fanout2303 (.X(net2303),
    .A(_1250_));
 sg13g2_buf_4 fanout2304 (.X(net2304),
    .A(_2745_));
 sg13g2_buf_8 fanout2305 (.A(_3461_),
    .X(net2305));
 sg13g2_buf_8 fanout2306 (.A(net2307),
    .X(net2306));
 sg13g2_buf_8 fanout2307 (.A(_3453_),
    .X(net2307));
 sg13g2_buf_8 fanout2308 (.A(_3450_),
    .X(net2308));
 sg13g2_buf_8 fanout2309 (.A(_3449_),
    .X(net2309));
 sg13g2_buf_4 fanout2310 (.X(net2310),
    .A(_3449_));
 sg13g2_buf_4 fanout2311 (.X(net2311),
    .A(net2312));
 sg13g2_buf_8 fanout2312 (.A(_3051_),
    .X(net2312));
 sg13g2_buf_4 fanout2313 (.X(net2313),
    .A(net2317));
 sg13g2_buf_4 fanout2314 (.X(net2314),
    .A(net2317));
 sg13g2_buf_4 fanout2315 (.X(net2315),
    .A(net2316));
 sg13g2_buf_4 fanout2316 (.X(net2316),
    .A(net2317));
 sg13g2_buf_4 fanout2317 (.X(net2317),
    .A(_3050_));
 sg13g2_buf_4 fanout2318 (.X(net2318),
    .A(net2319));
 sg13g2_buf_4 fanout2319 (.X(net2319),
    .A(net2320));
 sg13g2_buf_8 fanout2320 (.A(_3049_),
    .X(net2320));
 sg13g2_buf_2 fanout2321 (.A(net2322),
    .X(net2321));
 sg13g2_buf_2 fanout2322 (.A(net2323),
    .X(net2322));
 sg13g2_buf_4 fanout2323 (.X(net2323),
    .A(net2324));
 sg13g2_buf_2 fanout2324 (.A(_3049_),
    .X(net2324));
 sg13g2_buf_4 fanout2325 (.X(net2325),
    .A(net2327));
 sg13g2_buf_4 fanout2326 (.X(net2326),
    .A(net2327));
 sg13g2_buf_8 fanout2327 (.A(_3040_),
    .X(net2327));
 sg13g2_buf_4 fanout2328 (.X(net2328),
    .A(net2329));
 sg13g2_buf_8 fanout2329 (.A(_3039_),
    .X(net2329));
 sg13g2_buf_4 fanout2330 (.X(net2330),
    .A(_3016_));
 sg13g2_buf_4 fanout2331 (.X(net2331),
    .A(_3016_));
 sg13g2_buf_4 fanout2332 (.X(net2332),
    .A(net2334));
 sg13g2_buf_2 fanout2333 (.A(net2334),
    .X(net2333));
 sg13g2_buf_8 fanout2334 (.A(_3015_),
    .X(net2334));
 sg13g2_buf_4 fanout2335 (.X(net2335),
    .A(_3015_));
 sg13g2_buf_8 fanout2336 (.A(net2337),
    .X(net2336));
 sg13g2_buf_8 fanout2337 (.A(_2537_),
    .X(net2337));
 sg13g2_buf_4 fanout2338 (.X(net2338),
    .A(net2339));
 sg13g2_buf_4 fanout2339 (.X(net2339),
    .A(net2340));
 sg13g2_buf_8 fanout2340 (.A(_2526_),
    .X(net2340));
 sg13g2_buf_8 fanout2341 (.A(_2185_),
    .X(net2341));
 sg13g2_buf_4 fanout2342 (.X(net2342),
    .A(net2343));
 sg13g2_buf_4 fanout2343 (.X(net2343),
    .A(net2344));
 sg13g2_buf_8 fanout2344 (.A(_2174_),
    .X(net2344));
 sg13g2_buf_4 fanout2345 (.X(net2345),
    .A(net2348));
 sg13g2_buf_2 fanout2346 (.A(net2348),
    .X(net2346));
 sg13g2_buf_4 fanout2347 (.X(net2347),
    .A(net2348));
 sg13g2_buf_2 fanout2348 (.A(_1998_),
    .X(net2348));
 sg13g2_buf_4 fanout2349 (.X(net2349),
    .A(net2350));
 sg13g2_buf_4 fanout2350 (.X(net2350),
    .A(_1987_));
 sg13g2_buf_4 fanout2351 (.X(net2351),
    .A(net2352));
 sg13g2_buf_4 fanout2352 (.X(net2352),
    .A(_1976_));
 sg13g2_buf_8 fanout2353 (.A(_1965_),
    .X(net2353));
 sg13g2_buf_4 fanout2354 (.X(net2354),
    .A(_1965_));
 sg13g2_buf_4 fanout2355 (.X(net2355),
    .A(_1954_));
 sg13g2_buf_8 fanout2356 (.A(_1943_),
    .X(net2356));
 sg13g2_buf_4 fanout2357 (.X(net2357),
    .A(_1833_));
 sg13g2_buf_8 fanout2358 (.A(_1822_),
    .X(net2358));
 sg13g2_buf_4 fanout2359 (.X(net2359),
    .A(_1822_));
 sg13g2_buf_4 fanout2360 (.X(net2360),
    .A(net2361));
 sg13g2_buf_4 fanout2361 (.X(net2361),
    .A(net2365));
 sg13g2_buf_4 fanout2362 (.X(net2362),
    .A(net2365));
 sg13g2_buf_4 fanout2363 (.X(net2363),
    .A(net2365));
 sg13g2_buf_4 fanout2364 (.X(net2364),
    .A(net2365));
 sg13g2_buf_4 fanout2365 (.X(net2365),
    .A(_1767_));
 sg13g2_buf_4 fanout2366 (.X(net2366),
    .A(net2368));
 sg13g2_buf_2 fanout2367 (.A(net2368),
    .X(net2367));
 sg13g2_buf_2 fanout2368 (.A(net2369),
    .X(net2368));
 sg13g2_buf_4 fanout2369 (.X(net2369),
    .A(_1756_));
 sg13g2_buf_4 fanout2370 (.X(net2370),
    .A(net2371));
 sg13g2_buf_2 fanout2371 (.A(net2372),
    .X(net2371));
 sg13g2_buf_4 fanout2372 (.X(net2372),
    .A(_1756_));
 sg13g2_buf_4 fanout2373 (.X(net2373),
    .A(_1723_));
 sg13g2_buf_4 fanout2374 (.X(net2374),
    .A(_1723_));
 sg13g2_buf_4 fanout2375 (.X(net2375),
    .A(_1712_));
 sg13g2_buf_4 fanout2376 (.X(net2376),
    .A(net2387));
 sg13g2_buf_2 fanout2377 (.A(net2387),
    .X(net2377));
 sg13g2_buf_4 fanout2378 (.X(net2378),
    .A(net2379));
 sg13g2_buf_4 fanout2379 (.X(net2379),
    .A(net2381));
 sg13g2_buf_4 fanout2380 (.X(net2380),
    .A(net2381));
 sg13g2_buf_2 fanout2381 (.A(net2387),
    .X(net2381));
 sg13g2_buf_4 fanout2382 (.X(net2382),
    .A(net2387));
 sg13g2_buf_2 fanout2383 (.A(net2386),
    .X(net2383));
 sg13g2_buf_4 fanout2384 (.X(net2384),
    .A(net2385));
 sg13g2_buf_4 fanout2385 (.X(net2385),
    .A(net2386));
 sg13g2_buf_4 fanout2386 (.X(net2386),
    .A(net2387));
 sg13g2_buf_8 fanout2387 (.A(_1206_),
    .X(net2387));
 sg13g2_buf_4 fanout2388 (.X(net2388),
    .A(net2389));
 sg13g2_buf_2 fanout2389 (.A(net2390),
    .X(net2389));
 sg13g2_buf_4 fanout2390 (.X(net2390),
    .A(net2394));
 sg13g2_buf_2 fanout2391 (.A(net2393),
    .X(net2391));
 sg13g2_buf_2 fanout2392 (.A(net2393),
    .X(net2392));
 sg13g2_buf_4 fanout2393 (.X(net2393),
    .A(net2394));
 sg13g2_buf_2 fanout2394 (.A(_1195_),
    .X(net2394));
 sg13g2_buf_4 fanout2395 (.X(net2395),
    .A(net2401));
 sg13g2_buf_4 fanout2396 (.X(net2396),
    .A(net2401));
 sg13g2_buf_4 fanout2397 (.X(net2397),
    .A(net2398));
 sg13g2_buf_4 fanout2398 (.X(net2398),
    .A(net2401));
 sg13g2_buf_4 fanout2399 (.X(net2399),
    .A(net2401));
 sg13g2_buf_2 fanout2400 (.A(net2401),
    .X(net2400));
 sg13g2_buf_4 fanout2401 (.X(net2401),
    .A(_1195_));
 sg13g2_buf_4 fanout2402 (.X(net2402),
    .A(net2406));
 sg13g2_buf_4 fanout2403 (.X(net2403),
    .A(net2406));
 sg13g2_buf_8 fanout2404 (.A(net2406),
    .X(net2404));
 sg13g2_buf_2 fanout2405 (.A(net2406),
    .X(net2405));
 sg13g2_buf_4 fanout2406 (.X(net2406),
    .A(_2163_));
 sg13g2_buf_4 fanout2407 (.X(net2407),
    .A(net2408));
 sg13g2_buf_4 fanout2408 (.X(net2408),
    .A(net2409));
 sg13g2_buf_8 fanout2409 (.A(_2152_),
    .X(net2409));
 sg13g2_buf_2 fanout2410 (.A(net2411),
    .X(net2410));
 sg13g2_buf_2 fanout2411 (.A(net2413),
    .X(net2411));
 sg13g2_buf_4 fanout2412 (.X(net2412),
    .A(net2413));
 sg13g2_buf_2 fanout2413 (.A(net2415),
    .X(net2413));
 sg13g2_buf_4 fanout2414 (.X(net2414),
    .A(net2415));
 sg13g2_buf_2 fanout2415 (.A(_2152_),
    .X(net2415));
 sg13g2_buf_4 fanout2416 (.X(net2416),
    .A(net2417));
 sg13g2_buf_4 fanout2417 (.X(net2417),
    .A(net2420));
 sg13g2_buf_4 fanout2418 (.X(net2418),
    .A(net2419));
 sg13g2_buf_4 fanout2419 (.X(net2419),
    .A(net2420));
 sg13g2_buf_8 fanout2420 (.A(_2141_),
    .X(net2420));
 sg13g2_buf_4 fanout2421 (.X(net2421),
    .A(net2423));
 sg13g2_buf_2 fanout2422 (.A(net2423),
    .X(net2422));
 sg13g2_buf_4 fanout2423 (.X(net2423),
    .A(net2424));
 sg13g2_buf_2 fanout2424 (.A(_2130_),
    .X(net2424));
 sg13g2_buf_4 fanout2425 (.X(net2425),
    .A(net2427));
 sg13g2_buf_4 fanout2426 (.X(net2426),
    .A(net2427));
 sg13g2_buf_4 fanout2427 (.X(net2427),
    .A(net2428));
 sg13g2_buf_4 fanout2428 (.X(net2428),
    .A(_2130_));
 sg13g2_buf_4 fanout2429 (.X(net2429),
    .A(net2433));
 sg13g2_buf_2 fanout2430 (.A(net2433),
    .X(net2430));
 sg13g2_buf_4 fanout2431 (.X(net2431),
    .A(net2433));
 sg13g2_buf_2 fanout2432 (.A(net2433),
    .X(net2432));
 sg13g2_buf_2 fanout2433 (.A(_2119_),
    .X(net2433));
 sg13g2_buf_4 fanout2434 (.X(net2434),
    .A(net2435));
 sg13g2_buf_4 fanout2435 (.X(net2435),
    .A(net2438));
 sg13g2_buf_4 fanout2436 (.X(net2436),
    .A(net2437));
 sg13g2_buf_4 fanout2437 (.X(net2437),
    .A(net2438));
 sg13g2_buf_2 fanout2438 (.A(_2119_),
    .X(net2438));
 sg13g2_buf_4 fanout2439 (.X(net2439),
    .A(net2441));
 sg13g2_buf_2 fanout2440 (.A(net2441),
    .X(net2440));
 sg13g2_buf_4 fanout2441 (.X(net2441),
    .A(net2442));
 sg13g2_buf_4 fanout2442 (.X(net2442),
    .A(net2450));
 sg13g2_buf_4 fanout2443 (.X(net2443),
    .A(net2444));
 sg13g2_buf_4 fanout2444 (.X(net2444),
    .A(net2447));
 sg13g2_buf_4 fanout2445 (.X(net2445),
    .A(net2447));
 sg13g2_buf_2 fanout2446 (.A(net2447),
    .X(net2446));
 sg13g2_buf_4 fanout2447 (.X(net2447),
    .A(net2450));
 sg13g2_buf_4 fanout2448 (.X(net2448),
    .A(net2449));
 sg13g2_buf_8 fanout2449 (.A(net2450),
    .X(net2449));
 sg13g2_buf_4 fanout2450 (.X(net2450),
    .A(_2108_));
 sg13g2_buf_4 fanout2451 (.X(net2451),
    .A(net2452));
 sg13g2_buf_4 fanout2452 (.X(net2452),
    .A(_1701_));
 sg13g2_buf_4 fanout2453 (.X(net2453),
    .A(_1690_));
 sg13g2_buf_4 fanout2454 (.X(net2454),
    .A(_1690_));
 sg13g2_buf_4 fanout2455 (.X(net2455),
    .A(net2457));
 sg13g2_buf_2 fanout2456 (.A(net2457),
    .X(net2456));
 sg13g2_buf_4 fanout2457 (.X(net2457),
    .A(_1668_));
 sg13g2_buf_4 fanout2458 (.X(net2458),
    .A(net2459));
 sg13g2_buf_4 fanout2459 (.X(net2459),
    .A(net2460));
 sg13g2_buf_4 fanout2460 (.X(net2460),
    .A(_1657_));
 sg13g2_buf_4 fanout2461 (.X(net2461),
    .A(net2464));
 sg13g2_buf_4 fanout2462 (.X(net2462),
    .A(net2463));
 sg13g2_buf_4 fanout2463 (.X(net2463),
    .A(net2464));
 sg13g2_buf_4 fanout2464 (.X(net2464),
    .A(net2469));
 sg13g2_buf_4 fanout2465 (.X(net2465),
    .A(net2466));
 sg13g2_buf_4 fanout2466 (.X(net2466),
    .A(net2469));
 sg13g2_buf_4 fanout2467 (.X(net2467),
    .A(net2469));
 sg13g2_buf_2 fanout2468 (.A(net2469),
    .X(net2468));
 sg13g2_buf_4 fanout2469 (.X(net2469),
    .A(_1360_));
 sg13g2_buf_4 fanout2470 (.X(net2470),
    .A(net2472));
 sg13g2_buf_2 fanout2471 (.A(net2472),
    .X(net2471));
 sg13g2_buf_4 fanout2472 (.X(net2472),
    .A(net2482));
 sg13g2_buf_4 fanout2473 (.X(net2473),
    .A(net2475));
 sg13g2_buf_4 fanout2474 (.X(net2474),
    .A(net2475));
 sg13g2_buf_4 fanout2475 (.X(net2475),
    .A(net2482));
 sg13g2_buf_4 fanout2476 (.X(net2476),
    .A(net2479));
 sg13g2_buf_2 fanout2477 (.A(net2479),
    .X(net2477));
 sg13g2_buf_4 fanout2478 (.X(net2478),
    .A(net2479));
 sg13g2_buf_2 fanout2479 (.A(net2482),
    .X(net2479));
 sg13g2_buf_4 fanout2480 (.X(net2480),
    .A(net2481));
 sg13g2_buf_4 fanout2481 (.X(net2481),
    .A(net2482));
 sg13g2_buf_8 fanout2482 (.A(_1349_),
    .X(net2482));
 sg13g2_buf_4 fanout2483 (.X(net2483),
    .A(net2486));
 sg13g2_buf_2 fanout2484 (.A(net2486),
    .X(net2484));
 sg13g2_buf_4 fanout2485 (.X(net2485),
    .A(net2486));
 sg13g2_buf_4 fanout2486 (.X(net2486),
    .A(net2492));
 sg13g2_buf_4 fanout2487 (.X(net2487),
    .A(net2488));
 sg13g2_buf_4 fanout2488 (.X(net2488),
    .A(net2489));
 sg13g2_buf_2 fanout2489 (.A(net2492),
    .X(net2489));
 sg13g2_buf_4 fanout2490 (.X(net2490),
    .A(net2492));
 sg13g2_buf_2 fanout2491 (.A(net2492),
    .X(net2491));
 sg13g2_buf_2 fanout2492 (.A(_1283_),
    .X(net2492));
 sg13g2_buf_4 fanout2493 (.X(net2493),
    .A(net2496));
 sg13g2_buf_4 fanout2494 (.X(net2494),
    .A(net2496));
 sg13g2_buf_1 fanout2495 (.A(net2496),
    .X(net2495));
 sg13g2_buf_4 fanout2496 (.X(net2496),
    .A(_1283_));
 sg13g2_buf_4 fanout2497 (.X(net2497),
    .A(net2500));
 sg13g2_buf_4 fanout2498 (.X(net2498),
    .A(net2500));
 sg13g2_buf_2 fanout2499 (.A(net2500),
    .X(net2499));
 sg13g2_buf_4 fanout2500 (.X(net2500),
    .A(_1283_));
 sg13g2_buf_4 fanout2501 (.X(net2501),
    .A(net2503));
 sg13g2_buf_2 fanout2502 (.A(net2503),
    .X(net2502));
 sg13g2_buf_2 fanout2503 (.A(net2505),
    .X(net2503));
 sg13g2_buf_4 fanout2504 (.X(net2504),
    .A(net2505));
 sg13g2_buf_4 fanout2505 (.X(net2505),
    .A(_1272_));
 sg13g2_buf_2 fanout2506 (.A(net2507),
    .X(net2506));
 sg13g2_buf_2 fanout2507 (.A(net2511),
    .X(net2507));
 sg13g2_buf_4 fanout2508 (.X(net2508),
    .A(net2511));
 sg13g2_buf_1 fanout2509 (.A(net2511),
    .X(net2509));
 sg13g2_buf_4 fanout2510 (.X(net2510),
    .A(net2511));
 sg13g2_buf_4 fanout2511 (.X(net2511),
    .A(_1272_));
 sg13g2_buf_4 fanout2512 (.X(net2512),
    .A(net2514));
 sg13g2_buf_4 fanout2513 (.X(net2513),
    .A(net2519));
 sg13g2_buf_2 fanout2514 (.A(net2519),
    .X(net2514));
 sg13g2_buf_4 fanout2515 (.X(net2515),
    .A(net2517));
 sg13g2_buf_2 fanout2516 (.A(net2517),
    .X(net2516));
 sg13g2_buf_4 fanout2517 (.X(net2517),
    .A(net2518));
 sg13g2_buf_4 fanout2518 (.X(net2518),
    .A(net2519));
 sg13g2_buf_4 fanout2519 (.X(net2519),
    .A(_1272_));
 sg13g2_buf_4 fanout2520 (.X(net2520),
    .A(net2525));
 sg13g2_buf_4 fanout2521 (.X(net2521),
    .A(net2525));
 sg13g2_buf_4 fanout2522 (.X(net2522),
    .A(net2524));
 sg13g2_buf_4 fanout2523 (.X(net2523),
    .A(net2524));
 sg13g2_buf_2 fanout2524 (.A(net2525),
    .X(net2524));
 sg13g2_buf_4 fanout2525 (.X(net2525),
    .A(_1338_));
 sg13g2_buf_4 fanout2526 (.X(net2526),
    .A(net2528));
 sg13g2_buf_2 fanout2527 (.A(net2528),
    .X(net2527));
 sg13g2_buf_4 fanout2528 (.X(net2528),
    .A(_1338_));
 sg13g2_buf_4 fanout2529 (.X(net2529),
    .A(net2530));
 sg13g2_buf_4 fanout2530 (.X(net2530),
    .A(net2531));
 sg13g2_buf_4 fanout2531 (.X(net2531),
    .A(net2537));
 sg13g2_buf_4 fanout2532 (.X(net2532),
    .A(net2537));
 sg13g2_buf_2 fanout2533 (.A(net2537),
    .X(net2533));
 sg13g2_buf_4 fanout2534 (.X(net2534),
    .A(net2536));
 sg13g2_buf_2 fanout2535 (.A(net2536),
    .X(net2535));
 sg13g2_buf_2 fanout2536 (.A(net2537),
    .X(net2536));
 sg13g2_buf_2 fanout2537 (.A(_1338_),
    .X(net2537));
 sg13g2_buf_2 fanout2538 (.A(net2540),
    .X(net2538));
 sg13g2_buf_4 fanout2539 (.X(net2539),
    .A(net2540));
 sg13g2_buf_2 fanout2540 (.A(net2543),
    .X(net2540));
 sg13g2_buf_4 fanout2541 (.X(net2541),
    .A(net2542));
 sg13g2_buf_4 fanout2542 (.X(net2542),
    .A(net2543));
 sg13g2_buf_2 fanout2543 (.A(_1327_),
    .X(net2543));
 sg13g2_buf_4 fanout2544 (.X(net2544),
    .A(net2547));
 sg13g2_buf_4 fanout2545 (.X(net2545),
    .A(net2546));
 sg13g2_buf_2 fanout2546 (.A(net2547),
    .X(net2546));
 sg13g2_buf_2 fanout2547 (.A(_1327_),
    .X(net2547));
 sg13g2_buf_4 fanout2548 (.X(net2548),
    .A(net2552));
 sg13g2_buf_4 fanout2549 (.X(net2549),
    .A(net2551));
 sg13g2_buf_4 fanout2550 (.X(net2550),
    .A(net2551));
 sg13g2_buf_2 fanout2551 (.A(net2552),
    .X(net2551));
 sg13g2_buf_2 fanout2552 (.A(net2558),
    .X(net2552));
 sg13g2_buf_4 fanout2553 (.X(net2553),
    .A(net2558));
 sg13g2_buf_4 fanout2554 (.X(net2554),
    .A(net2557));
 sg13g2_buf_2 fanout2555 (.A(net2556),
    .X(net2555));
 sg13g2_buf_4 fanout2556 (.X(net2556),
    .A(net2557));
 sg13g2_buf_2 fanout2557 (.A(net2558),
    .X(net2557));
 sg13g2_buf_4 fanout2558 (.X(net2558),
    .A(_1327_));
 sg13g2_buf_4 fanout2559 (.X(net2559),
    .A(net2568));
 sg13g2_buf_4 fanout2560 (.X(net2560),
    .A(net2568));
 sg13g2_buf_2 fanout2561 (.A(net2562),
    .X(net2561));
 sg13g2_buf_4 fanout2562 (.X(net2562),
    .A(net2568));
 sg13g2_buf_4 fanout2563 (.X(net2563),
    .A(net2564));
 sg13g2_buf_4 fanout2564 (.X(net2564),
    .A(net2567));
 sg13g2_buf_4 fanout2565 (.X(net2565),
    .A(net2567));
 sg13g2_buf_1 fanout2566 (.A(net2567),
    .X(net2566));
 sg13g2_buf_2 fanout2567 (.A(net2568),
    .X(net2567));
 sg13g2_buf_4 fanout2568 (.X(net2568),
    .A(_1316_));
 sg13g2_buf_2 fanout2569 (.A(net2570),
    .X(net2569));
 sg13g2_buf_4 fanout2570 (.X(net2570),
    .A(net2573));
 sg13g2_buf_4 fanout2571 (.X(net2571),
    .A(net2573));
 sg13g2_buf_2 fanout2572 (.A(net2573),
    .X(net2572));
 sg13g2_buf_2 fanout2573 (.A(_1316_),
    .X(net2573));
 sg13g2_buf_4 fanout2574 (.X(net2574),
    .A(net2577));
 sg13g2_buf_4 fanout2575 (.X(net2575),
    .A(net2576));
 sg13g2_buf_4 fanout2576 (.X(net2576),
    .A(net2577));
 sg13g2_buf_4 fanout2577 (.X(net2577),
    .A(_1316_));
 sg13g2_buf_4 fanout2578 (.X(net2578),
    .A(net2580));
 sg13g2_buf_2 fanout2579 (.A(net2580),
    .X(net2579));
 sg13g2_buf_2 fanout2580 (.A(net2591),
    .X(net2580));
 sg13g2_buf_2 fanout2581 (.A(net2582),
    .X(net2581));
 sg13g2_buf_1 fanout2582 (.A(net2583),
    .X(net2582));
 sg13g2_buf_2 fanout2583 (.A(net2584),
    .X(net2583));
 sg13g2_buf_4 fanout2584 (.X(net2584),
    .A(net2591));
 sg13g2_buf_2 fanout2585 (.A(net2586),
    .X(net2585));
 sg13g2_buf_2 fanout2586 (.A(net2590),
    .X(net2586));
 sg13g2_buf_2 fanout2587 (.A(net2590),
    .X(net2587));
 sg13g2_buf_4 fanout2588 (.X(net2588),
    .A(net2589));
 sg13g2_buf_4 fanout2589 (.X(net2589),
    .A(net2590));
 sg13g2_buf_2 fanout2590 (.A(net2591),
    .X(net2590));
 sg13g2_buf_2 fanout2591 (.A(_1305_),
    .X(net2591));
 sg13g2_buf_4 fanout2592 (.X(net2592),
    .A(net2593));
 sg13g2_buf_4 fanout2593 (.X(net2593),
    .A(net2596));
 sg13g2_buf_4 fanout2594 (.X(net2594),
    .A(net2595));
 sg13g2_buf_4 fanout2595 (.X(net2595),
    .A(net2596));
 sg13g2_buf_4 fanout2596 (.X(net2596),
    .A(_1305_));
 sg13g2_buf_4 fanout2597 (.X(net2597),
    .A(net2600));
 sg13g2_buf_2 fanout2598 (.A(net2599),
    .X(net2598));
 sg13g2_buf_2 fanout2599 (.A(net2600),
    .X(net2599));
 sg13g2_buf_2 fanout2600 (.A(net2601),
    .X(net2600));
 sg13g2_buf_4 fanout2601 (.X(net2601),
    .A(_1305_));
 sg13g2_buf_2 fanout2602 (.A(_0658_),
    .X(net2602));
 sg13g2_buf_2 fanout2603 (.A(net2604),
    .X(net2603));
 sg13g2_buf_4 fanout2604 (.X(net2604),
    .A(\pix_y[6] ));
 sg13g2_buf_2 fanout2605 (.A(net164),
    .X(net2605));
 sg13g2_buf_2 fanout2606 (.A(\pix_y[5] ),
    .X(net2606));
 sg13g2_buf_4 fanout2607 (.X(net2607),
    .A(\pix_y[4] ));
 sg13g2_buf_2 fanout2608 (.A(net2609),
    .X(net2608));
 sg13g2_buf_2 fanout2609 (.A(\pix_y[3] ),
    .X(net2609));
 sg13g2_buf_2 fanout2610 (.A(net2611),
    .X(net2610));
 sg13g2_buf_2 fanout2611 (.A(\pix_y[2] ),
    .X(net2611));
 sg13g2_buf_2 fanout2612 (.A(\pix_y[1] ),
    .X(net2612));
 sg13g2_buf_4 fanout2613 (.X(net2613),
    .A(\pix_y[0] ));
 sg13g2_buf_2 fanout2614 (.A(net2615),
    .X(net2614));
 sg13g2_buf_4 fanout2615 (.X(net2615),
    .A(dir_y));
 sg13g2_buf_4 fanout2616 (.X(net2616),
    .A(net2617));
 sg13g2_buf_4 fanout2617 (.X(net2617),
    .A(dir_x));
 sg13g2_buf_2 fanout2618 (.A(net184),
    .X(net2618));
 sg13g2_buf_4 fanout2619 (.X(net2619),
    .A(net159));
 sg13g2_buf_4 fanout2620 (.X(net2620),
    .A(net136));
 sg13g2_buf_2 fanout2621 (.A(net163),
    .X(net2621));
 sg13g2_buf_4 fanout2622 (.X(net2622),
    .A(_0878_));
 sg13g2_buf_2 fanout2623 (.A(net2624),
    .X(net2623));
 sg13g2_buf_1 fanout2624 (.A(net2625),
    .X(net2624));
 sg13g2_buf_2 fanout2625 (.A(net2626),
    .X(net2625));
 sg13g2_buf_4 fanout2626 (.X(net2626),
    .A(net1));
 sg13g2_buf_4 fanout2627 (.X(net2627),
    .A(net2629));
 sg13g2_buf_1 fanout2628 (.A(net2629),
    .X(net2628));
 sg13g2_buf_2 fanout2629 (.A(net1),
    .X(net2629));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_tielo tt_um_arud4172_ROOTS_vga_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0014_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0008_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold3 (.A(_2984_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0011_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0049_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0009_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0070_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0010_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0062_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0002_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0047_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0012_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0037_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0013_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0027_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold16 (.A(\prev_y[6] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold17 (.A(\prev_y[9] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0061_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold19 (.A(\frame_divider[1] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold20 (.A(_2953_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold21 (.A(\prev_y[4] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0056_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold23 (.A(\prev_y[3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0005_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0048_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold26 (.A(\prev_y[8] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold27 (.A(\prev_y[5] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0057_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold29 (.A(\prev_y[2] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold30 (.A(\prev_y[7] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold31 (.A(\prev_y[1] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0053_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold33 (.A(\prev_y[0] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0052_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold35 (.A(\logo_top[9] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold36 (.A(\frame_counter[7] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0069_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold38 (.A(\logo_left[1] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold39 (.A(\logo_top[1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold40 (.A(\pix_x[2] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold41 (.A(_2747_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold42 (.A(\pix_x[9] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold43 (.A(_2758_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold44 (.A(\pix_x[6] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold45 (.A(_1020_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0000_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold47 (.A(\frame_counter[4] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0066_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold49 (.A(\color_index[2] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0051_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold51 (.A(\color_index[1] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold52 (.A(_2933_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold53 (.A(\pix_x[1] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold54 (.A(_2746_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold55 (.A(\logo_left[8] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0035_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold57 (.A(\frame_counter[3] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0065_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold59 (.A(\frame_counter[2] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0064_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold61 (.A(\logo_top[8] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold62 (.A(\frame_counter[5] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0067_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold64 (.A(\logo_left[9] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0036_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold66 (.A(\pix_y[9] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold67 (.A(\pix_x[7] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold68 (.A(_2756_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold69 (.A(\pix_x[3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold70 (.A(_2748_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold71 (.A(\pix_x[5] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold72 (.A(\pix_y[5] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold73 (.A(\logo_top[2] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold74 (.A(\logo_top[7] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0044_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold76 (.A(\logo_left[4] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0031_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold78 (.A(\logo_left[2] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold79 (.A(\logo_top[6] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold80 (.A(\pix_x[4] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold81 (.A(\pix_y[7] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold82 (.A(\logo_top[5] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold83 (.A(\logo_top[3] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold84 (.A(\logo_left[5] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold85 (.A(\logo_top[4] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold86 (.A(\frame_counter[6] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold87 (.A(\frame_counter[0] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold88 (.A(_2945_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0063_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pix_x[7] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold91 (.A(\color_index[0] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold92 (.A(\logo_left[3] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold93 (.A(\color_index[1] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold94 (.A(\color_index[2] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold95 (.A(\pix_x[1] ),
    .X(net187));
 sg13g2_antennanp ANTENNA_1 (.A(_0688_));
 sg13g2_antennanp ANTENNA_2 (.A(_1406_));
 sg13g2_antennanp ANTENNA_3 (.A(_1406_));
 sg13g2_antennanp ANTENNA_4 (.A(_1857_));
 sg13g2_antennanp ANTENNA_5 (.A(_3299_));
 sg13g2_antennanp ANTENNA_6 (.A(_3299_));
 sg13g2_antennanp ANTENNA_7 (.A(_3299_));
 sg13g2_antennanp ANTENNA_8 (.A(_3419_));
 sg13g2_antennanp ANTENNA_9 (.A(_3419_));
 sg13g2_antennanp ANTENNA_10 (.A(_3419_));
 sg13g2_antennanp ANTENNA_11 (.A(_3419_));
 sg13g2_antennanp ANTENNA_12 (.A(_3419_));
 sg13g2_antennanp ANTENNA_13 (.A(_3419_));
 sg13g2_antennanp ANTENNA_14 (.A(_3419_));
 sg13g2_antennanp ANTENNA_15 (.A(_3419_));
 sg13g2_antennanp ANTENNA_16 (.A(net2157));
 sg13g2_antennanp ANTENNA_17 (.A(net2157));
 sg13g2_antennanp ANTENNA_18 (.A(net2157));
 sg13g2_antennanp ANTENNA_19 (.A(net2157));
 sg13g2_antennanp ANTENNA_20 (.A(net2387));
 sg13g2_antennanp ANTENNA_21 (.A(net2387));
 sg13g2_antennanp ANTENNA_22 (.A(net2387));
 sg13g2_antennanp ANTENNA_23 (.A(net2387));
 sg13g2_antennanp ANTENNA_24 (.A(net2387));
 sg13g2_antennanp ANTENNA_25 (.A(net2387));
 sg13g2_antennanp ANTENNA_26 (.A(_0688_));
 sg13g2_antennanp ANTENNA_27 (.A(_1406_));
 sg13g2_antennanp ANTENNA_28 (.A(_1406_));
 sg13g2_antennanp ANTENNA_29 (.A(_1857_));
 sg13g2_antennanp ANTENNA_30 (.A(_3299_));
 sg13g2_antennanp ANTENNA_31 (.A(_3299_));
 sg13g2_antennanp ANTENNA_32 (.A(_3299_));
 sg13g2_antennanp ANTENNA_33 (.A(_3411_));
 sg13g2_antennanp ANTENNA_34 (.A(_3411_));
 sg13g2_antennanp ANTENNA_35 (.A(_3411_));
 sg13g2_antennanp ANTENNA_36 (.A(_3411_));
 sg13g2_antennanp ANTENNA_37 (.A(_3411_));
 sg13g2_antennanp ANTENNA_38 (.A(_3411_));
 sg13g2_antennanp ANTENNA_39 (.A(net2387));
 sg13g2_antennanp ANTENNA_40 (.A(net2387));
 sg13g2_antennanp ANTENNA_41 (.A(net2387));
 sg13g2_antennanp ANTENNA_42 (.A(net2387));
 sg13g2_antennanp ANTENNA_43 (.A(net2387));
 sg13g2_antennanp ANTENNA_44 (.A(net2387));
 sg13g2_antennanp ANTENNA_45 (.A(net2387));
 sg13g2_antennanp ANTENNA_46 (.A(net2387));
 sg13g2_antennanp ANTENNA_47 (.A(net2387));
 sg13g2_antennanp ANTENNA_48 (.A(net2387));
 sg13g2_antennanp ANTENNA_49 (.A(_0688_));
 sg13g2_antennanp ANTENNA_50 (.A(_1406_));
 sg13g2_antennanp ANTENNA_51 (.A(_1406_));
 sg13g2_antennanp ANTENNA_52 (.A(_1857_));
 sg13g2_antennanp ANTENNA_53 (.A(net2387));
 sg13g2_antennanp ANTENNA_54 (.A(net2387));
 sg13g2_antennanp ANTENNA_55 (.A(net2387));
 sg13g2_antennanp ANTENNA_56 (.A(net2387));
 sg13g2_antennanp ANTENNA_57 (.A(net2387));
 sg13g2_antennanp ANTENNA_58 (.A(net2387));
 sg13g2_antennanp ANTENNA_59 (.A(net2387));
 sg13g2_antennanp ANTENNA_60 (.A(net2387));
 sg13g2_antennanp ANTENNA_61 (.A(net2387));
 sg13g2_antennanp ANTENNA_62 (.A(net2387));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_4 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_decap_4 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_4 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_261 ();
 sg13g2_decap_8 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_decap_4 FILLER_6_282 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_decap_4 FILLER_6_292 ();
 sg13g2_fill_2 FILLER_6_296 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_fill_2 FILLER_6_339 ();
 sg13g2_fill_1 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_4 FILLER_6_358 ();
 sg13g2_fill_1 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_decap_8 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_6_414 ();
 sg13g2_fill_2 FILLER_6_421 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_536 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_4 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_4 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_151 ();
 sg13g2_decap_4 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_203 ();
 sg13g2_fill_2 FILLER_7_208 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_fill_2 FILLER_7_224 ();
 sg13g2_decap_4 FILLER_7_234 ();
 sg13g2_fill_2 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_255 ();
 sg13g2_fill_1 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_289 ();
 sg13g2_decap_4 FILLER_7_296 ();
 sg13g2_fill_1 FILLER_7_300 ();
 sg13g2_decap_8 FILLER_7_307 ();
 sg13g2_fill_2 FILLER_7_314 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_decap_4 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_fill_2 FILLER_7_360 ();
 sg13g2_fill_1 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_fill_2 FILLER_7_386 ();
 sg13g2_fill_2 FILLER_7_399 ();
 sg13g2_fill_1 FILLER_7_401 ();
 sg13g2_decap_4 FILLER_7_412 ();
 sg13g2_fill_1 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_decap_8 FILLER_7_429 ();
 sg13g2_decap_4 FILLER_7_436 ();
 sg13g2_decap_8 FILLER_7_445 ();
 sg13g2_decap_8 FILLER_7_452 ();
 sg13g2_decap_8 FILLER_7_459 ();
 sg13g2_fill_1 FILLER_7_466 ();
 sg13g2_decap_8 FILLER_7_479 ();
 sg13g2_decap_8 FILLER_7_486 ();
 sg13g2_decap_8 FILLER_7_493 ();
 sg13g2_decap_8 FILLER_7_500 ();
 sg13g2_fill_2 FILLER_7_507 ();
 sg13g2_fill_1 FILLER_7_509 ();
 sg13g2_decap_4 FILLER_7_514 ();
 sg13g2_fill_2 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_528 ();
 sg13g2_fill_2 FILLER_7_535 ();
 sg13g2_decap_8 FILLER_7_542 ();
 sg13g2_decap_8 FILLER_7_549 ();
 sg13g2_decap_8 FILLER_7_556 ();
 sg13g2_decap_8 FILLER_7_563 ();
 sg13g2_decap_8 FILLER_7_570 ();
 sg13g2_decap_8 FILLER_7_577 ();
 sg13g2_decap_8 FILLER_7_584 ();
 sg13g2_decap_8 FILLER_7_591 ();
 sg13g2_decap_8 FILLER_7_598 ();
 sg13g2_decap_8 FILLER_7_605 ();
 sg13g2_decap_8 FILLER_7_612 ();
 sg13g2_decap_8 FILLER_7_619 ();
 sg13g2_decap_8 FILLER_7_626 ();
 sg13g2_decap_8 FILLER_7_633 ();
 sg13g2_decap_8 FILLER_7_640 ();
 sg13g2_decap_8 FILLER_7_647 ();
 sg13g2_decap_8 FILLER_7_654 ();
 sg13g2_decap_8 FILLER_7_661 ();
 sg13g2_decap_8 FILLER_7_668 ();
 sg13g2_decap_8 FILLER_7_675 ();
 sg13g2_decap_8 FILLER_7_682 ();
 sg13g2_decap_8 FILLER_7_689 ();
 sg13g2_decap_8 FILLER_7_696 ();
 sg13g2_decap_8 FILLER_7_703 ();
 sg13g2_decap_8 FILLER_7_710 ();
 sg13g2_decap_8 FILLER_7_717 ();
 sg13g2_decap_8 FILLER_7_724 ();
 sg13g2_decap_8 FILLER_7_731 ();
 sg13g2_decap_8 FILLER_7_738 ();
 sg13g2_decap_8 FILLER_7_745 ();
 sg13g2_decap_8 FILLER_7_752 ();
 sg13g2_decap_8 FILLER_7_759 ();
 sg13g2_decap_8 FILLER_7_766 ();
 sg13g2_decap_8 FILLER_7_773 ();
 sg13g2_decap_8 FILLER_7_780 ();
 sg13g2_decap_8 FILLER_7_787 ();
 sg13g2_decap_8 FILLER_7_794 ();
 sg13g2_decap_8 FILLER_7_801 ();
 sg13g2_decap_8 FILLER_7_808 ();
 sg13g2_decap_8 FILLER_7_815 ();
 sg13g2_decap_8 FILLER_7_822 ();
 sg13g2_decap_8 FILLER_7_829 ();
 sg13g2_decap_8 FILLER_7_836 ();
 sg13g2_decap_8 FILLER_7_843 ();
 sg13g2_decap_8 FILLER_7_850 ();
 sg13g2_decap_4 FILLER_7_857 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_decap_4 FILLER_8_129 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_143 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_fill_1 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_176 ();
 sg13g2_decap_4 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_fill_2 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_198 ();
 sg13g2_decap_8 FILLER_8_204 ();
 sg13g2_decap_4 FILLER_8_211 ();
 sg13g2_fill_1 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_246 ();
 sg13g2_decap_8 FILLER_8_255 ();
 sg13g2_decap_8 FILLER_8_262 ();
 sg13g2_decap_4 FILLER_8_285 ();
 sg13g2_decap_4 FILLER_8_293 ();
 sg13g2_fill_1 FILLER_8_297 ();
 sg13g2_fill_2 FILLER_8_311 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_4 FILLER_8_363 ();
 sg13g2_fill_2 FILLER_8_367 ();
 sg13g2_fill_2 FILLER_8_374 ();
 sg13g2_fill_1 FILLER_8_376 ();
 sg13g2_fill_2 FILLER_8_382 ();
 sg13g2_fill_1 FILLER_8_384 ();
 sg13g2_fill_2 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_403 ();
 sg13g2_decap_4 FILLER_8_416 ();
 sg13g2_fill_1 FILLER_8_426 ();
 sg13g2_decap_4 FILLER_8_432 ();
 sg13g2_fill_1 FILLER_8_467 ();
 sg13g2_fill_2 FILLER_8_486 ();
 sg13g2_fill_1 FILLER_8_488 ();
 sg13g2_fill_2 FILLER_8_512 ();
 sg13g2_fill_1 FILLER_8_514 ();
 sg13g2_decap_4 FILLER_8_520 ();
 sg13g2_fill_2 FILLER_8_531 ();
 sg13g2_fill_2 FILLER_8_541 ();
 sg13g2_decap_4 FILLER_8_559 ();
 sg13g2_decap_8 FILLER_8_571 ();
 sg13g2_decap_8 FILLER_8_578 ();
 sg13g2_decap_8 FILLER_8_585 ();
 sg13g2_decap_8 FILLER_8_592 ();
 sg13g2_decap_8 FILLER_8_599 ();
 sg13g2_decap_8 FILLER_8_606 ();
 sg13g2_decap_8 FILLER_8_613 ();
 sg13g2_decap_8 FILLER_8_620 ();
 sg13g2_decap_8 FILLER_8_627 ();
 sg13g2_decap_8 FILLER_8_634 ();
 sg13g2_decap_8 FILLER_8_641 ();
 sg13g2_decap_8 FILLER_8_648 ();
 sg13g2_decap_8 FILLER_8_655 ();
 sg13g2_decap_8 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_669 ();
 sg13g2_decap_8 FILLER_8_676 ();
 sg13g2_decap_8 FILLER_8_683 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_8 FILLER_8_697 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_732 ();
 sg13g2_decap_8 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_8 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_767 ();
 sg13g2_decap_8 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_4 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_4 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_136 ();
 sg13g2_decap_4 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_152 ();
 sg13g2_decap_4 FILLER_9_180 ();
 sg13g2_fill_1 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_4 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_fill_2 FILLER_9_262 ();
 sg13g2_fill_1 FILLER_9_264 ();
 sg13g2_fill_2 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_4 FILLER_9_302 ();
 sg13g2_fill_1 FILLER_9_306 ();
 sg13g2_fill_2 FILLER_9_317 ();
 sg13g2_decap_4 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_328 ();
 sg13g2_decap_4 FILLER_9_342 ();
 sg13g2_fill_2 FILLER_9_346 ();
 sg13g2_decap_4 FILLER_9_353 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_decap_4 FILLER_9_369 ();
 sg13g2_decap_4 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_decap_4 FILLER_9_416 ();
 sg13g2_decap_8 FILLER_9_430 ();
 sg13g2_decap_4 FILLER_9_437 ();
 sg13g2_fill_1 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_4 FILLER_9_466 ();
 sg13g2_decap_8 FILLER_9_481 ();
 sg13g2_fill_2 FILLER_9_488 ();
 sg13g2_decap_8 FILLER_9_495 ();
 sg13g2_decap_8 FILLER_9_502 ();
 sg13g2_fill_2 FILLER_9_509 ();
 sg13g2_fill_1 FILLER_9_511 ();
 sg13g2_fill_2 FILLER_9_517 ();
 sg13g2_fill_1 FILLER_9_519 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_4 FILLER_9_544 ();
 sg13g2_fill_1 FILLER_9_548 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_fill_2 FILLER_9_567 ();
 sg13g2_fill_1 FILLER_9_569 ();
 sg13g2_decap_8 FILLER_9_578 ();
 sg13g2_decap_8 FILLER_9_585 ();
 sg13g2_decap_8 FILLER_9_592 ();
 sg13g2_decap_8 FILLER_9_599 ();
 sg13g2_decap_8 FILLER_9_606 ();
 sg13g2_decap_8 FILLER_9_613 ();
 sg13g2_decap_8 FILLER_9_620 ();
 sg13g2_decap_8 FILLER_9_627 ();
 sg13g2_decap_8 FILLER_9_634 ();
 sg13g2_decap_8 FILLER_9_641 ();
 sg13g2_decap_8 FILLER_9_648 ();
 sg13g2_decap_8 FILLER_9_655 ();
 sg13g2_decap_8 FILLER_9_662 ();
 sg13g2_decap_8 FILLER_9_669 ();
 sg13g2_decap_8 FILLER_9_676 ();
 sg13g2_decap_8 FILLER_9_683 ();
 sg13g2_decap_8 FILLER_9_690 ();
 sg13g2_decap_8 FILLER_9_697 ();
 sg13g2_decap_8 FILLER_9_704 ();
 sg13g2_decap_8 FILLER_9_711 ();
 sg13g2_decap_8 FILLER_9_718 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_decap_8 FILLER_9_732 ();
 sg13g2_decap_8 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_746 ();
 sg13g2_decap_8 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_760 ();
 sg13g2_decap_8 FILLER_9_767 ();
 sg13g2_decap_8 FILLER_9_774 ();
 sg13g2_decap_8 FILLER_9_781 ();
 sg13g2_decap_8 FILLER_9_788 ();
 sg13g2_decap_8 FILLER_9_795 ();
 sg13g2_decap_8 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_809 ();
 sg13g2_decap_8 FILLER_9_816 ();
 sg13g2_decap_8 FILLER_9_823 ();
 sg13g2_decap_8 FILLER_9_830 ();
 sg13g2_decap_8 FILLER_9_837 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_decap_8 FILLER_9_851 ();
 sg13g2_decap_4 FILLER_9_858 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_fill_2 FILLER_10_56 ();
 sg13g2_fill_1 FILLER_10_58 ();
 sg13g2_fill_1 FILLER_10_67 ();
 sg13g2_decap_4 FILLER_10_74 ();
 sg13g2_fill_1 FILLER_10_78 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_decap_4 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_decap_4 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_232 ();
 sg13g2_decap_4 FILLER_10_239 ();
 sg13g2_fill_2 FILLER_10_243 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_fill_2 FILLER_10_277 ();
 sg13g2_fill_2 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_301 ();
 sg13g2_decap_4 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_4 FILLER_10_367 ();
 sg13g2_fill_2 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_fill_2 FILLER_10_388 ();
 sg13g2_fill_1 FILLER_10_390 ();
 sg13g2_fill_2 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_436 ();
 sg13g2_decap_8 FILLER_10_443 ();
 sg13g2_decap_8 FILLER_10_450 ();
 sg13g2_fill_1 FILLER_10_457 ();
 sg13g2_decap_8 FILLER_10_475 ();
 sg13g2_fill_2 FILLER_10_482 ();
 sg13g2_fill_1 FILLER_10_484 ();
 sg13g2_fill_2 FILLER_10_503 ();
 sg13g2_fill_1 FILLER_10_505 ();
 sg13g2_decap_4 FILLER_10_510 ();
 sg13g2_fill_2 FILLER_10_514 ();
 sg13g2_decap_8 FILLER_10_521 ();
 sg13g2_fill_2 FILLER_10_528 ();
 sg13g2_fill_1 FILLER_10_530 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_fill_1 FILLER_10_546 ();
 sg13g2_fill_2 FILLER_10_551 ();
 sg13g2_fill_1 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_565 ();
 sg13g2_decap_4 FILLER_10_572 ();
 sg13g2_fill_1 FILLER_10_576 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_fill_2 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_642 ();
 sg13g2_decap_4 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_653 ();
 sg13g2_decap_8 FILLER_10_660 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_decap_8 FILLER_10_674 ();
 sg13g2_decap_8 FILLER_10_681 ();
 sg13g2_decap_8 FILLER_10_688 ();
 sg13g2_decap_8 FILLER_10_695 ();
 sg13g2_decap_8 FILLER_10_702 ();
 sg13g2_decap_8 FILLER_10_709 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_decap_8 FILLER_10_723 ();
 sg13g2_decap_8 FILLER_10_730 ();
 sg13g2_decap_8 FILLER_10_737 ();
 sg13g2_decap_8 FILLER_10_744 ();
 sg13g2_decap_8 FILLER_10_751 ();
 sg13g2_decap_8 FILLER_10_758 ();
 sg13g2_decap_8 FILLER_10_765 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_8 FILLER_10_842 ();
 sg13g2_decap_8 FILLER_10_849 ();
 sg13g2_decap_4 FILLER_10_856 ();
 sg13g2_fill_2 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_4 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_48 ();
 sg13g2_decap_8 FILLER_11_55 ();
 sg13g2_decap_4 FILLER_11_62 ();
 sg13g2_decap_8 FILLER_11_71 ();
 sg13g2_decap_8 FILLER_11_78 ();
 sg13g2_decap_4 FILLER_11_85 ();
 sg13g2_decap_8 FILLER_11_99 ();
 sg13g2_fill_1 FILLER_11_106 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_decap_4 FILLER_11_123 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_decap_4 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_143 ();
 sg13g2_decap_4 FILLER_11_150 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_fill_2 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_4 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_4 FILLER_11_234 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_4 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_fill_1 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_4 FILLER_11_333 ();
 sg13g2_decap_4 FILLER_11_351 ();
 sg13g2_fill_1 FILLER_11_355 ();
 sg13g2_decap_4 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_4 FILLER_11_393 ();
 sg13g2_fill_1 FILLER_11_397 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_decap_8 FILLER_11_428 ();
 sg13g2_fill_2 FILLER_11_435 ();
 sg13g2_decap_4 FILLER_11_440 ();
 sg13g2_fill_2 FILLER_11_444 ();
 sg13g2_decap_8 FILLER_11_451 ();
 sg13g2_fill_1 FILLER_11_458 ();
 sg13g2_decap_8 FILLER_11_486 ();
 sg13g2_fill_1 FILLER_11_493 ();
 sg13g2_fill_2 FILLER_11_511 ();
 sg13g2_decap_4 FILLER_11_541 ();
 sg13g2_fill_1 FILLER_11_545 ();
 sg13g2_fill_1 FILLER_11_555 ();
 sg13g2_fill_2 FILLER_11_561 ();
 sg13g2_decap_8 FILLER_11_573 ();
 sg13g2_decap_8 FILLER_11_597 ();
 sg13g2_decap_8 FILLER_11_604 ();
 sg13g2_decap_8 FILLER_11_611 ();
 sg13g2_fill_2 FILLER_11_618 ();
 sg13g2_fill_2 FILLER_11_625 ();
 sg13g2_decap_4 FILLER_11_649 ();
 sg13g2_fill_1 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_4 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_58 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_fill_2 FILLER_12_80 ();
 sg13g2_decap_4 FILLER_12_98 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_decap_4 FILLER_12_143 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_decap_8 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_183 ();
 sg13g2_decap_4 FILLER_12_192 ();
 sg13g2_fill_1 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_4 FILLER_12_210 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_fill_2 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_fill_2 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_fill_2 FILLER_12_353 ();
 sg13g2_fill_1 FILLER_12_355 ();
 sg13g2_fill_2 FILLER_12_361 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_decap_4 FILLER_12_369 ();
 sg13g2_fill_1 FILLER_12_373 ();
 sg13g2_decap_4 FILLER_12_382 ();
 sg13g2_fill_1 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_410 ();
 sg13g2_fill_1 FILLER_12_425 ();
 sg13g2_decap_8 FILLER_12_453 ();
 sg13g2_decap_4 FILLER_12_460 ();
 sg13g2_decap_8 FILLER_12_468 ();
 sg13g2_decap_8 FILLER_12_475 ();
 sg13g2_fill_2 FILLER_12_482 ();
 sg13g2_fill_1 FILLER_12_484 ();
 sg13g2_decap_4 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_502 ();
 sg13g2_decap_8 FILLER_12_509 ();
 sg13g2_decap_4 FILLER_12_516 ();
 sg13g2_fill_1 FILLER_12_520 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_fill_2 FILLER_12_532 ();
 sg13g2_fill_1 FILLER_12_534 ();
 sg13g2_decap_4 FILLER_12_541 ();
 sg13g2_decap_8 FILLER_12_549 ();
 sg13g2_fill_1 FILLER_12_556 ();
 sg13g2_decap_8 FILLER_12_565 ();
 sg13g2_decap_8 FILLER_12_572 ();
 sg13g2_decap_8 FILLER_12_579 ();
 sg13g2_fill_1 FILLER_12_586 ();
 sg13g2_decap_8 FILLER_12_592 ();
 sg13g2_fill_1 FILLER_12_599 ();
 sg13g2_fill_1 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_4 FILLER_12_637 ();
 sg13g2_fill_1 FILLER_12_647 ();
 sg13g2_decap_8 FILLER_12_654 ();
 sg13g2_fill_2 FILLER_12_661 ();
 sg13g2_decap_8 FILLER_12_667 ();
 sg13g2_fill_2 FILLER_12_674 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_fill_1 FILLER_12_691 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_4 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_4 FILLER_13_67 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_decap_8 FILLER_13_83 ();
 sg13g2_decap_8 FILLER_13_90 ();
 sg13g2_decap_8 FILLER_13_97 ();
 sg13g2_decap_8 FILLER_13_104 ();
 sg13g2_decap_8 FILLER_13_111 ();
 sg13g2_decap_8 FILLER_13_118 ();
 sg13g2_decap_4 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_129 ();
 sg13g2_decap_8 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_fill_2 FILLER_13_151 ();
 sg13g2_decap_4 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_decap_4 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_fill_2 FILLER_13_196 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_decap_8 FILLER_13_205 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_decap_4 FILLER_13_219 ();
 sg13g2_decap_4 FILLER_13_242 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_fill_2 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_298 ();
 sg13g2_fill_2 FILLER_13_307 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_4 FILLER_13_354 ();
 sg13g2_fill_2 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_fill_2 FILLER_13_400 ();
 sg13g2_fill_1 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_8 FILLER_13_430 ();
 sg13g2_decap_4 FILLER_13_437 ();
 sg13g2_fill_2 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_451 ();
 sg13g2_fill_2 FILLER_13_458 ();
 sg13g2_fill_1 FILLER_13_460 ();
 sg13g2_fill_2 FILLER_13_479 ();
 sg13g2_fill_1 FILLER_13_481 ();
 sg13g2_fill_2 FILLER_13_487 ();
 sg13g2_decap_8 FILLER_13_505 ();
 sg13g2_decap_4 FILLER_13_512 ();
 sg13g2_fill_1 FILLER_13_516 ();
 sg13g2_fill_2 FILLER_13_528 ();
 sg13g2_fill_1 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_555 ();
 sg13g2_decap_8 FILLER_13_562 ();
 sg13g2_decap_4 FILLER_13_569 ();
 sg13g2_fill_1 FILLER_13_573 ();
 sg13g2_decap_8 FILLER_13_605 ();
 sg13g2_decap_8 FILLER_13_612 ();
 sg13g2_fill_2 FILLER_13_619 ();
 sg13g2_fill_1 FILLER_13_621 ();
 sg13g2_decap_8 FILLER_13_627 ();
 sg13g2_fill_1 FILLER_13_634 ();
 sg13g2_fill_2 FILLER_13_647 ();
 sg13g2_fill_1 FILLER_13_649 ();
 sg13g2_decap_4 FILLER_13_658 ();
 sg13g2_fill_2 FILLER_13_662 ();
 sg13g2_fill_2 FILLER_13_670 ();
 sg13g2_fill_1 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_712 ();
 sg13g2_decap_8 FILLER_13_719 ();
 sg13g2_fill_2 FILLER_13_726 ();
 sg13g2_decap_8 FILLER_13_736 ();
 sg13g2_decap_8 FILLER_13_743 ();
 sg13g2_decap_8 FILLER_13_750 ();
 sg13g2_decap_8 FILLER_13_757 ();
 sg13g2_decap_8 FILLER_13_764 ();
 sg13g2_decap_8 FILLER_13_771 ();
 sg13g2_decap_8 FILLER_13_778 ();
 sg13g2_decap_8 FILLER_13_785 ();
 sg13g2_decap_8 FILLER_13_792 ();
 sg13g2_decap_8 FILLER_13_799 ();
 sg13g2_decap_8 FILLER_13_806 ();
 sg13g2_decap_8 FILLER_13_813 ();
 sg13g2_decap_8 FILLER_13_820 ();
 sg13g2_decap_8 FILLER_13_827 ();
 sg13g2_decap_8 FILLER_13_834 ();
 sg13g2_decap_8 FILLER_13_841 ();
 sg13g2_decap_8 FILLER_13_848 ();
 sg13g2_decap_8 FILLER_13_855 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_40 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_decap_8 FILLER_14_54 ();
 sg13g2_decap_4 FILLER_14_61 ();
 sg13g2_fill_1 FILLER_14_65 ();
 sg13g2_decap_4 FILLER_14_78 ();
 sg13g2_decap_4 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_fill_2 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_125 ();
 sg13g2_decap_8 FILLER_14_146 ();
 sg13g2_fill_2 FILLER_14_153 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_fill_2 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_fill_1 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_4 FILLER_14_217 ();
 sg13g2_fill_2 FILLER_14_221 ();
 sg13g2_decap_4 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_231 ();
 sg13g2_decap_4 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_fill_2 FILLER_14_268 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_4 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_371 ();
 sg13g2_fill_1 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_fill_2 FILLER_14_387 ();
 sg13g2_decap_4 FILLER_14_398 ();
 sg13g2_fill_1 FILLER_14_407 ();
 sg13g2_decap_4 FILLER_14_414 ();
 sg13g2_fill_2 FILLER_14_423 ();
 sg13g2_decap_4 FILLER_14_439 ();
 sg13g2_decap_8 FILLER_14_457 ();
 sg13g2_fill_1 FILLER_14_464 ();
 sg13g2_decap_8 FILLER_14_471 ();
 sg13g2_decap_4 FILLER_14_478 ();
 sg13g2_fill_1 FILLER_14_482 ();
 sg13g2_decap_8 FILLER_14_487 ();
 sg13g2_fill_2 FILLER_14_494 ();
 sg13g2_fill_1 FILLER_14_496 ();
 sg13g2_decap_4 FILLER_14_508 ();
 sg13g2_fill_1 FILLER_14_512 ();
 sg13g2_decap_4 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_527 ();
 sg13g2_decap_8 FILLER_14_534 ();
 sg13g2_decap_4 FILLER_14_541 ();
 sg13g2_fill_2 FILLER_14_545 ();
 sg13g2_decap_4 FILLER_14_559 ();
 sg13g2_fill_2 FILLER_14_563 ();
 sg13g2_fill_2 FILLER_14_587 ();
 sg13g2_decap_8 FILLER_14_594 ();
 sg13g2_decap_8 FILLER_14_601 ();
 sg13g2_decap_4 FILLER_14_608 ();
 sg13g2_fill_1 FILLER_14_612 ();
 sg13g2_decap_4 FILLER_14_627 ();
 sg13g2_decap_8 FILLER_14_639 ();
 sg13g2_decap_8 FILLER_14_646 ();
 sg13g2_fill_2 FILLER_14_653 ();
 sg13g2_decap_4 FILLER_14_663 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_fill_2 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_fill_1 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_712 ();
 sg13g2_decap_4 FILLER_14_719 ();
 sg13g2_fill_2 FILLER_14_723 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_fill_1 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_835 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_8 FILLER_14_849 ();
 sg13g2_decap_4 FILLER_14_856 ();
 sg13g2_fill_2 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_44 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_51 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_decap_4 FILLER_15_64 ();
 sg13g2_fill_2 FILLER_15_68 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_fill_2 FILLER_15_134 ();
 sg13g2_decap_4 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_decap_8 FILLER_15_198 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_256 ();
 sg13g2_fill_1 FILLER_15_258 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_decap_4 FILLER_15_309 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_fill_2 FILLER_15_364 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_fill_1 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_fill_1 FILLER_15_397 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_fill_1 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_fill_2 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_479 ();
 sg13g2_fill_2 FILLER_15_486 ();
 sg13g2_decap_4 FILLER_15_496 ();
 sg13g2_fill_2 FILLER_15_505 ();
 sg13g2_decap_8 FILLER_15_513 ();
 sg13g2_fill_1 FILLER_15_520 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_fill_2 FILLER_15_550 ();
 sg13g2_fill_1 FILLER_15_552 ();
 sg13g2_fill_1 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_566 ();
 sg13g2_decap_4 FILLER_15_573 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_4 FILLER_15_588 ();
 sg13g2_fill_2 FILLER_15_592 ();
 sg13g2_decap_4 FILLER_15_600 ();
 sg13g2_fill_2 FILLER_15_604 ();
 sg13g2_fill_1 FILLER_15_611 ();
 sg13g2_decap_8 FILLER_15_618 ();
 sg13g2_decap_8 FILLER_15_625 ();
 sg13g2_decap_8 FILLER_15_632 ();
 sg13g2_fill_2 FILLER_15_639 ();
 sg13g2_fill_1 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_652 ();
 sg13g2_fill_1 FILLER_15_659 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_fill_2 FILLER_15_676 ();
 sg13g2_fill_1 FILLER_15_678 ();
 sg13g2_fill_2 FILLER_15_691 ();
 sg13g2_fill_1 FILLER_15_693 ();
 sg13g2_fill_1 FILLER_15_709 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_decap_8 FILLER_15_753 ();
 sg13g2_decap_8 FILLER_15_760 ();
 sg13g2_decap_4 FILLER_15_767 ();
 sg13g2_fill_2 FILLER_15_771 ();
 sg13g2_decap_8 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_8 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_816 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_4 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_18 ();
 sg13g2_decap_4 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_fill_2 FILLER_16_37 ();
 sg13g2_decap_4 FILLER_16_50 ();
 sg13g2_fill_2 FILLER_16_54 ();
 sg13g2_decap_4 FILLER_16_68 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_decap_8 FILLER_16_86 ();
 sg13g2_decap_8 FILLER_16_93 ();
 sg13g2_decap_8 FILLER_16_100 ();
 sg13g2_decap_8 FILLER_16_107 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_fill_2 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_128 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_fill_1 FILLER_16_137 ();
 sg13g2_decap_4 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_162 ();
 sg13g2_decap_4 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_decap_4 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_208 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_4 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_333 ();
 sg13g2_fill_2 FILLER_16_352 ();
 sg13g2_fill_1 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_fill_2 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_431 ();
 sg13g2_fill_1 FILLER_16_433 ();
 sg13g2_decap_4 FILLER_16_457 ();
 sg13g2_fill_1 FILLER_16_461 ();
 sg13g2_decap_8 FILLER_16_472 ();
 sg13g2_decap_4 FILLER_16_479 ();
 sg13g2_fill_2 FILLER_16_489 ();
 sg13g2_fill_1 FILLER_16_491 ();
 sg13g2_decap_8 FILLER_16_508 ();
 sg13g2_decap_4 FILLER_16_515 ();
 sg13g2_fill_1 FILLER_16_519 ();
 sg13g2_fill_2 FILLER_16_526 ();
 sg13g2_fill_1 FILLER_16_528 ();
 sg13g2_fill_2 FILLER_16_541 ();
 sg13g2_fill_1 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_550 ();
 sg13g2_fill_1 FILLER_16_557 ();
 sg13g2_fill_2 FILLER_16_576 ();
 sg13g2_fill_2 FILLER_16_583 ();
 sg13g2_fill_1 FILLER_16_585 ();
 sg13g2_decap_8 FILLER_16_607 ();
 sg13g2_decap_8 FILLER_16_614 ();
 sg13g2_decap_4 FILLER_16_621 ();
 sg13g2_fill_2 FILLER_16_625 ();
 sg13g2_fill_1 FILLER_16_640 ();
 sg13g2_fill_2 FILLER_16_656 ();
 sg13g2_decap_4 FILLER_16_672 ();
 sg13g2_fill_1 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_696 ();
 sg13g2_decap_4 FILLER_16_703 ();
 sg13g2_fill_1 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_713 ();
 sg13g2_decap_8 FILLER_16_720 ();
 sg13g2_decap_8 FILLER_16_727 ();
 sg13g2_decap_4 FILLER_16_734 ();
 sg13g2_fill_2 FILLER_16_738 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_fill_2 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_797 ();
 sg13g2_decap_8 FILLER_16_804 ();
 sg13g2_decap_8 FILLER_16_811 ();
 sg13g2_decap_8 FILLER_16_818 ();
 sg13g2_decap_8 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_832 ();
 sg13g2_decap_8 FILLER_16_839 ();
 sg13g2_decap_8 FILLER_16_846 ();
 sg13g2_decap_8 FILLER_16_853 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_22 ();
 sg13g2_decap_8 FILLER_17_29 ();
 sg13g2_decap_8 FILLER_17_36 ();
 sg13g2_decap_8 FILLER_17_43 ();
 sg13g2_decap_8 FILLER_17_50 ();
 sg13g2_decap_8 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_79 ();
 sg13g2_decap_4 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_100 ();
 sg13g2_decap_8 FILLER_17_107 ();
 sg13g2_fill_2 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_122 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_158 ();
 sg13g2_fill_2 FILLER_17_165 ();
 sg13g2_fill_1 FILLER_17_167 ();
 sg13g2_fill_2 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_194 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_4 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_fill_1 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_fill_1 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_4 FILLER_17_365 ();
 sg13g2_fill_1 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_392 ();
 sg13g2_decap_4 FILLER_17_431 ();
 sg13g2_fill_2 FILLER_17_435 ();
 sg13g2_fill_2 FILLER_17_443 ();
 sg13g2_fill_2 FILLER_17_456 ();
 sg13g2_fill_1 FILLER_17_458 ();
 sg13g2_fill_2 FILLER_17_474 ();
 sg13g2_decap_8 FILLER_17_492 ();
 sg13g2_decap_8 FILLER_17_499 ();
 sg13g2_decap_4 FILLER_17_506 ();
 sg13g2_decap_8 FILLER_17_521 ();
 sg13g2_decap_8 FILLER_17_528 ();
 sg13g2_fill_1 FILLER_17_540 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_4 FILLER_17_572 ();
 sg13g2_decap_4 FILLER_17_584 ();
 sg13g2_fill_2 FILLER_17_588 ();
 sg13g2_decap_4 FILLER_17_604 ();
 sg13g2_fill_1 FILLER_17_608 ();
 sg13g2_fill_1 FILLER_17_617 ();
 sg13g2_decap_8 FILLER_17_636 ();
 sg13g2_decap_8 FILLER_17_643 ();
 sg13g2_decap_8 FILLER_17_650 ();
 sg13g2_decap_8 FILLER_17_657 ();
 sg13g2_fill_2 FILLER_17_664 ();
 sg13g2_fill_1 FILLER_17_666 ();
 sg13g2_decap_8 FILLER_17_674 ();
 sg13g2_decap_4 FILLER_17_681 ();
 sg13g2_fill_1 FILLER_17_685 ();
 sg13g2_decap_8 FILLER_17_691 ();
 sg13g2_fill_1 FILLER_17_703 ();
 sg13g2_fill_2 FILLER_17_711 ();
 sg13g2_fill_1 FILLER_17_713 ();
 sg13g2_decap_8 FILLER_17_719 ();
 sg13g2_fill_2 FILLER_17_726 ();
 sg13g2_fill_1 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_737 ();
 sg13g2_fill_2 FILLER_17_747 ();
 sg13g2_fill_1 FILLER_17_749 ();
 sg13g2_fill_2 FILLER_17_765 ();
 sg13g2_fill_1 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_773 ();
 sg13g2_decap_8 FILLER_17_780 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_decap_8 FILLER_17_794 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_decap_8 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_decap_8 FILLER_17_836 ();
 sg13g2_decap_8 FILLER_17_843 ();
 sg13g2_decap_8 FILLER_17_850 ();
 sg13g2_decap_4 FILLER_17_857 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_23 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_fill_2 FILLER_18_73 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_decap_8 FILLER_18_89 ();
 sg13g2_decap_4 FILLER_18_96 ();
 sg13g2_decap_4 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_decap_4 FILLER_18_129 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_decap_4 FILLER_18_145 ();
 sg13g2_decap_8 FILLER_18_159 ();
 sg13g2_decap_4 FILLER_18_166 ();
 sg13g2_fill_2 FILLER_18_170 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_4 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_282 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_4 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_fill_2 FILLER_18_402 ();
 sg13g2_fill_1 FILLER_18_404 ();
 sg13g2_decap_8 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_8 FILLER_18_425 ();
 sg13g2_decap_8 FILLER_18_432 ();
 sg13g2_decap_8 FILLER_18_439 ();
 sg13g2_decap_8 FILLER_18_446 ();
 sg13g2_decap_8 FILLER_18_453 ();
 sg13g2_decap_8 FILLER_18_460 ();
 sg13g2_fill_1 FILLER_18_478 ();
 sg13g2_decap_8 FILLER_18_485 ();
 sg13g2_decap_8 FILLER_18_492 ();
 sg13g2_fill_2 FILLER_18_508 ();
 sg13g2_fill_1 FILLER_18_510 ();
 sg13g2_decap_8 FILLER_18_527 ();
 sg13g2_decap_4 FILLER_18_565 ();
 sg13g2_fill_1 FILLER_18_569 ();
 sg13g2_decap_4 FILLER_18_576 ();
 sg13g2_decap_8 FILLER_18_586 ();
 sg13g2_fill_1 FILLER_18_593 ();
 sg13g2_decap_8 FILLER_18_600 ();
 sg13g2_decap_8 FILLER_18_607 ();
 sg13g2_decap_4 FILLER_18_614 ();
 sg13g2_fill_2 FILLER_18_618 ();
 sg13g2_decap_4 FILLER_18_634 ();
 sg13g2_fill_2 FILLER_18_638 ();
 sg13g2_fill_2 FILLER_18_657 ();
 sg13g2_decap_8 FILLER_18_676 ();
 sg13g2_fill_2 FILLER_18_683 ();
 sg13g2_fill_1 FILLER_18_685 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_fill_1 FILLER_18_710 ();
 sg13g2_fill_2 FILLER_18_717 ();
 sg13g2_fill_1 FILLER_18_736 ();
 sg13g2_decap_8 FILLER_18_755 ();
 sg13g2_decap_4 FILLER_18_778 ();
 sg13g2_fill_1 FILLER_18_782 ();
 sg13g2_decap_4 FILLER_18_789 ();
 sg13g2_fill_2 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_18_849 ();
 sg13g2_decap_4 FILLER_18_856 ();
 sg13g2_fill_2 FILLER_18_860 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_fill_1 FILLER_19_48 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_decap_8 FILLER_19_66 ();
 sg13g2_decap_8 FILLER_19_85 ();
 sg13g2_decap_4 FILLER_19_92 ();
 sg13g2_decap_8 FILLER_19_107 ();
 sg13g2_decap_4 FILLER_19_114 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_decap_4 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_decap_4 FILLER_19_150 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_decap_4 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_184 ();
 sg13g2_decap_4 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_decap_8 FILLER_19_278 ();
 sg13g2_decap_4 FILLER_19_296 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_decap_4 FILLER_19_327 ();
 sg13g2_fill_2 FILLER_19_331 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_decap_4 FILLER_19_349 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_decap_4 FILLER_19_365 ();
 sg13g2_decap_4 FILLER_19_380 ();
 sg13g2_fill_2 FILLER_19_384 ();
 sg13g2_fill_2 FILLER_19_391 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_decap_4 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_19_451 ();
 sg13g2_fill_2 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_468 ();
 sg13g2_decap_4 FILLER_19_475 ();
 sg13g2_decap_8 FILLER_19_485 ();
 sg13g2_decap_8 FILLER_19_492 ();
 sg13g2_fill_2 FILLER_19_499 ();
 sg13g2_fill_1 FILLER_19_501 ();
 sg13g2_decap_8 FILLER_19_513 ();
 sg13g2_fill_1 FILLER_19_520 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_fill_1 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_548 ();
 sg13g2_decap_8 FILLER_19_565 ();
 sg13g2_decap_4 FILLER_19_572 ();
 sg13g2_decap_4 FILLER_19_594 ();
 sg13g2_fill_2 FILLER_19_603 ();
 sg13g2_fill_1 FILLER_19_605 ();
 sg13g2_decap_8 FILLER_19_611 ();
 sg13g2_decap_8 FILLER_19_618 ();
 sg13g2_fill_1 FILLER_19_625 ();
 sg13g2_decap_4 FILLER_19_631 ();
 sg13g2_fill_1 FILLER_19_635 ();
 sg13g2_fill_1 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_4 FILLER_19_676 ();
 sg13g2_decap_8 FILLER_19_696 ();
 sg13g2_fill_1 FILLER_19_703 ();
 sg13g2_decap_4 FILLER_19_709 ();
 sg13g2_fill_2 FILLER_19_713 ();
 sg13g2_decap_8 FILLER_19_720 ();
 sg13g2_fill_1 FILLER_19_727 ();
 sg13g2_decap_8 FILLER_19_748 ();
 sg13g2_fill_2 FILLER_19_755 ();
 sg13g2_fill_1 FILLER_19_766 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_4 FILLER_19_784 ();
 sg13g2_fill_1 FILLER_19_788 ();
 sg13g2_decap_8 FILLER_19_807 ();
 sg13g2_decap_4 FILLER_19_814 ();
 sg13g2_fill_2 FILLER_19_818 ();
 sg13g2_decap_8 FILLER_19_828 ();
 sg13g2_decap_8 FILLER_19_835 ();
 sg13g2_decap_8 FILLER_19_842 ();
 sg13g2_decap_8 FILLER_19_849 ();
 sg13g2_decap_4 FILLER_19_856 ();
 sg13g2_fill_2 FILLER_19_860 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_24 ();
 sg13g2_fill_1 FILLER_20_31 ();
 sg13g2_decap_8 FILLER_20_59 ();
 sg13g2_fill_1 FILLER_20_76 ();
 sg13g2_decap_8 FILLER_20_87 ();
 sg13g2_fill_2 FILLER_20_94 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_decap_4 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_decap_4 FILLER_20_158 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_decap_4 FILLER_20_187 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_decap_4 FILLER_20_198 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_decap_4 FILLER_20_237 ();
 sg13g2_decap_4 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_273 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_293 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_341 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_decap_4 FILLER_20_396 ();
 sg13g2_fill_2 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_decap_8 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_20_446 ();
 sg13g2_fill_2 FILLER_20_453 ();
 sg13g2_decap_4 FILLER_20_461 ();
 sg13g2_fill_2 FILLER_20_478 ();
 sg13g2_fill_1 FILLER_20_500 ();
 sg13g2_decap_8 FILLER_20_506 ();
 sg13g2_fill_2 FILLER_20_513 ();
 sg13g2_fill_2 FILLER_20_521 ();
 sg13g2_fill_1 FILLER_20_523 ();
 sg13g2_decap_8 FILLER_20_538 ();
 sg13g2_decap_8 FILLER_20_545 ();
 sg13g2_decap_4 FILLER_20_552 ();
 sg13g2_fill_2 FILLER_20_556 ();
 sg13g2_decap_8 FILLER_20_563 ();
 sg13g2_decap_4 FILLER_20_570 ();
 sg13g2_fill_2 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_fill_2 FILLER_20_588 ();
 sg13g2_fill_1 FILLER_20_590 ();
 sg13g2_fill_2 FILLER_20_615 ();
 sg13g2_fill_1 FILLER_20_617 ();
 sg13g2_fill_2 FILLER_20_636 ();
 sg13g2_fill_1 FILLER_20_638 ();
 sg13g2_fill_2 FILLER_20_653 ();
 sg13g2_decap_8 FILLER_20_661 ();
 sg13g2_decap_4 FILLER_20_668 ();
 sg13g2_fill_1 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_687 ();
 sg13g2_decap_8 FILLER_20_694 ();
 sg13g2_fill_2 FILLER_20_701 ();
 sg13g2_fill_1 FILLER_20_708 ();
 sg13g2_decap_4 FILLER_20_721 ();
 sg13g2_fill_2 FILLER_20_725 ();
 sg13g2_decap_4 FILLER_20_733 ();
 sg13g2_fill_1 FILLER_20_737 ();
 sg13g2_decap_8 FILLER_20_747 ();
 sg13g2_fill_1 FILLER_20_754 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_decap_8 FILLER_20_785 ();
 sg13g2_decap_4 FILLER_20_792 ();
 sg13g2_fill_1 FILLER_20_796 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_30 ();
 sg13g2_decap_4 FILLER_21_37 ();
 sg13g2_decap_4 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_4 FILLER_21_67 ();
 sg13g2_decap_4 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_86 ();
 sg13g2_decap_8 FILLER_21_96 ();
 sg13g2_decap_4 FILLER_21_103 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_decap_4 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_fill_2 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_4 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_353 ();
 sg13g2_decap_4 FILLER_21_367 ();
 sg13g2_fill_1 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_4 FILLER_21_395 ();
 sg13g2_decap_4 FILLER_21_417 ();
 sg13g2_fill_1 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_21_443 ();
 sg13g2_decap_4 FILLER_21_450 ();
 sg13g2_fill_1 FILLER_21_454 ();
 sg13g2_decap_4 FILLER_21_460 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_4 FILLER_21_483 ();
 sg13g2_fill_1 FILLER_21_498 ();
 sg13g2_decap_8 FILLER_21_507 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_decap_4 FILLER_21_521 ();
 sg13g2_decap_4 FILLER_21_538 ();
 sg13g2_decap_4 FILLER_21_550 ();
 sg13g2_fill_2 FILLER_21_571 ();
 sg13g2_fill_1 FILLER_21_573 ();
 sg13g2_decap_8 FILLER_21_586 ();
 sg13g2_fill_1 FILLER_21_593 ();
 sg13g2_fill_1 FILLER_21_599 ();
 sg13g2_decap_8 FILLER_21_624 ();
 sg13g2_decap_8 FILLER_21_631 ();
 sg13g2_decap_8 FILLER_21_638 ();
 sg13g2_decap_8 FILLER_21_645 ();
 sg13g2_decap_4 FILLER_21_652 ();
 sg13g2_fill_2 FILLER_21_656 ();
 sg13g2_decap_8 FILLER_21_666 ();
 sg13g2_fill_1 FILLER_21_673 ();
 sg13g2_fill_1 FILLER_21_680 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_fill_1 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_716 ();
 sg13g2_decap_8 FILLER_21_723 ();
 sg13g2_decap_8 FILLER_21_730 ();
 sg13g2_decap_4 FILLER_21_737 ();
 sg13g2_decap_8 FILLER_21_755 ();
 sg13g2_decap_8 FILLER_21_762 ();
 sg13g2_fill_2 FILLER_21_769 ();
 sg13g2_decap_8 FILLER_21_792 ();
 sg13g2_decap_8 FILLER_21_799 ();
 sg13g2_fill_2 FILLER_21_812 ();
 sg13g2_fill_1 FILLER_21_814 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_decap_8 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_850 ();
 sg13g2_decap_4 FILLER_21_857 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_11 ();
 sg13g2_fill_1 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_45 ();
 sg13g2_fill_1 FILLER_22_47 ();
 sg13g2_decap_8 FILLER_22_52 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_fill_2 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_1 FILLER_22_147 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_174 ();
 sg13g2_decap_8 FILLER_22_181 ();
 sg13g2_decap_4 FILLER_22_188 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_208 ();
 sg13g2_decap_4 FILLER_22_216 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_271 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_370 ();
 sg13g2_fill_1 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_fill_2 FILLER_22_424 ();
 sg13g2_decap_8 FILLER_22_439 ();
 sg13g2_decap_8 FILLER_22_446 ();
 sg13g2_decap_4 FILLER_22_453 ();
 sg13g2_fill_2 FILLER_22_468 ();
 sg13g2_fill_1 FILLER_22_470 ();
 sg13g2_decap_4 FILLER_22_484 ();
 sg13g2_fill_2 FILLER_22_488 ();
 sg13g2_decap_8 FILLER_22_509 ();
 sg13g2_fill_1 FILLER_22_516 ();
 sg13g2_decap_8 FILLER_22_523 ();
 sg13g2_fill_2 FILLER_22_534 ();
 sg13g2_decap_8 FILLER_22_544 ();
 sg13g2_decap_4 FILLER_22_551 ();
 sg13g2_fill_2 FILLER_22_555 ();
 sg13g2_decap_8 FILLER_22_571 ();
 sg13g2_fill_1 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_592 ();
 sg13g2_fill_1 FILLER_22_599 ();
 sg13g2_decap_4 FILLER_22_608 ();
 sg13g2_decap_8 FILLER_22_617 ();
 sg13g2_decap_4 FILLER_22_624 ();
 sg13g2_fill_2 FILLER_22_628 ();
 sg13g2_fill_2 FILLER_22_643 ();
 sg13g2_fill_1 FILLER_22_645 ();
 sg13g2_decap_4 FILLER_22_654 ();
 sg13g2_decap_4 FILLER_22_663 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_fill_1 FILLER_22_679 ();
 sg13g2_fill_2 FILLER_22_705 ();
 sg13g2_fill_1 FILLER_22_707 ();
 sg13g2_fill_2 FILLER_22_721 ();
 sg13g2_fill_1 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_743 ();
 sg13g2_fill_2 FILLER_22_750 ();
 sg13g2_fill_1 FILLER_22_752 ();
 sg13g2_decap_4 FILLER_22_762 ();
 sg13g2_fill_1 FILLER_22_766 ();
 sg13g2_decap_8 FILLER_22_771 ();
 sg13g2_decap_8 FILLER_22_778 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_820 ();
 sg13g2_fill_1 FILLER_22_827 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_57 ();
 sg13g2_decap_8 FILLER_23_64 ();
 sg13g2_fill_2 FILLER_23_75 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_87 ();
 sg13g2_decap_4 FILLER_23_94 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_4 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_145 ();
 sg13g2_decap_8 FILLER_23_152 ();
 sg13g2_decap_4 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_decap_4 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_213 ();
 sg13g2_decap_4 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_decap_4 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_decap_4 FILLER_23_308 ();
 sg13g2_fill_2 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_decap_4 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_416 ();
 sg13g2_fill_2 FILLER_23_423 ();
 sg13g2_fill_1 FILLER_23_425 ();
 sg13g2_fill_2 FILLER_23_431 ();
 sg13g2_fill_1 FILLER_23_433 ();
 sg13g2_decap_4 FILLER_23_442 ();
 sg13g2_fill_2 FILLER_23_446 ();
 sg13g2_fill_2 FILLER_23_465 ();
 sg13g2_fill_1 FILLER_23_467 ();
 sg13g2_decap_8 FILLER_23_478 ();
 sg13g2_decap_4 FILLER_23_485 ();
 sg13g2_decap_4 FILLER_23_494 ();
 sg13g2_fill_2 FILLER_23_502 ();
 sg13g2_fill_1 FILLER_23_504 ();
 sg13g2_decap_4 FILLER_23_513 ();
 sg13g2_fill_2 FILLER_23_517 ();
 sg13g2_fill_2 FILLER_23_524 ();
 sg13g2_fill_1 FILLER_23_526 ();
 sg13g2_fill_1 FILLER_23_533 ();
 sg13g2_fill_1 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_551 ();
 sg13g2_fill_1 FILLER_23_558 ();
 sg13g2_decap_8 FILLER_23_564 ();
 sg13g2_decap_4 FILLER_23_575 ();
 sg13g2_fill_1 FILLER_23_579 ();
 sg13g2_fill_2 FILLER_23_584 ();
 sg13g2_fill_1 FILLER_23_586 ();
 sg13g2_decap_8 FILLER_23_593 ();
 sg13g2_fill_1 FILLER_23_600 ();
 sg13g2_decap_8 FILLER_23_627 ();
 sg13g2_fill_2 FILLER_23_634 ();
 sg13g2_decap_4 FILLER_23_642 ();
 sg13g2_fill_2 FILLER_23_646 ();
 sg13g2_decap_4 FILLER_23_657 ();
 sg13g2_decap_8 FILLER_23_667 ();
 sg13g2_decap_4 FILLER_23_674 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_fill_1 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_713 ();
 sg13g2_decap_8 FILLER_23_720 ();
 sg13g2_fill_2 FILLER_23_727 ();
 sg13g2_decap_8 FILLER_23_740 ();
 sg13g2_decap_4 FILLER_23_747 ();
 sg13g2_fill_2 FILLER_23_751 ();
 sg13g2_fill_1 FILLER_23_757 ();
 sg13g2_decap_4 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_790 ();
 sg13g2_decap_8 FILLER_23_802 ();
 sg13g2_decap_4 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_821 ();
 sg13g2_decap_8 FILLER_23_828 ();
 sg13g2_decap_8 FILLER_23_835 ();
 sg13g2_decap_8 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_849 ();
 sg13g2_decap_4 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_32 ();
 sg13g2_decap_4 FILLER_24_54 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_89 ();
 sg13g2_decap_4 FILLER_24_96 ();
 sg13g2_decap_8 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_125 ();
 sg13g2_decap_8 FILLER_24_132 ();
 sg13g2_decap_4 FILLER_24_139 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_decap_4 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_decap_4 FILLER_24_192 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_decap_4 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_fill_2 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_24_425 ();
 sg13g2_decap_4 FILLER_24_439 ();
 sg13g2_fill_1 FILLER_24_443 ();
 sg13g2_decap_8 FILLER_24_454 ();
 sg13g2_decap_4 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_475 ();
 sg13g2_decap_8 FILLER_24_482 ();
 sg13g2_fill_1 FILLER_24_489 ();
 sg13g2_decap_8 FILLER_24_495 ();
 sg13g2_decap_8 FILLER_24_502 ();
 sg13g2_decap_8 FILLER_24_509 ();
 sg13g2_fill_2 FILLER_24_524 ();
 sg13g2_fill_1 FILLER_24_526 ();
 sg13g2_decap_8 FILLER_24_538 ();
 sg13g2_decap_8 FILLER_24_545 ();
 sg13g2_fill_2 FILLER_24_552 ();
 sg13g2_fill_1 FILLER_24_554 ();
 sg13g2_fill_1 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_573 ();
 sg13g2_decap_8 FILLER_24_601 ();
 sg13g2_decap_8 FILLER_24_608 ();
 sg13g2_fill_2 FILLER_24_615 ();
 sg13g2_decap_8 FILLER_24_632 ();
 sg13g2_decap_4 FILLER_24_639 ();
 sg13g2_fill_2 FILLER_24_643 ();
 sg13g2_decap_8 FILLER_24_657 ();
 sg13g2_fill_2 FILLER_24_675 ();
 sg13g2_decap_8 FILLER_24_692 ();
 sg13g2_fill_2 FILLER_24_699 ();
 sg13g2_decap_4 FILLER_24_726 ();
 sg13g2_fill_1 FILLER_24_730 ();
 sg13g2_fill_1 FILLER_24_736 ();
 sg13g2_decap_8 FILLER_24_750 ();
 sg13g2_fill_2 FILLER_24_757 ();
 sg13g2_fill_1 FILLER_24_759 ();
 sg13g2_decap_8 FILLER_24_769 ();
 sg13g2_decap_4 FILLER_24_776 ();
 sg13g2_fill_2 FILLER_24_780 ();
 sg13g2_decap_4 FILLER_24_787 ();
 sg13g2_fill_1 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_808 ();
 sg13g2_decap_4 FILLER_24_815 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_fill_1 FILLER_24_847 ();
 sg13g2_decap_4 FILLER_24_856 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_23 ();
 sg13g2_decap_8 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_46 ();
 sg13g2_decap_4 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_57 ();
 sg13g2_decap_8 FILLER_25_66 ();
 sg13g2_decap_8 FILLER_25_73 ();
 sg13g2_decap_4 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_89 ();
 sg13g2_decap_8 FILLER_25_96 ();
 sg13g2_decap_4 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_decap_4 FILLER_25_166 ();
 sg13g2_decap_4 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_4 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_4 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_decap_4 FILLER_25_346 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_4 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_398 ();
 sg13g2_fill_1 FILLER_25_400 ();
 sg13g2_decap_4 FILLER_25_407 ();
 sg13g2_fill_2 FILLER_25_411 ();
 sg13g2_fill_2 FILLER_25_421 ();
 sg13g2_fill_1 FILLER_25_423 ();
 sg13g2_decap_8 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_25_436 ();
 sg13g2_fill_2 FILLER_25_443 ();
 sg13g2_fill_2 FILLER_25_450 ();
 sg13g2_fill_1 FILLER_25_452 ();
 sg13g2_fill_2 FILLER_25_465 ();
 sg13g2_decap_8 FILLER_25_472 ();
 sg13g2_fill_1 FILLER_25_479 ();
 sg13g2_fill_2 FILLER_25_485 ();
 sg13g2_fill_1 FILLER_25_487 ();
 sg13g2_decap_8 FILLER_25_493 ();
 sg13g2_fill_1 FILLER_25_514 ();
 sg13g2_decap_4 FILLER_25_523 ();
 sg13g2_fill_1 FILLER_25_527 ();
 sg13g2_fill_2 FILLER_25_533 ();
 sg13g2_fill_1 FILLER_25_535 ();
 sg13g2_decap_8 FILLER_25_541 ();
 sg13g2_fill_2 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_576 ();
 sg13g2_fill_1 FILLER_25_583 ();
 sg13g2_decap_4 FILLER_25_593 ();
 sg13g2_fill_1 FILLER_25_597 ();
 sg13g2_decap_8 FILLER_25_607 ();
 sg13g2_fill_1 FILLER_25_614 ();
 sg13g2_decap_8 FILLER_25_620 ();
 sg13g2_fill_1 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_fill_1 FILLER_25_658 ();
 sg13g2_fill_1 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_684 ();
 sg13g2_fill_1 FILLER_25_691 ();
 sg13g2_decap_8 FILLER_25_704 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_4 FILLER_25_718 ();
 sg13g2_decap_8 FILLER_25_738 ();
 sg13g2_decap_8 FILLER_25_745 ();
 sg13g2_fill_1 FILLER_25_752 ();
 sg13g2_decap_8 FILLER_25_771 ();
 sg13g2_decap_8 FILLER_25_778 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_fill_2 FILLER_25_800 ();
 sg13g2_fill_1 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_fill_2 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_855 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_16 ();
 sg13g2_decap_4 FILLER_26_23 ();
 sg13g2_fill_1 FILLER_26_27 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_2 FILLER_26_45 ();
 sg13g2_decap_8 FILLER_26_58 ();
 sg13g2_fill_1 FILLER_26_75 ();
 sg13g2_fill_2 FILLER_26_86 ();
 sg13g2_decap_8 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_decap_8 FILLER_26_141 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_decap_4 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_4 FILLER_26_186 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_257 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_fill_1 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_338 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_4 FILLER_26_384 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_4 FILLER_26_420 ();
 sg13g2_fill_1 FILLER_26_424 ();
 sg13g2_decap_8 FILLER_26_444 ();
 sg13g2_decap_8 FILLER_26_451 ();
 sg13g2_decap_8 FILLER_26_458 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_4 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_498 ();
 sg13g2_decap_8 FILLER_26_505 ();
 sg13g2_decap_4 FILLER_26_512 ();
 sg13g2_decap_8 FILLER_26_538 ();
 sg13g2_decap_8 FILLER_26_545 ();
 sg13g2_decap_4 FILLER_26_552 ();
 sg13g2_fill_2 FILLER_26_556 ();
 sg13g2_decap_8 FILLER_26_566 ();
 sg13g2_decap_8 FILLER_26_573 ();
 sg13g2_fill_2 FILLER_26_580 ();
 sg13g2_fill_1 FILLER_26_582 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_fill_2 FILLER_26_602 ();
 sg13g2_fill_1 FILLER_26_604 ();
 sg13g2_decap_8 FILLER_26_625 ();
 sg13g2_decap_8 FILLER_26_632 ();
 sg13g2_decap_8 FILLER_26_639 ();
 sg13g2_fill_1 FILLER_26_646 ();
 sg13g2_decap_8 FILLER_26_652 ();
 sg13g2_fill_2 FILLER_26_659 ();
 sg13g2_fill_1 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_678 ();
 sg13g2_fill_2 FILLER_26_685 ();
 sg13g2_fill_1 FILLER_26_687 ();
 sg13g2_fill_1 FILLER_26_701 ();
 sg13g2_decap_8 FILLER_26_710 ();
 sg13g2_fill_2 FILLER_26_717 ();
 sg13g2_decap_8 FILLER_26_724 ();
 sg13g2_fill_2 FILLER_26_731 ();
 sg13g2_decap_4 FILLER_26_738 ();
 sg13g2_fill_2 FILLER_26_742 ();
 sg13g2_fill_2 FILLER_26_753 ();
 sg13g2_fill_1 FILLER_26_755 ();
 sg13g2_decap_8 FILLER_26_767 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_4 FILLER_26_829 ();
 sg13g2_fill_2 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_843 ();
 sg13g2_decap_4 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_20 ();
 sg13g2_decap_4 FILLER_27_27 ();
 sg13g2_fill_1 FILLER_27_31 ();
 sg13g2_decap_8 FILLER_27_44 ();
 sg13g2_decap_8 FILLER_27_51 ();
 sg13g2_decap_8 FILLER_27_64 ();
 sg13g2_decap_4 FILLER_27_71 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_decap_8 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_decap_4 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_4 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_decap_4 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_fill_2 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_decap_4 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_348 ();
 sg13g2_decap_8 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_fill_2 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_4 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_8 FILLER_27_432 ();
 sg13g2_decap_8 FILLER_27_439 ();
 sg13g2_decap_4 FILLER_27_446 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_465 ();
 sg13g2_fill_1 FILLER_27_467 ();
 sg13g2_decap_8 FILLER_27_473 ();
 sg13g2_decap_4 FILLER_27_480 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_fill_1 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_517 ();
 sg13g2_decap_4 FILLER_27_524 ();
 sg13g2_fill_1 FILLER_27_528 ();
 sg13g2_fill_2 FILLER_27_539 ();
 sg13g2_fill_1 FILLER_27_541 ();
 sg13g2_decap_8 FILLER_27_547 ();
 sg13g2_decap_4 FILLER_27_570 ();
 sg13g2_fill_2 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_600 ();
 sg13g2_fill_1 FILLER_27_607 ();
 sg13g2_decap_4 FILLER_27_614 ();
 sg13g2_fill_1 FILLER_27_646 ();
 sg13g2_decap_8 FILLER_27_656 ();
 sg13g2_decap_8 FILLER_27_663 ();
 sg13g2_fill_2 FILLER_27_670 ();
 sg13g2_fill_1 FILLER_27_677 ();
 sg13g2_fill_2 FILLER_27_682 ();
 sg13g2_decap_4 FILLER_27_692 ();
 sg13g2_fill_1 FILLER_27_696 ();
 sg13g2_decap_4 FILLER_27_702 ();
 sg13g2_fill_2 FILLER_27_706 ();
 sg13g2_decap_8 FILLER_27_713 ();
 sg13g2_decap_8 FILLER_27_720 ();
 sg13g2_decap_4 FILLER_27_727 ();
 sg13g2_fill_1 FILLER_27_731 ();
 sg13g2_decap_8 FILLER_27_744 ();
 sg13g2_decap_8 FILLER_27_751 ();
 sg13g2_decap_8 FILLER_27_758 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_fill_1 FILLER_27_778 ();
 sg13g2_fill_2 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_4 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_fill_1 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_832 ();
 sg13g2_decap_4 FILLER_27_839 ();
 sg13g2_fill_2 FILLER_27_843 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_4 FILLER_27_858 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_decap_4 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_71 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_84 ();
 sg13g2_decap_4 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_113 ();
 sg13g2_decap_8 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_decap_4 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_229 ();
 sg13g2_decap_4 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_decap_8 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_4 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_324 ();
 sg13g2_decap_4 FILLER_28_331 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_fill_1 FILLER_28_394 ();
 sg13g2_fill_1 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_fill_1 FILLER_28_430 ();
 sg13g2_fill_2 FILLER_28_444 ();
 sg13g2_decap_4 FILLER_28_455 ();
 sg13g2_fill_2 FILLER_28_459 ();
 sg13g2_fill_2 FILLER_28_485 ();
 sg13g2_fill_1 FILLER_28_493 ();
 sg13g2_decap_8 FILLER_28_502 ();
 sg13g2_decap_8 FILLER_28_509 ();
 sg13g2_decap_4 FILLER_28_516 ();
 sg13g2_fill_1 FILLER_28_520 ();
 sg13g2_fill_1 FILLER_28_526 ();
 sg13g2_decap_4 FILLER_28_535 ();
 sg13g2_decap_8 FILLER_28_547 ();
 sg13g2_fill_2 FILLER_28_554 ();
 sg13g2_fill_1 FILLER_28_556 ();
 sg13g2_fill_1 FILLER_28_561 ();
 sg13g2_decap_8 FILLER_28_566 ();
 sg13g2_decap_8 FILLER_28_573 ();
 sg13g2_decap_4 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_599 ();
 sg13g2_decap_4 FILLER_28_606 ();
 sg13g2_fill_2 FILLER_28_610 ();
 sg13g2_fill_2 FILLER_28_616 ();
 sg13g2_fill_1 FILLER_28_618 ();
 sg13g2_decap_8 FILLER_28_624 ();
 sg13g2_decap_4 FILLER_28_631 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_4 FILLER_28_650 ();
 sg13g2_fill_1 FILLER_28_654 ();
 sg13g2_decap_8 FILLER_28_671 ();
 sg13g2_fill_2 FILLER_28_678 ();
 sg13g2_fill_1 FILLER_28_680 ();
 sg13g2_decap_8 FILLER_28_691 ();
 sg13g2_decap_8 FILLER_28_698 ();
 sg13g2_decap_8 FILLER_28_705 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_4 FILLER_28_741 ();
 sg13g2_fill_2 FILLER_28_745 ();
 sg13g2_fill_2 FILLER_28_789 ();
 sg13g2_decap_8 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_806 ();
 sg13g2_fill_1 FILLER_28_813 ();
 sg13g2_fill_2 FILLER_28_823 ();
 sg13g2_fill_1 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_831 ();
 sg13g2_fill_2 FILLER_28_838 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_27 ();
 sg13g2_fill_2 FILLER_29_38 ();
 sg13g2_decap_4 FILLER_29_54 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_decap_4 FILLER_29_110 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_decap_4 FILLER_29_137 ();
 sg13g2_fill_2 FILLER_29_141 ();
 sg13g2_fill_2 FILLER_29_165 ();
 sg13g2_fill_1 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_197 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_2 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_decap_4 FILLER_29_246 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_decap_4 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_decap_4 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_378 ();
 sg13g2_decap_4 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_409 ();
 sg13g2_decap_8 FILLER_29_416 ();
 sg13g2_fill_2 FILLER_29_423 ();
 sg13g2_decap_4 FILLER_29_433 ();
 sg13g2_fill_2 FILLER_29_437 ();
 sg13g2_decap_8 FILLER_29_444 ();
 sg13g2_fill_2 FILLER_29_451 ();
 sg13g2_decap_8 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_466 ();
 sg13g2_decap_8 FILLER_29_478 ();
 sg13g2_fill_2 FILLER_29_485 ();
 sg13g2_decap_8 FILLER_29_493 ();
 sg13g2_decap_4 FILLER_29_504 ();
 sg13g2_fill_1 FILLER_29_508 ();
 sg13g2_decap_4 FILLER_29_515 ();
 sg13g2_fill_1 FILLER_29_519 ();
 sg13g2_decap_4 FILLER_29_525 ();
 sg13g2_fill_1 FILLER_29_529 ();
 sg13g2_decap_8 FILLER_29_535 ();
 sg13g2_fill_2 FILLER_29_542 ();
 sg13g2_decap_4 FILLER_29_552 ();
 sg13g2_fill_1 FILLER_29_556 ();
 sg13g2_decap_8 FILLER_29_570 ();
 sg13g2_fill_2 FILLER_29_577 ();
 sg13g2_decap_8 FILLER_29_596 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_4 FILLER_29_616 ();
 sg13g2_decap_4 FILLER_29_631 ();
 sg13g2_fill_1 FILLER_29_635 ();
 sg13g2_decap_8 FILLER_29_641 ();
 sg13g2_fill_1 FILLER_29_652 ();
 sg13g2_decap_4 FILLER_29_658 ();
 sg13g2_fill_2 FILLER_29_662 ();
 sg13g2_decap_4 FILLER_29_669 ();
 sg13g2_fill_1 FILLER_29_673 ();
 sg13g2_fill_2 FILLER_29_683 ();
 sg13g2_fill_1 FILLER_29_685 ();
 sg13g2_decap_8 FILLER_29_694 ();
 sg13g2_fill_1 FILLER_29_701 ();
 sg13g2_decap_4 FILLER_29_712 ();
 sg13g2_decap_8 FILLER_29_726 ();
 sg13g2_decap_4 FILLER_29_733 ();
 sg13g2_fill_2 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_fill_1 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_fill_2 FILLER_29_786 ();
 sg13g2_fill_1 FILLER_29_788 ();
 sg13g2_decap_4 FILLER_29_794 ();
 sg13g2_fill_2 FILLER_29_798 ();
 sg13g2_fill_2 FILLER_29_806 ();
 sg13g2_fill_1 FILLER_29_808 ();
 sg13g2_decap_8 FILLER_29_827 ();
 sg13g2_fill_2 FILLER_29_834 ();
 sg13g2_decap_8 FILLER_29_841 ();
 sg13g2_decap_8 FILLER_29_848 ();
 sg13g2_decap_8 FILLER_29_855 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_26 ();
 sg13g2_decap_4 FILLER_30_33 ();
 sg13g2_fill_1 FILLER_30_37 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_62 ();
 sg13g2_decap_8 FILLER_30_69 ();
 sg13g2_fill_2 FILLER_30_76 ();
 sg13g2_decap_8 FILLER_30_88 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_111 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_decap_8 FILLER_30_125 ();
 sg13g2_decap_8 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_decap_4 FILLER_30_146 ();
 sg13g2_decap_8 FILLER_30_166 ();
 sg13g2_decap_4 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_decap_8 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_239 ();
 sg13g2_decap_4 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_decap_8 FILLER_30_292 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_decap_4 FILLER_30_309 ();
 sg13g2_fill_2 FILLER_30_313 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_4 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_30_416 ();
 sg13g2_fill_1 FILLER_30_423 ();
 sg13g2_decap_4 FILLER_30_438 ();
 sg13g2_decap_8 FILLER_30_447 ();
 sg13g2_fill_2 FILLER_30_454 ();
 sg13g2_fill_1 FILLER_30_456 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_fill_2 FILLER_30_474 ();
 sg13g2_decap_4 FILLER_30_484 ();
 sg13g2_fill_1 FILLER_30_505 ();
 sg13g2_fill_1 FILLER_30_519 ();
 sg13g2_decap_8 FILLER_30_565 ();
 sg13g2_decap_8 FILLER_30_572 ();
 sg13g2_decap_4 FILLER_30_589 ();
 sg13g2_fill_2 FILLER_30_593 ();
 sg13g2_fill_1 FILLER_30_599 ();
 sg13g2_fill_2 FILLER_30_608 ();
 sg13g2_decap_8 FILLER_30_622 ();
 sg13g2_fill_1 FILLER_30_629 ();
 sg13g2_decap_4 FILLER_30_643 ();
 sg13g2_decap_4 FILLER_30_655 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_4 FILLER_30_679 ();
 sg13g2_fill_1 FILLER_30_683 ();
 sg13g2_decap_8 FILLER_30_695 ();
 sg13g2_decap_4 FILLER_30_702 ();
 sg13g2_fill_2 FILLER_30_706 ();
 sg13g2_fill_1 FILLER_30_713 ();
 sg13g2_decap_8 FILLER_30_722 ();
 sg13g2_fill_1 FILLER_30_729 ();
 sg13g2_fill_1 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_751 ();
 sg13g2_fill_2 FILLER_30_758 ();
 sg13g2_decap_4 FILLER_30_778 ();
 sg13g2_fill_2 FILLER_30_782 ();
 sg13g2_decap_4 FILLER_30_794 ();
 sg13g2_decap_4 FILLER_30_811 ();
 sg13g2_fill_2 FILLER_30_815 ();
 sg13g2_fill_1 FILLER_30_832 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_24 ();
 sg13g2_fill_2 FILLER_31_31 ();
 sg13g2_fill_1 FILLER_31_38 ();
 sg13g2_decap_8 FILLER_31_44 ();
 sg13g2_decap_4 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_fill_2 FILLER_31_60 ();
 sg13g2_decap_4 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_90 ();
 sg13g2_fill_1 FILLER_31_97 ();
 sg13g2_decap_8 FILLER_31_106 ();
 sg13g2_decap_8 FILLER_31_113 ();
 sg13g2_decap_8 FILLER_31_132 ();
 sg13g2_decap_8 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_decap_4 FILLER_31_247 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_273 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_4 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_418 ();
 sg13g2_decap_8 FILLER_31_433 ();
 sg13g2_decap_4 FILLER_31_440 ();
 sg13g2_fill_2 FILLER_31_444 ();
 sg13g2_fill_2 FILLER_31_463 ();
 sg13g2_fill_1 FILLER_31_465 ();
 sg13g2_decap_8 FILLER_31_485 ();
 sg13g2_decap_8 FILLER_31_492 ();
 sg13g2_decap_8 FILLER_31_499 ();
 sg13g2_decap_8 FILLER_31_506 ();
 sg13g2_decap_8 FILLER_31_513 ();
 sg13g2_decap_8 FILLER_31_520 ();
 sg13g2_decap_4 FILLER_31_527 ();
 sg13g2_decap_8 FILLER_31_536 ();
 sg13g2_decap_8 FILLER_31_543 ();
 sg13g2_decap_8 FILLER_31_550 ();
 sg13g2_fill_2 FILLER_31_557 ();
 sg13g2_decap_8 FILLER_31_582 ();
 sg13g2_decap_8 FILLER_31_589 ();
 sg13g2_decap_8 FILLER_31_596 ();
 sg13g2_decap_4 FILLER_31_603 ();
 sg13g2_fill_1 FILLER_31_607 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_fill_1 FILLER_31_629 ();
 sg13g2_decap_8 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_645 ();
 sg13g2_decap_8 FILLER_31_652 ();
 sg13g2_fill_2 FILLER_31_659 ();
 sg13g2_fill_2 FILLER_31_666 ();
 sg13g2_fill_2 FILLER_31_674 ();
 sg13g2_fill_1 FILLER_31_676 ();
 sg13g2_decap_4 FILLER_31_692 ();
 sg13g2_fill_2 FILLER_31_696 ();
 sg13g2_decap_4 FILLER_31_706 ();
 sg13g2_fill_2 FILLER_31_710 ();
 sg13g2_decap_8 FILLER_31_717 ();
 sg13g2_decap_8 FILLER_31_724 ();
 sg13g2_decap_4 FILLER_31_731 ();
 sg13g2_fill_2 FILLER_31_740 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_fill_1 FILLER_31_769 ();
 sg13g2_decap_8 FILLER_31_780 ();
 sg13g2_fill_2 FILLER_31_787 ();
 sg13g2_fill_1 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_fill_2 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_823 ();
 sg13g2_decap_8 FILLER_31_830 ();
 sg13g2_decap_4 FILLER_31_837 ();
 sg13g2_fill_1 FILLER_31_841 ();
 sg13g2_decap_8 FILLER_31_851 ();
 sg13g2_decap_4 FILLER_31_858 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_23 ();
 sg13g2_fill_1 FILLER_32_25 ();
 sg13g2_fill_2 FILLER_32_37 ();
 sg13g2_decap_8 FILLER_32_54 ();
 sg13g2_decap_4 FILLER_32_61 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_fill_2 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_82 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_95 ();
 sg13g2_decap_4 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_117 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_4 FILLER_32_185 ();
 sg13g2_decap_4 FILLER_32_210 ();
 sg13g2_decap_4 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_4 FILLER_32_284 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_1 FILLER_32_313 ();
 sg13g2_decap_8 FILLER_32_335 ();
 sg13g2_decap_4 FILLER_32_342 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_366 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_decap_4 FILLER_32_416 ();
 sg13g2_fill_2 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_430 ();
 sg13g2_fill_1 FILLER_32_432 ();
 sg13g2_decap_8 FILLER_32_438 ();
 sg13g2_decap_8 FILLER_32_445 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_fill_2 FILLER_32_478 ();
 sg13g2_fill_2 FILLER_32_486 ();
 sg13g2_fill_1 FILLER_32_488 ();
 sg13g2_decap_8 FILLER_32_516 ();
 sg13g2_fill_2 FILLER_32_523 ();
 sg13g2_fill_1 FILLER_32_525 ();
 sg13g2_decap_4 FILLER_32_540 ();
 sg13g2_fill_2 FILLER_32_544 ();
 sg13g2_decap_8 FILLER_32_559 ();
 sg13g2_decap_4 FILLER_32_566 ();
 sg13g2_fill_2 FILLER_32_570 ();
 sg13g2_fill_1 FILLER_32_591 ();
 sg13g2_decap_8 FILLER_32_601 ();
 sg13g2_decap_8 FILLER_32_608 ();
 sg13g2_fill_1 FILLER_32_615 ();
 sg13g2_decap_8 FILLER_32_628 ();
 sg13g2_fill_2 FILLER_32_635 ();
 sg13g2_fill_2 FILLER_32_657 ();
 sg13g2_decap_4 FILLER_32_664 ();
 sg13g2_fill_2 FILLER_32_668 ();
 sg13g2_decap_8 FILLER_32_675 ();
 sg13g2_fill_2 FILLER_32_682 ();
 sg13g2_fill_1 FILLER_32_684 ();
 sg13g2_decap_4 FILLER_32_696 ();
 sg13g2_fill_1 FILLER_32_700 ();
 sg13g2_fill_2 FILLER_32_736 ();
 sg13g2_decap_8 FILLER_32_750 ();
 sg13g2_fill_1 FILLER_32_757 ();
 sg13g2_fill_2 FILLER_32_764 ();
 sg13g2_fill_1 FILLER_32_766 ();
 sg13g2_fill_1 FILLER_32_775 ();
 sg13g2_decap_4 FILLER_32_792 ();
 sg13g2_decap_8 FILLER_32_809 ();
 sg13g2_fill_2 FILLER_32_816 ();
 sg13g2_fill_1 FILLER_32_818 ();
 sg13g2_fill_2 FILLER_32_835 ();
 sg13g2_fill_1 FILLER_32_837 ();
 sg13g2_decap_8 FILLER_32_852 ();
 sg13g2_fill_2 FILLER_32_859 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_18 ();
 sg13g2_decap_8 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_32 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_fill_2 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_4 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_64 ();
 sg13g2_decap_8 FILLER_33_82 ();
 sg13g2_decap_4 FILLER_33_89 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_116 ();
 sg13g2_decap_4 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_4 FILLER_33_214 ();
 sg13g2_decap_4 FILLER_33_223 ();
 sg13g2_fill_2 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_264 ();
 sg13g2_decap_8 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_4 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_4 FILLER_33_421 ();
 sg13g2_fill_1 FILLER_33_425 ();
 sg13g2_decap_8 FILLER_33_445 ();
 sg13g2_decap_8 FILLER_33_452 ();
 sg13g2_decap_8 FILLER_33_459 ();
 sg13g2_decap_4 FILLER_33_478 ();
 sg13g2_fill_1 FILLER_33_482 ();
 sg13g2_decap_8 FILLER_33_491 ();
 sg13g2_decap_8 FILLER_33_498 ();
 sg13g2_decap_4 FILLER_33_505 ();
 sg13g2_fill_2 FILLER_33_509 ();
 sg13g2_fill_2 FILLER_33_519 ();
 sg13g2_decap_8 FILLER_33_538 ();
 sg13g2_fill_2 FILLER_33_545 ();
 sg13g2_decap_4 FILLER_33_552 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_4 FILLER_33_595 ();
 sg13g2_fill_2 FILLER_33_599 ();
 sg13g2_decap_8 FILLER_33_612 ();
 sg13g2_decap_8 FILLER_33_619 ();
 sg13g2_decap_4 FILLER_33_626 ();
 sg13g2_fill_2 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_646 ();
 sg13g2_fill_1 FILLER_33_653 ();
 sg13g2_decap_4 FILLER_33_660 ();
 sg13g2_fill_2 FILLER_33_664 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_fill_1 FILLER_33_686 ();
 sg13g2_decap_4 FILLER_33_693 ();
 sg13g2_fill_2 FILLER_33_697 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_4 FILLER_33_714 ();
 sg13g2_fill_2 FILLER_33_718 ();
 sg13g2_decap_8 FILLER_33_725 ();
 sg13g2_decap_8 FILLER_33_732 ();
 sg13g2_decap_4 FILLER_33_739 ();
 sg13g2_decap_8 FILLER_33_748 ();
 sg13g2_decap_4 FILLER_33_755 ();
 sg13g2_fill_1 FILLER_33_759 ();
 sg13g2_decap_8 FILLER_33_769 ();
 sg13g2_decap_8 FILLER_33_776 ();
 sg13g2_decap_4 FILLER_33_783 ();
 sg13g2_fill_2 FILLER_33_787 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_fill_2 FILLER_33_816 ();
 sg13g2_fill_1 FILLER_33_818 ();
 sg13g2_decap_8 FILLER_33_823 ();
 sg13g2_decap_4 FILLER_33_830 ();
 sg13g2_fill_2 FILLER_33_834 ();
 sg13g2_decap_4 FILLER_33_858 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_27 ();
 sg13g2_fill_1 FILLER_34_45 ();
 sg13g2_decap_4 FILLER_34_52 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_decap_8 FILLER_34_79 ();
 sg13g2_decap_4 FILLER_34_86 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_decap_4 FILLER_34_107 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_131 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_decap_4 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_decap_4 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_decap_4 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_decap_8 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_decap_4 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_fill_1 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_fill_2 FILLER_34_396 ();
 sg13g2_fill_1 FILLER_34_398 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_414 ();
 sg13g2_decap_8 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_34_430 ();
 sg13g2_decap_4 FILLER_34_437 ();
 sg13g2_decap_8 FILLER_34_466 ();
 sg13g2_fill_2 FILLER_34_473 ();
 sg13g2_fill_2 FILLER_34_479 ();
 sg13g2_fill_1 FILLER_34_481 ();
 sg13g2_decap_8 FILLER_34_487 ();
 sg13g2_fill_1 FILLER_34_494 ();
 sg13g2_decap_8 FILLER_34_515 ();
 sg13g2_fill_1 FILLER_34_522 ();
 sg13g2_decap_4 FILLER_34_531 ();
 sg13g2_fill_2 FILLER_34_535 ();
 sg13g2_decap_8 FILLER_34_542 ();
 sg13g2_decap_4 FILLER_34_549 ();
 sg13g2_fill_1 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_565 ();
 sg13g2_fill_2 FILLER_34_572 ();
 sg13g2_fill_1 FILLER_34_574 ();
 sg13g2_decap_4 FILLER_34_597 ();
 sg13g2_fill_1 FILLER_34_601 ();
 sg13g2_fill_2 FILLER_34_606 ();
 sg13g2_decap_8 FILLER_34_625 ();
 sg13g2_decap_4 FILLER_34_632 ();
 sg13g2_fill_1 FILLER_34_636 ();
 sg13g2_fill_2 FILLER_34_650 ();
 sg13g2_decap_8 FILLER_34_657 ();
 sg13g2_decap_8 FILLER_34_664 ();
 sg13g2_fill_2 FILLER_34_677 ();
 sg13g2_decap_4 FILLER_34_683 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_fill_1 FILLER_34_705 ();
 sg13g2_fill_1 FILLER_34_711 ();
 sg13g2_decap_4 FILLER_34_717 ();
 sg13g2_decap_8 FILLER_34_737 ();
 sg13g2_fill_1 FILLER_34_759 ();
 sg13g2_decap_4 FILLER_34_781 ();
 sg13g2_fill_2 FILLER_34_785 ();
 sg13g2_decap_8 FILLER_34_800 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_fill_2 FILLER_34_814 ();
 sg13g2_decap_4 FILLER_34_837 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_decap_8 FILLER_35_29 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_decap_8 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_62 ();
 sg13g2_fill_2 FILLER_35_69 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_88 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_160 ();
 sg13g2_decap_4 FILLER_35_167 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_decap_4 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_212 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_decap_4 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_decap_8 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_4 FILLER_35_358 ();
 sg13g2_decap_4 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_4 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_411 ();
 sg13g2_decap_8 FILLER_35_435 ();
 sg13g2_decap_8 FILLER_35_442 ();
 sg13g2_decap_4 FILLER_35_449 ();
 sg13g2_decap_8 FILLER_35_457 ();
 sg13g2_fill_2 FILLER_35_464 ();
 sg13g2_fill_2 FILLER_35_474 ();
 sg13g2_fill_1 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_485 ();
 sg13g2_decap_4 FILLER_35_498 ();
 sg13g2_fill_1 FILLER_35_502 ();
 sg13g2_decap_8 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_521 ();
 sg13g2_decap_8 FILLER_35_528 ();
 sg13g2_decap_8 FILLER_35_561 ();
 sg13g2_decap_8 FILLER_35_568 ();
 sg13g2_fill_2 FILLER_35_575 ();
 sg13g2_decap_8 FILLER_35_583 ();
 sg13g2_decap_8 FILLER_35_590 ();
 sg13g2_decap_8 FILLER_35_608 ();
 sg13g2_decap_8 FILLER_35_615 ();
 sg13g2_fill_2 FILLER_35_622 ();
 sg13g2_fill_2 FILLER_35_628 ();
 sg13g2_fill_1 FILLER_35_630 ();
 sg13g2_fill_2 FILLER_35_641 ();
 sg13g2_fill_1 FILLER_35_643 ();
 sg13g2_decap_4 FILLER_35_649 ();
 sg13g2_fill_2 FILLER_35_653 ();
 sg13g2_decap_4 FILLER_35_666 ();
 sg13g2_fill_2 FILLER_35_670 ();
 sg13g2_fill_2 FILLER_35_677 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_fill_2 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_715 ();
 sg13g2_fill_2 FILLER_35_722 ();
 sg13g2_fill_1 FILLER_35_724 ();
 sg13g2_decap_4 FILLER_35_731 ();
 sg13g2_decap_4 FILLER_35_743 ();
 sg13g2_fill_2 FILLER_35_747 ();
 sg13g2_decap_8 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_774 ();
 sg13g2_decap_4 FILLER_35_781 ();
 sg13g2_fill_2 FILLER_35_790 ();
 sg13g2_fill_1 FILLER_35_792 ();
 sg13g2_decap_4 FILLER_35_807 ();
 sg13g2_fill_2 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_decap_8 FILLER_35_832 ();
 sg13g2_fill_2 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_852 ();
 sg13g2_fill_2 FILLER_35_859 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_31 ();
 sg13g2_decap_8 FILLER_36_37 ();
 sg13g2_fill_2 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_decap_4 FILLER_36_51 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_71 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_fill_2 FILLER_36_90 ();
 sg13g2_decap_4 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_100 ();
 sg13g2_decap_8 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_157 ();
 sg13g2_fill_1 FILLER_36_164 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_4 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_decap_4 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_313 ();
 sg13g2_decap_8 FILLER_36_320 ();
 sg13g2_decap_4 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_decap_4 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_decap_4 FILLER_36_397 ();
 sg13g2_fill_1 FILLER_36_401 ();
 sg13g2_decap_8 FILLER_36_408 ();
 sg13g2_decap_4 FILLER_36_415 ();
 sg13g2_fill_2 FILLER_36_419 ();
 sg13g2_fill_1 FILLER_36_426 ();
 sg13g2_decap_8 FILLER_36_435 ();
 sg13g2_fill_2 FILLER_36_442 ();
 sg13g2_fill_1 FILLER_36_444 ();
 sg13g2_decap_8 FILLER_36_473 ();
 sg13g2_decap_4 FILLER_36_480 ();
 sg13g2_fill_1 FILLER_36_484 ();
 sg13g2_decap_8 FILLER_36_493 ();
 sg13g2_decap_8 FILLER_36_500 ();
 sg13g2_decap_4 FILLER_36_507 ();
 sg13g2_fill_2 FILLER_36_511 ();
 sg13g2_fill_2 FILLER_36_521 ();
 sg13g2_decap_8 FILLER_36_531 ();
 sg13g2_fill_2 FILLER_36_538 ();
 sg13g2_decap_8 FILLER_36_544 ();
 sg13g2_decap_8 FILLER_36_551 ();
 sg13g2_decap_8 FILLER_36_558 ();
 sg13g2_decap_8 FILLER_36_565 ();
 sg13g2_fill_1 FILLER_36_572 ();
 sg13g2_decap_8 FILLER_36_589 ();
 sg13g2_decap_4 FILLER_36_596 ();
 sg13g2_fill_2 FILLER_36_600 ();
 sg13g2_decap_4 FILLER_36_612 ();
 sg13g2_decap_8 FILLER_36_622 ();
 sg13g2_fill_1 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_639 ();
 sg13g2_decap_8 FILLER_36_646 ();
 sg13g2_decap_8 FILLER_36_671 ();
 sg13g2_decap_4 FILLER_36_678 ();
 sg13g2_decap_8 FILLER_36_699 ();
 sg13g2_fill_2 FILLER_36_706 ();
 sg13g2_decap_8 FILLER_36_717 ();
 sg13g2_decap_8 FILLER_36_724 ();
 sg13g2_decap_4 FILLER_36_731 ();
 sg13g2_fill_2 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_741 ();
 sg13g2_decap_8 FILLER_36_748 ();
 sg13g2_decap_4 FILLER_36_755 ();
 sg13g2_fill_1 FILLER_36_759 ();
 sg13g2_fill_2 FILLER_36_770 ();
 sg13g2_fill_1 FILLER_36_772 ();
 sg13g2_fill_1 FILLER_36_778 ();
 sg13g2_fill_1 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_790 ();
 sg13g2_decap_4 FILLER_36_797 ();
 sg13g2_fill_2 FILLER_36_806 ();
 sg13g2_fill_1 FILLER_36_808 ();
 sg13g2_decap_8 FILLER_36_853 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_32 ();
 sg13g2_fill_1 FILLER_37_36 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_decap_8 FILLER_37_74 ();
 sg13g2_decap_8 FILLER_37_81 ();
 sg13g2_decap_4 FILLER_37_88 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_decap_4 FILLER_37_103 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_decap_8 FILLER_37_130 ();
 sg13g2_decap_4 FILLER_37_137 ();
 sg13g2_fill_1 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_156 ();
 sg13g2_decap_4 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_decap_4 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_212 ();
 sg13g2_decap_8 FILLER_37_227 ();
 sg13g2_decap_4 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_261 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_4 FILLER_37_365 ();
 sg13g2_fill_2 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_4 FILLER_37_392 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_4 FILLER_37_420 ();
 sg13g2_fill_2 FILLER_37_443 ();
 sg13g2_fill_1 FILLER_37_445 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_4 FILLER_37_483 ();
 sg13g2_fill_1 FILLER_37_487 ();
 sg13g2_decap_8 FILLER_37_494 ();
 sg13g2_decap_4 FILLER_37_501 ();
 sg13g2_fill_1 FILLER_37_505 ();
 sg13g2_decap_8 FILLER_37_523 ();
 sg13g2_decap_8 FILLER_37_530 ();
 sg13g2_decap_4 FILLER_37_537 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_decap_4 FILLER_37_563 ();
 sg13g2_fill_1 FILLER_37_567 ();
 sg13g2_decap_4 FILLER_37_579 ();
 sg13g2_fill_1 FILLER_37_583 ();
 sg13g2_fill_2 FILLER_37_592 ();
 sg13g2_fill_2 FILLER_37_625 ();
 sg13g2_fill_1 FILLER_37_627 ();
 sg13g2_decap_8 FILLER_37_646 ();
 sg13g2_fill_1 FILLER_37_653 ();
 sg13g2_decap_4 FILLER_37_663 ();
 sg13g2_fill_2 FILLER_37_667 ();
 sg13g2_decap_4 FILLER_37_679 ();
 sg13g2_fill_1 FILLER_37_683 ();
 sg13g2_decap_8 FILLER_37_689 ();
 sg13g2_decap_8 FILLER_37_696 ();
 sg13g2_decap_4 FILLER_37_725 ();
 sg13g2_fill_2 FILLER_37_729 ();
 sg13g2_fill_1 FILLER_37_738 ();
 sg13g2_decap_4 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_769 ();
 sg13g2_decap_4 FILLER_37_776 ();
 sg13g2_fill_1 FILLER_37_780 ();
 sg13g2_decap_4 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_801 ();
 sg13g2_decap_8 FILLER_37_808 ();
 sg13g2_fill_1 FILLER_37_815 ();
 sg13g2_fill_1 FILLER_37_820 ();
 sg13g2_decap_8 FILLER_37_831 ();
 sg13g2_fill_2 FILLER_37_838 ();
 sg13g2_decap_8 FILLER_37_844 ();
 sg13g2_decap_8 FILLER_37_851 ();
 sg13g2_decap_4 FILLER_37_858 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_11 ();
 sg13g2_fill_2 FILLER_38_22 ();
 sg13g2_fill_1 FILLER_38_24 ();
 sg13g2_decap_4 FILLER_38_35 ();
 sg13g2_decap_4 FILLER_38_47 ();
 sg13g2_fill_1 FILLER_38_51 ();
 sg13g2_fill_2 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_57 ();
 sg13g2_decap_8 FILLER_38_71 ();
 sg13g2_fill_1 FILLER_38_78 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_101 ();
 sg13g2_decap_8 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_decap_8 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_4 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_4 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_4 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_4 FILLER_38_358 ();
 sg13g2_fill_2 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_394 ();
 sg13g2_fill_1 FILLER_38_396 ();
 sg13g2_decap_8 FILLER_38_405 ();
 sg13g2_decap_8 FILLER_38_412 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_426 ();
 sg13g2_decap_8 FILLER_38_440 ();
 sg13g2_decap_8 FILLER_38_447 ();
 sg13g2_fill_2 FILLER_38_454 ();
 sg13g2_decap_8 FILLER_38_460 ();
 sg13g2_fill_2 FILLER_38_467 ();
 sg13g2_fill_1 FILLER_38_478 ();
 sg13g2_fill_1 FILLER_38_484 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_fill_2 FILLER_38_497 ();
 sg13g2_decap_4 FILLER_38_509 ();
 sg13g2_fill_1 FILLER_38_523 ();
 sg13g2_fill_1 FILLER_38_537 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_4 FILLER_38_553 ();
 sg13g2_fill_1 FILLER_38_557 ();
 sg13g2_fill_2 FILLER_38_563 ();
 sg13g2_decap_8 FILLER_38_589 ();
 sg13g2_decap_8 FILLER_38_596 ();
 sg13g2_decap_8 FILLER_38_603 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_decap_4 FILLER_38_617 ();
 sg13g2_fill_2 FILLER_38_621 ();
 sg13g2_fill_2 FILLER_38_629 ();
 sg13g2_fill_2 FILLER_38_636 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_4 FILLER_38_672 ();
 sg13g2_fill_2 FILLER_38_681 ();
 sg13g2_fill_1 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_697 ();
 sg13g2_fill_2 FILLER_38_704 ();
 sg13g2_fill_2 FILLER_38_711 ();
 sg13g2_decap_8 FILLER_38_718 ();
 sg13g2_decap_4 FILLER_38_725 ();
 sg13g2_fill_1 FILLER_38_737 ();
 sg13g2_decap_8 FILLER_38_744 ();
 sg13g2_decap_8 FILLER_38_751 ();
 sg13g2_decap_4 FILLER_38_758 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_fill_1 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_fill_2 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_fill_1 FILLER_38_830 ();
 sg13g2_decap_4 FILLER_38_838 ();
 sg13g2_fill_1 FILLER_38_842 ();
 sg13g2_fill_2 FILLER_38_859 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_18 ();
 sg13g2_fill_1 FILLER_39_25 ();
 sg13g2_decap_4 FILLER_39_31 ();
 sg13g2_fill_1 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_68 ();
 sg13g2_decap_4 FILLER_39_75 ();
 sg13g2_fill_2 FILLER_39_79 ();
 sg13g2_fill_1 FILLER_39_90 ();
 sg13g2_decap_4 FILLER_39_100 ();
 sg13g2_decap_8 FILLER_39_114 ();
 sg13g2_decap_4 FILLER_39_121 ();
 sg13g2_decap_8 FILLER_39_137 ();
 sg13g2_decap_8 FILLER_39_144 ();
 sg13g2_decap_8 FILLER_39_151 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_218 ();
 sg13g2_fill_2 FILLER_39_225 ();
 sg13g2_decap_4 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_247 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_decap_8 FILLER_39_293 ();
 sg13g2_decap_4 FILLER_39_305 ();
 sg13g2_fill_2 FILLER_39_319 ();
 sg13g2_fill_2 FILLER_39_326 ();
 sg13g2_fill_1 FILLER_39_328 ();
 sg13g2_fill_2 FILLER_39_339 ();
 sg13g2_fill_1 FILLER_39_341 ();
 sg13g2_decap_4 FILLER_39_359 ();
 sg13g2_fill_2 FILLER_39_363 ();
 sg13g2_fill_2 FILLER_39_384 ();
 sg13g2_fill_1 FILLER_39_386 ();
 sg13g2_fill_2 FILLER_39_398 ();
 sg13g2_fill_1 FILLER_39_400 ();
 sg13g2_fill_1 FILLER_39_406 ();
 sg13g2_decap_4 FILLER_39_416 ();
 sg13g2_decap_4 FILLER_39_433 ();
 sg13g2_fill_2 FILLER_39_437 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_fill_2 FILLER_39_462 ();
 sg13g2_fill_1 FILLER_39_464 ();
 sg13g2_fill_1 FILLER_39_470 ();
 sg13g2_decap_8 FILLER_39_486 ();
 sg13g2_decap_4 FILLER_39_499 ();
 sg13g2_decap_8 FILLER_39_509 ();
 sg13g2_decap_8 FILLER_39_516 ();
 sg13g2_decap_4 FILLER_39_523 ();
 sg13g2_fill_1 FILLER_39_527 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_4 FILLER_39_546 ();
 sg13g2_fill_1 FILLER_39_554 ();
 sg13g2_decap_8 FILLER_39_562 ();
 sg13g2_decap_4 FILLER_39_569 ();
 sg13g2_fill_1 FILLER_39_573 ();
 sg13g2_fill_2 FILLER_39_582 ();
 sg13g2_fill_1 FILLER_39_584 ();
 sg13g2_decap_8 FILLER_39_590 ();
 sg13g2_fill_1 FILLER_39_597 ();
 sg13g2_fill_1 FILLER_39_606 ();
 sg13g2_decap_8 FILLER_39_618 ();
 sg13g2_fill_2 FILLER_39_625 ();
 sg13g2_fill_1 FILLER_39_627 ();
 sg13g2_decap_8 FILLER_39_633 ();
 sg13g2_decap_8 FILLER_39_640 ();
 sg13g2_decap_8 FILLER_39_647 ();
 sg13g2_decap_8 FILLER_39_654 ();
 sg13g2_decap_8 FILLER_39_661 ();
 sg13g2_decap_8 FILLER_39_668 ();
 sg13g2_fill_2 FILLER_39_675 ();
 sg13g2_fill_2 FILLER_39_682 ();
 sg13g2_fill_1 FILLER_39_684 ();
 sg13g2_decap_8 FILLER_39_690 ();
 sg13g2_fill_2 FILLER_39_705 ();
 sg13g2_decap_8 FILLER_39_723 ();
 sg13g2_fill_2 FILLER_39_730 ();
 sg13g2_fill_1 FILLER_39_737 ();
 sg13g2_decap_4 FILLER_39_752 ();
 sg13g2_decap_4 FILLER_39_761 ();
 sg13g2_fill_1 FILLER_39_765 ();
 sg13g2_decap_4 FILLER_39_791 ();
 sg13g2_fill_1 FILLER_39_795 ();
 sg13g2_decap_8 FILLER_39_825 ();
 sg13g2_decap_8 FILLER_39_832 ();
 sg13g2_decap_8 FILLER_39_853 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_23 ();
 sg13g2_decap_8 FILLER_40_29 ();
 sg13g2_decap_4 FILLER_40_36 ();
 sg13g2_fill_2 FILLER_40_40 ();
 sg13g2_decap_8 FILLER_40_50 ();
 sg13g2_decap_8 FILLER_40_57 ();
 sg13g2_fill_1 FILLER_40_64 ();
 sg13g2_decap_8 FILLER_40_75 ();
 sg13g2_decap_8 FILLER_40_82 ();
 sg13g2_decap_8 FILLER_40_89 ();
 sg13g2_decap_4 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_108 ();
 sg13g2_fill_1 FILLER_40_110 ();
 sg13g2_decap_8 FILLER_40_142 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_fill_2 FILLER_40_164 ();
 sg13g2_fill_1 FILLER_40_166 ();
 sg13g2_decap_8 FILLER_40_187 ();
 sg13g2_decap_8 FILLER_40_194 ();
 sg13g2_decap_4 FILLER_40_201 ();
 sg13g2_fill_2 FILLER_40_205 ();
 sg13g2_decap_8 FILLER_40_221 ();
 sg13g2_decap_8 FILLER_40_228 ();
 sg13g2_decap_8 FILLER_40_235 ();
 sg13g2_fill_2 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_244 ();
 sg13g2_decap_8 FILLER_40_250 ();
 sg13g2_fill_1 FILLER_40_257 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_4 FILLER_40_273 ();
 sg13g2_fill_2 FILLER_40_277 ();
 sg13g2_decap_8 FILLER_40_285 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_fill_2 FILLER_40_315 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_323 ();
 sg13g2_decap_4 FILLER_40_329 ();
 sg13g2_fill_2 FILLER_40_333 ();
 sg13g2_decap_4 FILLER_40_341 ();
 sg13g2_fill_1 FILLER_40_345 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_4 FILLER_40_378 ();
 sg13g2_fill_2 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_fill_2 FILLER_40_397 ();
 sg13g2_decap_8 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_40_415 ();
 sg13g2_fill_2 FILLER_40_422 ();
 sg13g2_fill_1 FILLER_40_424 ();
 sg13g2_decap_4 FILLER_40_431 ();
 sg13g2_fill_2 FILLER_40_435 ();
 sg13g2_decap_8 FILLER_40_453 ();
 sg13g2_decap_8 FILLER_40_460 ();
 sg13g2_fill_2 FILLER_40_490 ();
 sg13g2_fill_1 FILLER_40_500 ();
 sg13g2_decap_4 FILLER_40_536 ();
 sg13g2_fill_1 FILLER_40_552 ();
 sg13g2_decap_8 FILLER_40_558 ();
 sg13g2_decap_4 FILLER_40_565 ();
 sg13g2_fill_1 FILLER_40_569 ();
 sg13g2_decap_8 FILLER_40_578 ();
 sg13g2_decap_8 FILLER_40_585 ();
 sg13g2_decap_8 FILLER_40_592 ();
 sg13g2_decap_4 FILLER_40_599 ();
 sg13g2_fill_2 FILLER_40_603 ();
 sg13g2_decap_4 FILLER_40_614 ();
 sg13g2_fill_1 FILLER_40_618 ();
 sg13g2_fill_1 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_642 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_695 ();
 sg13g2_decap_8 FILLER_40_702 ();
 sg13g2_decap_8 FILLER_40_718 ();
 sg13g2_decap_8 FILLER_40_725 ();
 sg13g2_decap_8 FILLER_40_732 ();
 sg13g2_fill_2 FILLER_40_739 ();
 sg13g2_fill_1 FILLER_40_741 ();
 sg13g2_fill_2 FILLER_40_750 ();
 sg13g2_fill_1 FILLER_40_752 ();
 sg13g2_fill_2 FILLER_40_763 ();
 sg13g2_fill_1 FILLER_40_765 ();
 sg13g2_decap_4 FILLER_40_771 ();
 sg13g2_decap_8 FILLER_40_780 ();
 sg13g2_decap_8 FILLER_40_787 ();
 sg13g2_decap_8 FILLER_40_794 ();
 sg13g2_decap_4 FILLER_40_801 ();
 sg13g2_fill_2 FILLER_40_805 ();
 sg13g2_fill_1 FILLER_40_811 ();
 sg13g2_decap_4 FILLER_40_826 ();
 sg13g2_fill_1 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_855 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_58 ();
 sg13g2_fill_1 FILLER_41_60 ();
 sg13g2_decap_4 FILLER_41_67 ();
 sg13g2_decap_4 FILLER_41_93 ();
 sg13g2_decap_8 FILLER_41_114 ();
 sg13g2_decap_4 FILLER_41_121 ();
 sg13g2_decap_8 FILLER_41_135 ();
 sg13g2_fill_2 FILLER_41_142 ();
 sg13g2_fill_2 FILLER_41_158 ();
 sg13g2_fill_2 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_fill_1 FILLER_41_182 ();
 sg13g2_fill_2 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_222 ();
 sg13g2_decap_4 FILLER_41_229 ();
 sg13g2_fill_2 FILLER_41_233 ();
 sg13g2_fill_1 FILLER_41_251 ();
 sg13g2_decap_8 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_fill_1 FILLER_41_308 ();
 sg13g2_fill_2 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_4 FILLER_41_362 ();
 sg13g2_decap_4 FILLER_41_387 ();
 sg13g2_decap_8 FILLER_41_395 ();
 sg13g2_decap_8 FILLER_41_410 ();
 sg13g2_decap_4 FILLER_41_417 ();
 sg13g2_fill_2 FILLER_41_421 ();
 sg13g2_decap_8 FILLER_41_442 ();
 sg13g2_fill_2 FILLER_41_449 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_4 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_509 ();
 sg13g2_decap_8 FILLER_41_516 ();
 sg13g2_decap_8 FILLER_41_523 ();
 sg13g2_fill_2 FILLER_41_530 ();
 sg13g2_decap_4 FILLER_41_543 ();
 sg13g2_fill_1 FILLER_41_547 ();
 sg13g2_fill_2 FILLER_41_553 ();
 sg13g2_fill_1 FILLER_41_555 ();
 sg13g2_fill_1 FILLER_41_561 ();
 sg13g2_decap_4 FILLER_41_570 ();
 sg13g2_fill_2 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_584 ();
 sg13g2_fill_1 FILLER_41_608 ();
 sg13g2_decap_8 FILLER_41_622 ();
 sg13g2_fill_1 FILLER_41_634 ();
 sg13g2_fill_2 FILLER_41_645 ();
 sg13g2_decap_8 FILLER_41_656 ();
 sg13g2_decap_4 FILLER_41_663 ();
 sg13g2_fill_2 FILLER_41_667 ();
 sg13g2_decap_8 FILLER_41_674 ();
 sg13g2_fill_2 FILLER_41_681 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_4 FILLER_41_703 ();
 sg13g2_fill_1 FILLER_41_707 ();
 sg13g2_fill_2 FILLER_41_724 ();
 sg13g2_fill_1 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_746 ();
 sg13g2_decap_8 FILLER_41_753 ();
 sg13g2_fill_2 FILLER_41_760 ();
 sg13g2_fill_1 FILLER_41_762 ();
 sg13g2_decap_4 FILLER_41_774 ();
 sg13g2_fill_1 FILLER_41_786 ();
 sg13g2_decap_8 FILLER_41_804 ();
 sg13g2_decap_8 FILLER_41_811 ();
 sg13g2_decap_4 FILLER_41_834 ();
 sg13g2_fill_1 FILLER_41_838 ();
 sg13g2_decap_4 FILLER_41_857 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_4 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_32 ();
 sg13g2_fill_2 FILLER_42_38 ();
 sg13g2_decap_8 FILLER_42_45 ();
 sg13g2_decap_8 FILLER_42_52 ();
 sg13g2_decap_8 FILLER_42_59 ();
 sg13g2_fill_1 FILLER_42_66 ();
 sg13g2_decap_8 FILLER_42_76 ();
 sg13g2_decap_4 FILLER_42_83 ();
 sg13g2_fill_1 FILLER_42_87 ();
 sg13g2_decap_4 FILLER_42_93 ();
 sg13g2_fill_2 FILLER_42_97 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_fill_2 FILLER_42_119 ();
 sg13g2_decap_4 FILLER_42_139 ();
 sg13g2_decap_4 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_152 ();
 sg13g2_decap_8 FILLER_42_158 ();
 sg13g2_decap_4 FILLER_42_165 ();
 sg13g2_decap_4 FILLER_42_179 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_fill_2 FILLER_42_192 ();
 sg13g2_decap_8 FILLER_42_199 ();
 sg13g2_decap_4 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_fill_2 FILLER_42_219 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_decap_4 FILLER_42_249 ();
 sg13g2_decap_4 FILLER_42_268 ();
 sg13g2_fill_2 FILLER_42_290 ();
 sg13g2_fill_1 FILLER_42_292 ();
 sg13g2_fill_2 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_313 ();
 sg13g2_decap_8 FILLER_42_325 ();
 sg13g2_fill_2 FILLER_42_332 ();
 sg13g2_fill_1 FILLER_42_334 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_fill_2 FILLER_42_378 ();
 sg13g2_fill_1 FILLER_42_380 ();
 sg13g2_fill_1 FILLER_42_393 ();
 sg13g2_decap_8 FILLER_42_409 ();
 sg13g2_decap_4 FILLER_42_422 ();
 sg13g2_fill_2 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_42_435 ();
 sg13g2_decap_8 FILLER_42_442 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_decap_4 FILLER_42_468 ();
 sg13g2_fill_2 FILLER_42_472 ();
 sg13g2_fill_2 FILLER_42_478 ();
 sg13g2_decap_8 FILLER_42_491 ();
 sg13g2_fill_2 FILLER_42_498 ();
 sg13g2_fill_1 FILLER_42_500 ();
 sg13g2_decap_8 FILLER_42_507 ();
 sg13g2_fill_2 FILLER_42_514 ();
 sg13g2_fill_1 FILLER_42_516 ();
 sg13g2_decap_4 FILLER_42_522 ();
 sg13g2_fill_1 FILLER_42_526 ();
 sg13g2_decap_8 FILLER_42_542 ();
 sg13g2_decap_8 FILLER_42_549 ();
 sg13g2_decap_8 FILLER_42_567 ();
 sg13g2_fill_2 FILLER_42_574 ();
 sg13g2_fill_2 FILLER_42_592 ();
 sg13g2_decap_8 FILLER_42_598 ();
 sg13g2_decap_4 FILLER_42_614 ();
 sg13g2_fill_2 FILLER_42_623 ();
 sg13g2_fill_1 FILLER_42_625 ();
 sg13g2_decap_8 FILLER_42_632 ();
 sg13g2_fill_1 FILLER_42_639 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_fill_2 FILLER_42_651 ();
 sg13g2_decap_4 FILLER_42_664 ();
 sg13g2_fill_1 FILLER_42_668 ();
 sg13g2_decap_8 FILLER_42_674 ();
 sg13g2_fill_2 FILLER_42_681 ();
 sg13g2_fill_1 FILLER_42_683 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_718 ();
 sg13g2_decap_4 FILLER_42_725 ();
 sg13g2_decap_8 FILLER_42_738 ();
 sg13g2_decap_4 FILLER_42_745 ();
 sg13g2_fill_1 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_4 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_fill_2 FILLER_42_784 ();
 sg13g2_fill_1 FILLER_42_786 ();
 sg13g2_fill_2 FILLER_42_792 ();
 sg13g2_decap_8 FILLER_42_802 ();
 sg13g2_decap_8 FILLER_42_809 ();
 sg13g2_fill_1 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_4 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_852 ();
 sg13g2_fill_2 FILLER_42_859 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_29 ();
 sg13g2_decap_8 FILLER_43_36 ();
 sg13g2_decap_4 FILLER_43_43 ();
 sg13g2_fill_2 FILLER_43_66 ();
 sg13g2_fill_1 FILLER_43_68 ();
 sg13g2_fill_1 FILLER_43_73 ();
 sg13g2_decap_4 FILLER_43_79 ();
 sg13g2_fill_2 FILLER_43_83 ();
 sg13g2_fill_2 FILLER_43_93 ();
 sg13g2_fill_1 FILLER_43_95 ();
 sg13g2_decap_4 FILLER_43_112 ();
 sg13g2_decap_4 FILLER_43_124 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_decap_8 FILLER_43_134 ();
 sg13g2_decap_4 FILLER_43_141 ();
 sg13g2_fill_2 FILLER_43_145 ();
 sg13g2_fill_1 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_174 ();
 sg13g2_decap_8 FILLER_43_183 ();
 sg13g2_decap_4 FILLER_43_190 ();
 sg13g2_fill_2 FILLER_43_194 ();
 sg13g2_fill_1 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_216 ();
 sg13g2_decap_8 FILLER_43_223 ();
 sg13g2_decap_8 FILLER_43_230 ();
 sg13g2_decap_4 FILLER_43_243 ();
 sg13g2_fill_2 FILLER_43_247 ();
 sg13g2_decap_4 FILLER_43_253 ();
 sg13g2_decap_8 FILLER_43_265 ();
 sg13g2_decap_8 FILLER_43_272 ();
 sg13g2_decap_8 FILLER_43_279 ();
 sg13g2_decap_8 FILLER_43_297 ();
 sg13g2_decap_8 FILLER_43_304 ();
 sg13g2_decap_8 FILLER_43_311 ();
 sg13g2_decap_8 FILLER_43_318 ();
 sg13g2_fill_1 FILLER_43_325 ();
 sg13g2_decap_8 FILLER_43_331 ();
 sg13g2_fill_1 FILLER_43_338 ();
 sg13g2_decap_8 FILLER_43_356 ();
 sg13g2_decap_8 FILLER_43_363 ();
 sg13g2_decap_8 FILLER_43_384 ();
 sg13g2_decap_8 FILLER_43_391 ();
 sg13g2_decap_8 FILLER_43_398 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_4 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_449 ();
 sg13g2_decap_8 FILLER_43_456 ();
 sg13g2_decap_4 FILLER_43_463 ();
 sg13g2_fill_2 FILLER_43_467 ();
 sg13g2_decap_4 FILLER_43_474 ();
 sg13g2_fill_1 FILLER_43_478 ();
 sg13g2_decap_8 FILLER_43_484 ();
 sg13g2_decap_4 FILLER_43_491 ();
 sg13g2_decap_4 FILLER_43_513 ();
 sg13g2_fill_1 FILLER_43_517 ();
 sg13g2_decap_8 FILLER_43_523 ();
 sg13g2_fill_2 FILLER_43_530 ();
 sg13g2_decap_8 FILLER_43_548 ();
 sg13g2_decap_8 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_562 ();
 sg13g2_fill_1 FILLER_43_580 ();
 sg13g2_decap_8 FILLER_43_591 ();
 sg13g2_decap_8 FILLER_43_598 ();
 sg13g2_decap_4 FILLER_43_605 ();
 sg13g2_decap_8 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_621 ();
 sg13g2_decap_4 FILLER_43_628 ();
 sg13g2_fill_1 FILLER_43_638 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_fill_2 FILLER_43_682 ();
 sg13g2_fill_1 FILLER_43_684 ();
 sg13g2_decap_8 FILLER_43_690 ();
 sg13g2_decap_8 FILLER_43_697 ();
 sg13g2_decap_8 FILLER_43_704 ();
 sg13g2_fill_2 FILLER_43_711 ();
 sg13g2_decap_4 FILLER_43_728 ();
 sg13g2_fill_1 FILLER_43_732 ();
 sg13g2_fill_1 FILLER_43_762 ();
 sg13g2_decap_8 FILLER_43_776 ();
 sg13g2_decap_8 FILLER_43_783 ();
 sg13g2_fill_2 FILLER_43_790 ();
 sg13g2_decap_8 FILLER_43_802 ();
 sg13g2_decap_4 FILLER_43_809 ();
 sg13g2_fill_2 FILLER_43_813 ();
 sg13g2_fill_2 FILLER_43_833 ();
 sg13g2_decap_4 FILLER_43_857 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_4 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_33 ();
 sg13g2_decap_4 FILLER_44_40 ();
 sg13g2_fill_1 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_67 ();
 sg13g2_decap_8 FILLER_44_74 ();
 sg13g2_fill_1 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_90 ();
 sg13g2_decap_4 FILLER_44_97 ();
 sg13g2_decap_8 FILLER_44_106 ();
 sg13g2_fill_2 FILLER_44_113 ();
 sg13g2_fill_1 FILLER_44_115 ();
 sg13g2_decap_8 FILLER_44_121 ();
 sg13g2_fill_2 FILLER_44_128 ();
 sg13g2_fill_1 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_136 ();
 sg13g2_decap_4 FILLER_44_143 ();
 sg13g2_fill_1 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_164 ();
 sg13g2_fill_2 FILLER_44_171 ();
 sg13g2_decap_8 FILLER_44_179 ();
 sg13g2_decap_4 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_200 ();
 sg13g2_fill_2 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_218 ();
 sg13g2_decap_4 FILLER_44_225 ();
 sg13g2_decap_8 FILLER_44_237 ();
 sg13g2_fill_2 FILLER_44_244 ();
 sg13g2_fill_1 FILLER_44_246 ();
 sg13g2_fill_1 FILLER_44_260 ();
 sg13g2_decap_8 FILLER_44_275 ();
 sg13g2_fill_2 FILLER_44_282 ();
 sg13g2_decap_4 FILLER_44_297 ();
 sg13g2_fill_1 FILLER_44_301 ();
 sg13g2_decap_4 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_332 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_4 FILLER_44_371 ();
 sg13g2_fill_1 FILLER_44_375 ();
 sg13g2_fill_1 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_397 ();
 sg13g2_decap_8 FILLER_44_404 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_decap_4 FILLER_44_431 ();
 sg13g2_fill_2 FILLER_44_435 ();
 sg13g2_decap_4 FILLER_44_449 ();
 sg13g2_fill_2 FILLER_44_461 ();
 sg13g2_fill_1 FILLER_44_463 ();
 sg13g2_decap_8 FILLER_44_478 ();
 sg13g2_decap_8 FILLER_44_501 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_fill_2 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_530 ();
 sg13g2_decap_8 FILLER_44_537 ();
 sg13g2_decap_8 FILLER_44_544 ();
 sg13g2_decap_4 FILLER_44_554 ();
 sg13g2_fill_1 FILLER_44_558 ();
 sg13g2_decap_8 FILLER_44_582 ();
 sg13g2_fill_1 FILLER_44_589 ();
 sg13g2_decap_4 FILLER_44_611 ();
 sg13g2_fill_2 FILLER_44_634 ();
 sg13g2_decap_8 FILLER_44_641 ();
 sg13g2_decap_8 FILLER_44_648 ();
 sg13g2_fill_2 FILLER_44_655 ();
 sg13g2_fill_1 FILLER_44_657 ();
 sg13g2_decap_4 FILLER_44_681 ();
 sg13g2_fill_1 FILLER_44_685 ();
 sg13g2_decap_8 FILLER_44_712 ();
 sg13g2_decap_4 FILLER_44_719 ();
 sg13g2_fill_1 FILLER_44_723 ();
 sg13g2_decap_8 FILLER_44_732 ();
 sg13g2_decap_8 FILLER_44_739 ();
 sg13g2_decap_8 FILLER_44_746 ();
 sg13g2_decap_8 FILLER_44_753 ();
 sg13g2_decap_4 FILLER_44_776 ();
 sg13g2_fill_2 FILLER_44_780 ();
 sg13g2_decap_8 FILLER_44_806 ();
 sg13g2_fill_2 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_815 ();
 sg13g2_decap_8 FILLER_44_821 ();
 sg13g2_decap_8 FILLER_44_828 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_4 FILLER_44_857 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_25 ();
 sg13g2_decap_4 FILLER_45_36 ();
 sg13g2_fill_2 FILLER_45_44 ();
 sg13g2_decap_4 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_65 ();
 sg13g2_fill_2 FILLER_45_72 ();
 sg13g2_fill_2 FILLER_45_94 ();
 sg13g2_decap_4 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_106 ();
 sg13g2_decap_4 FILLER_45_118 ();
 sg13g2_decap_8 FILLER_45_141 ();
 sg13g2_decap_4 FILLER_45_148 ();
 sg13g2_fill_2 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_165 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_decap_4 FILLER_45_186 ();
 sg13g2_decap_8 FILLER_45_208 ();
 sg13g2_decap_8 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_fill_1 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_4 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_295 ();
 sg13g2_decap_8 FILLER_45_310 ();
 sg13g2_decap_4 FILLER_45_317 ();
 sg13g2_fill_2 FILLER_45_321 ();
 sg13g2_fill_1 FILLER_45_333 ();
 sg13g2_fill_2 FILLER_45_348 ();
 sg13g2_decap_8 FILLER_45_355 ();
 sg13g2_decap_4 FILLER_45_362 ();
 sg13g2_fill_1 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_fill_1 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_405 ();
 sg13g2_decap_4 FILLER_45_423 ();
 sg13g2_fill_2 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_447 ();
 sg13g2_fill_2 FILLER_45_454 ();
 sg13g2_decap_8 FILLER_45_478 ();
 sg13g2_fill_2 FILLER_45_485 ();
 sg13g2_fill_2 FILLER_45_496 ();
 sg13g2_fill_1 FILLER_45_498 ();
 sg13g2_fill_1 FILLER_45_504 ();
 sg13g2_fill_2 FILLER_45_519 ();
 sg13g2_fill_2 FILLER_45_527 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_decap_8 FILLER_45_557 ();
 sg13g2_fill_1 FILLER_45_564 ();
 sg13g2_decap_8 FILLER_45_569 ();
 sg13g2_decap_8 FILLER_45_579 ();
 sg13g2_decap_8 FILLER_45_586 ();
 sg13g2_decap_4 FILLER_45_593 ();
 sg13g2_decap_8 FILLER_45_602 ();
 sg13g2_fill_2 FILLER_45_609 ();
 sg13g2_decap_8 FILLER_45_616 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_decap_4 FILLER_45_630 ();
 sg13g2_fill_1 FILLER_45_634 ();
 sg13g2_fill_1 FILLER_45_640 ();
 sg13g2_fill_2 FILLER_45_651 ();
 sg13g2_fill_1 FILLER_45_653 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_672 ();
 sg13g2_fill_1 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_707 ();
 sg13g2_fill_2 FILLER_45_714 ();
 sg13g2_fill_1 FILLER_45_716 ();
 sg13g2_fill_2 FILLER_45_723 ();
 sg13g2_decap_4 FILLER_45_730 ();
 sg13g2_decap_8 FILLER_45_750 ();
 sg13g2_decap_4 FILLER_45_757 ();
 sg13g2_fill_2 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_4 FILLER_45_786 ();
 sg13g2_fill_2 FILLER_45_790 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_decap_4 FILLER_45_807 ();
 sg13g2_decap_4 FILLER_45_824 ();
 sg13g2_decap_4 FILLER_45_833 ();
 sg13g2_decap_8 FILLER_45_848 ();
 sg13g2_decap_8 FILLER_45_855 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_23 ();
 sg13g2_fill_2 FILLER_46_33 ();
 sg13g2_fill_1 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_55 ();
 sg13g2_decap_8 FILLER_46_61 ();
 sg13g2_decap_8 FILLER_46_68 ();
 sg13g2_decap_8 FILLER_46_86 ();
 sg13g2_decap_4 FILLER_46_93 ();
 sg13g2_decap_8 FILLER_46_111 ();
 sg13g2_decap_4 FILLER_46_118 ();
 sg13g2_fill_2 FILLER_46_122 ();
 sg13g2_decap_8 FILLER_46_141 ();
 sg13g2_fill_2 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_160 ();
 sg13g2_decap_8 FILLER_46_167 ();
 sg13g2_fill_1 FILLER_46_174 ();
 sg13g2_decap_8 FILLER_46_187 ();
 sg13g2_decap_4 FILLER_46_194 ();
 sg13g2_fill_1 FILLER_46_198 ();
 sg13g2_fill_1 FILLER_46_208 ();
 sg13g2_fill_2 FILLER_46_214 ();
 sg13g2_fill_1 FILLER_46_216 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_decap_8 FILLER_46_237 ();
 sg13g2_fill_1 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_249 ();
 sg13g2_decap_8 FILLER_46_264 ();
 sg13g2_fill_2 FILLER_46_271 ();
 sg13g2_decap_8 FILLER_46_300 ();
 sg13g2_decap_8 FILLER_46_307 ();
 sg13g2_fill_1 FILLER_46_314 ();
 sg13g2_decap_8 FILLER_46_325 ();
 sg13g2_decap_8 FILLER_46_332 ();
 sg13g2_decap_4 FILLER_46_339 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_decap_4 FILLER_46_351 ();
 sg13g2_decap_8 FILLER_46_363 ();
 sg13g2_decap_4 FILLER_46_370 ();
 sg13g2_decap_8 FILLER_46_387 ();
 sg13g2_fill_2 FILLER_46_394 ();
 sg13g2_fill_1 FILLER_46_396 ();
 sg13g2_fill_1 FILLER_46_411 ();
 sg13g2_decap_8 FILLER_46_418 ();
 sg13g2_decap_4 FILLER_46_425 ();
 sg13g2_fill_1 FILLER_46_434 ();
 sg13g2_fill_2 FILLER_46_439 ();
 sg13g2_decap_8 FILLER_46_452 ();
 sg13g2_decap_4 FILLER_46_459 ();
 sg13g2_decap_8 FILLER_46_468 ();
 sg13g2_decap_8 FILLER_46_475 ();
 sg13g2_decap_4 FILLER_46_482 ();
 sg13g2_decap_8 FILLER_46_491 ();
 sg13g2_decap_4 FILLER_46_498 ();
 sg13g2_fill_1 FILLER_46_502 ();
 sg13g2_decap_8 FILLER_46_507 ();
 sg13g2_fill_2 FILLER_46_514 ();
 sg13g2_fill_1 FILLER_46_516 ();
 sg13g2_decap_8 FILLER_46_522 ();
 sg13g2_decap_8 FILLER_46_529 ();
 sg13g2_decap_8 FILLER_46_536 ();
 sg13g2_fill_1 FILLER_46_543 ();
 sg13g2_decap_8 FILLER_46_548 ();
 sg13g2_fill_1 FILLER_46_555 ();
 sg13g2_fill_1 FILLER_46_567 ();
 sg13g2_decap_4 FILLER_46_582 ();
 sg13g2_fill_2 FILLER_46_586 ();
 sg13g2_fill_2 FILLER_46_596 ();
 sg13g2_decap_4 FILLER_46_606 ();
 sg13g2_fill_2 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_641 ();
 sg13g2_decap_4 FILLER_46_648 ();
 sg13g2_fill_1 FILLER_46_652 ();
 sg13g2_decap_4 FILLER_46_659 ();
 sg13g2_decap_4 FILLER_46_672 ();
 sg13g2_fill_1 FILLER_46_676 ();
 sg13g2_fill_2 FILLER_46_686 ();
 sg13g2_fill_1 FILLER_46_688 ();
 sg13g2_fill_1 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_699 ();
 sg13g2_decap_4 FILLER_46_706 ();
 sg13g2_fill_1 FILLER_46_710 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_4 FILLER_46_742 ();
 sg13g2_fill_2 FILLER_46_746 ();
 sg13g2_fill_2 FILLER_46_759 ();
 sg13g2_fill_1 FILLER_46_761 ();
 sg13g2_fill_2 FILLER_46_773 ();
 sg13g2_decap_4 FILLER_46_795 ();
 sg13g2_decap_4 FILLER_46_805 ();
 sg13g2_fill_2 FILLER_46_809 ();
 sg13g2_decap_4 FILLER_46_818 ();
 sg13g2_fill_2 FILLER_46_822 ();
 sg13g2_fill_2 FILLER_46_839 ();
 sg13g2_decap_8 FILLER_46_852 ();
 sg13g2_fill_2 FILLER_46_859 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_18 ();
 sg13g2_decap_8 FILLER_47_32 ();
 sg13g2_decap_8 FILLER_47_39 ();
 sg13g2_decap_4 FILLER_47_51 ();
 sg13g2_fill_1 FILLER_47_55 ();
 sg13g2_decap_4 FILLER_47_62 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_fill_2 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_94 ();
 sg13g2_decap_4 FILLER_47_101 ();
 sg13g2_fill_1 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_116 ();
 sg13g2_decap_4 FILLER_47_123 ();
 sg13g2_fill_1 FILLER_47_127 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_decap_8 FILLER_47_143 ();
 sg13g2_fill_2 FILLER_47_165 ();
 sg13g2_decap_4 FILLER_47_174 ();
 sg13g2_decap_4 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_198 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_decap_4 FILLER_47_221 ();
 sg13g2_decap_8 FILLER_47_230 ();
 sg13g2_decap_8 FILLER_47_237 ();
 sg13g2_fill_1 FILLER_47_244 ();
 sg13g2_decap_4 FILLER_47_248 ();
 sg13g2_fill_2 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_277 ();
 sg13g2_decap_8 FILLER_47_284 ();
 sg13g2_decap_8 FILLER_47_296 ();
 sg13g2_decap_4 FILLER_47_303 ();
 sg13g2_fill_2 FILLER_47_313 ();
 sg13g2_decap_8 FILLER_47_341 ();
 sg13g2_decap_8 FILLER_47_348 ();
 sg13g2_fill_2 FILLER_47_365 ();
 sg13g2_fill_1 FILLER_47_367 ();
 sg13g2_decap_8 FILLER_47_373 ();
 sg13g2_fill_2 FILLER_47_394 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_fill_1 FILLER_47_409 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_4 FILLER_47_434 ();
 sg13g2_fill_2 FILLER_47_438 ();
 sg13g2_decap_8 FILLER_47_445 ();
 sg13g2_decap_4 FILLER_47_452 ();
 sg13g2_fill_2 FILLER_47_482 ();
 sg13g2_fill_1 FILLER_47_484 ();
 sg13g2_decap_4 FILLER_47_490 ();
 sg13g2_fill_2 FILLER_47_504 ();
 sg13g2_fill_1 FILLER_47_506 ();
 sg13g2_fill_2 FILLER_47_512 ();
 sg13g2_decap_8 FILLER_47_524 ();
 sg13g2_fill_1 FILLER_47_531 ();
 sg13g2_fill_1 FILLER_47_547 ();
 sg13g2_fill_1 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_586 ();
 sg13g2_decap_4 FILLER_47_593 ();
 sg13g2_fill_2 FILLER_47_597 ();
 sg13g2_fill_2 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_631 ();
 sg13g2_decap_8 FILLER_47_638 ();
 sg13g2_decap_8 FILLER_47_645 ();
 sg13g2_decap_4 FILLER_47_663 ();
 sg13g2_fill_1 FILLER_47_667 ();
 sg13g2_decap_4 FILLER_47_675 ();
 sg13g2_fill_2 FILLER_47_679 ();
 sg13g2_fill_2 FILLER_47_701 ();
 sg13g2_fill_1 FILLER_47_703 ();
 sg13g2_decap_8 FILLER_47_709 ();
 sg13g2_fill_2 FILLER_47_716 ();
 sg13g2_decap_8 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_730 ();
 sg13g2_decap_4 FILLER_47_737 ();
 sg13g2_fill_2 FILLER_47_741 ();
 sg13g2_decap_8 FILLER_47_759 ();
 sg13g2_fill_2 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_787 ();
 sg13g2_fill_1 FILLER_47_794 ();
 sg13g2_decap_4 FILLER_47_800 ();
 sg13g2_decap_8 FILLER_47_809 ();
 sg13g2_decap_8 FILLER_47_825 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_839 ();
 sg13g2_decap_4 FILLER_47_846 ();
 sg13g2_decap_4 FILLER_47_858 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_29 ();
 sg13g2_decap_4 FILLER_48_58 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_decap_4 FILLER_48_116 ();
 sg13g2_fill_1 FILLER_48_120 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_138 ();
 sg13g2_decap_4 FILLER_48_145 ();
 sg13g2_fill_2 FILLER_48_149 ();
 sg13g2_decap_8 FILLER_48_159 ();
 sg13g2_decap_8 FILLER_48_166 ();
 sg13g2_fill_2 FILLER_48_173 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_4 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_222 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_251 ();
 sg13g2_fill_1 FILLER_48_253 ();
 sg13g2_fill_2 FILLER_48_265 ();
 sg13g2_fill_2 FILLER_48_280 ();
 sg13g2_fill_1 FILLER_48_282 ();
 sg13g2_decap_4 FILLER_48_296 ();
 sg13g2_fill_2 FILLER_48_308 ();
 sg13g2_fill_1 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_328 ();
 sg13g2_decap_8 FILLER_48_335 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_48_370 ();
 sg13g2_decap_4 FILLER_48_381 ();
 sg13g2_fill_1 FILLER_48_385 ();
 sg13g2_fill_2 FILLER_48_391 ();
 sg13g2_fill_1 FILLER_48_393 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_4 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_4 FILLER_48_434 ();
 sg13g2_fill_1 FILLER_48_438 ();
 sg13g2_decap_4 FILLER_48_454 ();
 sg13g2_fill_1 FILLER_48_458 ();
 sg13g2_decap_8 FILLER_48_464 ();
 sg13g2_decap_4 FILLER_48_471 ();
 sg13g2_fill_1 FILLER_48_475 ();
 sg13g2_fill_2 FILLER_48_481 ();
 sg13g2_decap_8 FILLER_48_491 ();
 sg13g2_decap_8 FILLER_48_498 ();
 sg13g2_fill_1 FILLER_48_505 ();
 sg13g2_fill_2 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_523 ();
 sg13g2_fill_2 FILLER_48_530 ();
 sg13g2_fill_1 FILLER_48_532 ();
 sg13g2_decap_4 FILLER_48_540 ();
 sg13g2_fill_1 FILLER_48_544 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_4 FILLER_48_560 ();
 sg13g2_fill_1 FILLER_48_564 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_583 ();
 sg13g2_decap_4 FILLER_48_600 ();
 sg13g2_fill_2 FILLER_48_604 ();
 sg13g2_decap_8 FILLER_48_611 ();
 sg13g2_decap_8 FILLER_48_618 ();
 sg13g2_fill_2 FILLER_48_630 ();
 sg13g2_fill_1 FILLER_48_632 ();
 sg13g2_decap_8 FILLER_48_638 ();
 sg13g2_fill_1 FILLER_48_645 ();
 sg13g2_decap_4 FILLER_48_661 ();
 sg13g2_fill_1 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_676 ();
 sg13g2_fill_2 FILLER_48_683 ();
 sg13g2_fill_1 FILLER_48_685 ();
 sg13g2_decap_8 FILLER_48_691 ();
 sg13g2_decap_4 FILLER_48_698 ();
 sg13g2_fill_2 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_713 ();
 sg13g2_fill_2 FILLER_48_720 ();
 sg13g2_fill_1 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_781 ();
 sg13g2_fill_2 FILLER_48_788 ();
 sg13g2_decap_4 FILLER_48_799 ();
 sg13g2_fill_2 FILLER_48_813 ();
 sg13g2_fill_1 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_821 ();
 sg13g2_decap_8 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_846 ();
 sg13g2_decap_8 FILLER_48_853 ();
 sg13g2_fill_2 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_34 ();
 sg13g2_decap_8 FILLER_49_41 ();
 sg13g2_decap_8 FILLER_49_48 ();
 sg13g2_decap_8 FILLER_49_55 ();
 sg13g2_fill_1 FILLER_49_62 ();
 sg13g2_decap_8 FILLER_49_73 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_fill_1 FILLER_49_82 ();
 sg13g2_decap_8 FILLER_49_87 ();
 sg13g2_decap_8 FILLER_49_94 ();
 sg13g2_decap_8 FILLER_49_101 ();
 sg13g2_fill_2 FILLER_49_108 ();
 sg13g2_decap_4 FILLER_49_114 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_fill_1 FILLER_49_129 ();
 sg13g2_decap_4 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_162 ();
 sg13g2_decap_8 FILLER_49_169 ();
 sg13g2_fill_2 FILLER_49_176 ();
 sg13g2_fill_1 FILLER_49_178 ();
 sg13g2_decap_8 FILLER_49_194 ();
 sg13g2_decap_4 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_232 ();
 sg13g2_decap_8 FILLER_49_239 ();
 sg13g2_decap_4 FILLER_49_246 ();
 sg13g2_fill_1 FILLER_49_250 ();
 sg13g2_decap_8 FILLER_49_265 ();
 sg13g2_decap_4 FILLER_49_272 ();
 sg13g2_fill_1 FILLER_49_276 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_decap_8 FILLER_49_288 ();
 sg13g2_decap_8 FILLER_49_295 ();
 sg13g2_decap_8 FILLER_49_302 ();
 sg13g2_decap_8 FILLER_49_309 ();
 sg13g2_decap_8 FILLER_49_316 ();
 sg13g2_fill_2 FILLER_49_323 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_4 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_decap_4 FILLER_49_366 ();
 sg13g2_fill_2 FILLER_49_370 ();
 sg13g2_fill_2 FILLER_49_387 ();
 sg13g2_fill_1 FILLER_49_389 ();
 sg13g2_fill_2 FILLER_49_404 ();
 sg13g2_decap_4 FILLER_49_419 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_fill_1 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_470 ();
 sg13g2_decap_8 FILLER_49_477 ();
 sg13g2_decap_4 FILLER_49_484 ();
 sg13g2_decap_8 FILLER_49_499 ();
 sg13g2_fill_1 FILLER_49_506 ();
 sg13g2_decap_8 FILLER_49_513 ();
 sg13g2_fill_2 FILLER_49_520 ();
 sg13g2_decap_8 FILLER_49_534 ();
 sg13g2_decap_8 FILLER_49_541 ();
 sg13g2_decap_8 FILLER_49_548 ();
 sg13g2_fill_1 FILLER_49_555 ();
 sg13g2_decap_4 FILLER_49_560 ();
 sg13g2_fill_1 FILLER_49_564 ();
 sg13g2_fill_2 FILLER_49_571 ();
 sg13g2_fill_1 FILLER_49_573 ();
 sg13g2_decap_4 FILLER_49_586 ();
 sg13g2_fill_2 FILLER_49_590 ();
 sg13g2_decap_8 FILLER_49_611 ();
 sg13g2_decap_4 FILLER_49_618 ();
 sg13g2_fill_1 FILLER_49_622 ();
 sg13g2_decap_4 FILLER_49_633 ();
 sg13g2_fill_2 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_4 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_4 FILLER_49_672 ();
 sg13g2_decap_4 FILLER_49_684 ();
 sg13g2_fill_1 FILLER_49_688 ();
 sg13g2_fill_1 FILLER_49_698 ();
 sg13g2_fill_2 FILLER_49_704 ();
 sg13g2_decap_8 FILLER_49_717 ();
 sg13g2_fill_2 FILLER_49_724 ();
 sg13g2_decap_4 FILLER_49_743 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_fill_2 FILLER_49_770 ();
 sg13g2_fill_1 FILLER_49_811 ();
 sg13g2_decap_8 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_4 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_18 ();
 sg13g2_fill_2 FILLER_50_32 ();
 sg13g2_fill_1 FILLER_50_34 ();
 sg13g2_decap_8 FILLER_50_43 ();
 sg13g2_decap_8 FILLER_50_50 ();
 sg13g2_decap_4 FILLER_50_57 ();
 sg13g2_fill_2 FILLER_50_61 ();
 sg13g2_fill_2 FILLER_50_68 ();
 sg13g2_decap_4 FILLER_50_76 ();
 sg13g2_fill_1 FILLER_50_80 ();
 sg13g2_decap_4 FILLER_50_96 ();
 sg13g2_fill_1 FILLER_50_100 ();
 sg13g2_fill_2 FILLER_50_107 ();
 sg13g2_fill_1 FILLER_50_109 ();
 sg13g2_fill_2 FILLER_50_120 ();
 sg13g2_decap_8 FILLER_50_129 ();
 sg13g2_decap_4 FILLER_50_136 ();
 sg13g2_decap_4 FILLER_50_145 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_decap_4 FILLER_50_164 ();
 sg13g2_fill_2 FILLER_50_181 ();
 sg13g2_decap_8 FILLER_50_192 ();
 sg13g2_fill_2 FILLER_50_199 ();
 sg13g2_fill_1 FILLER_50_201 ();
 sg13g2_decap_8 FILLER_50_219 ();
 sg13g2_decap_4 FILLER_50_226 ();
 sg13g2_fill_1 FILLER_50_230 ();
 sg13g2_decap_8 FILLER_50_247 ();
 sg13g2_decap_4 FILLER_50_254 ();
 sg13g2_fill_1 FILLER_50_258 ();
 sg13g2_fill_2 FILLER_50_264 ();
 sg13g2_fill_1 FILLER_50_291 ();
 sg13g2_decap_4 FILLER_50_310 ();
 sg13g2_fill_2 FILLER_50_314 ();
 sg13g2_decap_8 FILLER_50_321 ();
 sg13g2_decap_8 FILLER_50_328 ();
 sg13g2_decap_8 FILLER_50_335 ();
 sg13g2_decap_4 FILLER_50_342 ();
 sg13g2_fill_2 FILLER_50_346 ();
 sg13g2_decap_8 FILLER_50_375 ();
 sg13g2_decap_8 FILLER_50_382 ();
 sg13g2_decap_8 FILLER_50_389 ();
 sg13g2_decap_8 FILLER_50_396 ();
 sg13g2_decap_8 FILLER_50_403 ();
 sg13g2_decap_8 FILLER_50_416 ();
 sg13g2_decap_8 FILLER_50_423 ();
 sg13g2_decap_4 FILLER_50_430 ();
 sg13g2_fill_1 FILLER_50_434 ();
 sg13g2_decap_8 FILLER_50_445 ();
 sg13g2_decap_8 FILLER_50_452 ();
 sg13g2_fill_1 FILLER_50_459 ();
 sg13g2_fill_1 FILLER_50_477 ();
 sg13g2_decap_8 FILLER_50_491 ();
 sg13g2_decap_4 FILLER_50_498 ();
 sg13g2_fill_2 FILLER_50_502 ();
 sg13g2_decap_8 FILLER_50_514 ();
 sg13g2_fill_2 FILLER_50_521 ();
 sg13g2_fill_1 FILLER_50_523 ();
 sg13g2_fill_1 FILLER_50_541 ();
 sg13g2_decap_4 FILLER_50_547 ();
 sg13g2_decap_8 FILLER_50_566 ();
 sg13g2_decap_8 FILLER_50_573 ();
 sg13g2_decap_8 FILLER_50_580 ();
 sg13g2_decap_8 FILLER_50_587 ();
 sg13g2_fill_1 FILLER_50_594 ();
 sg13g2_decap_4 FILLER_50_613 ();
 sg13g2_fill_2 FILLER_50_617 ();
 sg13g2_decap_8 FILLER_50_640 ();
 sg13g2_decap_8 FILLER_50_647 ();
 sg13g2_decap_8 FILLER_50_659 ();
 sg13g2_decap_8 FILLER_50_666 ();
 sg13g2_decap_8 FILLER_50_687 ();
 sg13g2_decap_8 FILLER_50_694 ();
 sg13g2_decap_8 FILLER_50_701 ();
 sg13g2_decap_8 FILLER_50_708 ();
 sg13g2_decap_4 FILLER_50_715 ();
 sg13g2_fill_2 FILLER_50_724 ();
 sg13g2_fill_2 FILLER_50_734 ();
 sg13g2_fill_1 FILLER_50_736 ();
 sg13g2_decap_8 FILLER_50_742 ();
 sg13g2_decap_4 FILLER_50_749 ();
 sg13g2_fill_1 FILLER_50_753 ();
 sg13g2_fill_2 FILLER_50_759 ();
 sg13g2_decap_8 FILLER_50_771 ();
 sg13g2_decap_8 FILLER_50_778 ();
 sg13g2_decap_8 FILLER_50_785 ();
 sg13g2_decap_8 FILLER_50_792 ();
 sg13g2_decap_8 FILLER_50_799 ();
 sg13g2_decap_4 FILLER_50_806 ();
 sg13g2_fill_2 FILLER_50_810 ();
 sg13g2_decap_8 FILLER_50_817 ();
 sg13g2_decap_8 FILLER_50_824 ();
 sg13g2_decap_8 FILLER_50_831 ();
 sg13g2_decap_8 FILLER_50_838 ();
 sg13g2_decap_8 FILLER_50_845 ();
 sg13g2_decap_8 FILLER_50_852 ();
 sg13g2_fill_2 FILLER_50_859 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_4 FILLER_51_35 ();
 sg13g2_fill_1 FILLER_51_39 ();
 sg13g2_fill_2 FILLER_51_80 ();
 sg13g2_fill_1 FILLER_51_87 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_136 ();
 sg13g2_fill_2 FILLER_51_143 ();
 sg13g2_decap_4 FILLER_51_150 ();
 sg13g2_decap_8 FILLER_51_158 ();
 sg13g2_decap_8 FILLER_51_165 ();
 sg13g2_decap_8 FILLER_51_172 ();
 sg13g2_fill_2 FILLER_51_179 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_decap_8 FILLER_51_186 ();
 sg13g2_decap_8 FILLER_51_193 ();
 sg13g2_decap_4 FILLER_51_200 ();
 sg13g2_fill_2 FILLER_51_204 ();
 sg13g2_decap_4 FILLER_51_229 ();
 sg13g2_fill_2 FILLER_51_233 ();
 sg13g2_decap_8 FILLER_51_258 ();
 sg13g2_decap_4 FILLER_51_265 ();
 sg13g2_decap_8 FILLER_51_274 ();
 sg13g2_decap_8 FILLER_51_281 ();
 sg13g2_decap_8 FILLER_51_288 ();
 sg13g2_fill_2 FILLER_51_295 ();
 sg13g2_decap_8 FILLER_51_305 ();
 sg13g2_decap_8 FILLER_51_312 ();
 sg13g2_decap_4 FILLER_51_339 ();
 sg13g2_decap_8 FILLER_51_355 ();
 sg13g2_decap_8 FILLER_51_362 ();
 sg13g2_decap_4 FILLER_51_369 ();
 sg13g2_fill_1 FILLER_51_373 ();
 sg13g2_fill_1 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_388 ();
 sg13g2_decap_8 FILLER_51_395 ();
 sg13g2_fill_1 FILLER_51_402 ();
 sg13g2_fill_2 FILLER_51_416 ();
 sg13g2_fill_1 FILLER_51_418 ();
 sg13g2_decap_4 FILLER_51_424 ();
 sg13g2_fill_1 FILLER_51_428 ();
 sg13g2_fill_2 FILLER_51_443 ();
 sg13g2_fill_1 FILLER_51_445 ();
 sg13g2_fill_2 FILLER_51_454 ();
 sg13g2_decap_8 FILLER_51_464 ();
 sg13g2_fill_1 FILLER_51_471 ();
 sg13g2_fill_1 FILLER_51_476 ();
 sg13g2_decap_4 FILLER_51_482 ();
 sg13g2_decap_8 FILLER_51_492 ();
 sg13g2_decap_8 FILLER_51_516 ();
 sg13g2_fill_2 FILLER_51_523 ();
 sg13g2_decap_4 FILLER_51_542 ();
 sg13g2_fill_2 FILLER_51_557 ();
 sg13g2_fill_1 FILLER_51_559 ();
 sg13g2_fill_1 FILLER_51_573 ();
 sg13g2_decap_8 FILLER_51_579 ();
 sg13g2_decap_8 FILLER_51_586 ();
 sg13g2_fill_1 FILLER_51_593 ();
 sg13g2_fill_2 FILLER_51_598 ();
 sg13g2_fill_1 FILLER_51_600 ();
 sg13g2_decap_8 FILLER_51_606 ();
 sg13g2_decap_8 FILLER_51_613 ();
 sg13g2_decap_4 FILLER_51_620 ();
 sg13g2_decap_4 FILLER_51_636 ();
 sg13g2_fill_1 FILLER_51_640 ();
 sg13g2_fill_2 FILLER_51_667 ();
 sg13g2_fill_1 FILLER_51_669 ();
 sg13g2_decap_8 FILLER_51_676 ();
 sg13g2_decap_8 FILLER_51_690 ();
 sg13g2_decap_4 FILLER_51_697 ();
 sg13g2_decap_4 FILLER_51_711 ();
 sg13g2_fill_2 FILLER_51_731 ();
 sg13g2_fill_1 FILLER_51_733 ();
 sg13g2_decap_8 FILLER_51_747 ();
 sg13g2_decap_8 FILLER_51_754 ();
 sg13g2_decap_8 FILLER_51_761 ();
 sg13g2_decap_4 FILLER_51_768 ();
 sg13g2_fill_2 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_8 FILLER_51_804 ();
 sg13g2_decap_4 FILLER_51_811 ();
 sg13g2_fill_1 FILLER_51_815 ();
 sg13g2_decap_8 FILLER_51_820 ();
 sg13g2_decap_8 FILLER_51_835 ();
 sg13g2_decap_8 FILLER_51_842 ();
 sg13g2_decap_8 FILLER_51_849 ();
 sg13g2_decap_4 FILLER_51_856 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_4 FILLER_52_49 ();
 sg13g2_fill_2 FILLER_52_53 ();
 sg13g2_decap_4 FILLER_52_59 ();
 sg13g2_decap_4 FILLER_52_67 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_decap_8 FILLER_52_87 ();
 sg13g2_fill_2 FILLER_52_94 ();
 sg13g2_fill_1 FILLER_52_96 ();
 sg13g2_decap_8 FILLER_52_115 ();
 sg13g2_fill_2 FILLER_52_132 ();
 sg13g2_fill_2 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_147 ();
 sg13g2_fill_2 FILLER_52_188 ();
 sg13g2_fill_1 FILLER_52_190 ();
 sg13g2_decap_8 FILLER_52_204 ();
 sg13g2_fill_2 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_213 ();
 sg13g2_decap_8 FILLER_52_230 ();
 sg13g2_decap_4 FILLER_52_237 ();
 sg13g2_decap_8 FILLER_52_246 ();
 sg13g2_decap_8 FILLER_52_253 ();
 sg13g2_decap_4 FILLER_52_260 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_2 FILLER_52_272 ();
 sg13g2_fill_1 FILLER_52_274 ();
 sg13g2_decap_8 FILLER_52_285 ();
 sg13g2_fill_1 FILLER_52_292 ();
 sg13g2_fill_2 FILLER_52_303 ();
 sg13g2_decap_4 FILLER_52_322 ();
 sg13g2_fill_1 FILLER_52_326 ();
 sg13g2_decap_8 FILLER_52_332 ();
 sg13g2_fill_2 FILLER_52_339 ();
 sg13g2_decap_4 FILLER_52_346 ();
 sg13g2_fill_2 FILLER_52_350 ();
 sg13g2_decap_4 FILLER_52_365 ();
 sg13g2_fill_2 FILLER_52_369 ();
 sg13g2_decap_4 FILLER_52_388 ();
 sg13g2_decap_4 FILLER_52_409 ();
 sg13g2_decap_8 FILLER_52_417 ();
 sg13g2_fill_1 FILLER_52_424 ();
 sg13g2_decap_8 FILLER_52_431 ();
 sg13g2_decap_4 FILLER_52_438 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_fill_2 FILLER_52_467 ();
 sg13g2_fill_1 FILLER_52_469 ();
 sg13g2_fill_2 FILLER_52_487 ();
 sg13g2_fill_1 FILLER_52_489 ();
 sg13g2_decap_8 FILLER_52_509 ();
 sg13g2_fill_1 FILLER_52_516 ();
 sg13g2_decap_8 FILLER_52_536 ();
 sg13g2_decap_8 FILLER_52_543 ();
 sg13g2_fill_1 FILLER_52_550 ();
 sg13g2_decap_8 FILLER_52_556 ();
 sg13g2_decap_4 FILLER_52_563 ();
 sg13g2_fill_2 FILLER_52_567 ();
 sg13g2_fill_2 FILLER_52_574 ();
 sg13g2_decap_4 FILLER_52_587 ();
 sg13g2_fill_1 FILLER_52_591 ();
 sg13g2_decap_4 FILLER_52_618 ();
 sg13g2_decap_8 FILLER_52_626 ();
 sg13g2_fill_1 FILLER_52_633 ();
 sg13g2_decap_8 FILLER_52_647 ();
 sg13g2_decap_8 FILLER_52_654 ();
 sg13g2_fill_1 FILLER_52_661 ();
 sg13g2_decap_4 FILLER_52_667 ();
 sg13g2_fill_1 FILLER_52_671 ();
 sg13g2_decap_4 FILLER_52_680 ();
 sg13g2_fill_2 FILLER_52_684 ();
 sg13g2_decap_4 FILLER_52_692 ();
 sg13g2_fill_1 FILLER_52_696 ();
 sg13g2_decap_8 FILLER_52_703 ();
 sg13g2_decap_8 FILLER_52_710 ();
 sg13g2_decap_4 FILLER_52_717 ();
 sg13g2_fill_1 FILLER_52_721 ();
 sg13g2_decap_8 FILLER_52_727 ();
 sg13g2_fill_2 FILLER_52_734 ();
 sg13g2_fill_1 FILLER_52_736 ();
 sg13g2_fill_1 FILLER_52_773 ();
 sg13g2_decap_4 FILLER_52_783 ();
 sg13g2_fill_1 FILLER_52_787 ();
 sg13g2_fill_2 FILLER_52_810 ();
 sg13g2_fill_1 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_818 ();
 sg13g2_decap_8 FILLER_52_825 ();
 sg13g2_decap_8 FILLER_52_832 ();
 sg13g2_decap_8 FILLER_52_839 ();
 sg13g2_decap_8 FILLER_52_846 ();
 sg13g2_decap_8 FILLER_52_853 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_4 FILLER_53_21 ();
 sg13g2_fill_2 FILLER_53_29 ();
 sg13g2_fill_2 FILLER_53_44 ();
 sg13g2_fill_2 FILLER_53_54 ();
 sg13g2_decap_4 FILLER_53_69 ();
 sg13g2_fill_2 FILLER_53_73 ();
 sg13g2_decap_8 FILLER_53_83 ();
 sg13g2_fill_1 FILLER_53_90 ();
 sg13g2_decap_8 FILLER_53_117 ();
 sg13g2_fill_1 FILLER_53_124 ();
 sg13g2_decap_8 FILLER_53_138 ();
 sg13g2_fill_2 FILLER_53_145 ();
 sg13g2_fill_1 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_153 ();
 sg13g2_decap_8 FILLER_53_160 ();
 sg13g2_decap_8 FILLER_53_167 ();
 sg13g2_decap_8 FILLER_53_174 ();
 sg13g2_fill_1 FILLER_53_190 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_fill_2 FILLER_53_203 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_decap_8 FILLER_53_212 ();
 sg13g2_decap_8 FILLER_53_219 ();
 sg13g2_fill_2 FILLER_53_226 ();
 sg13g2_fill_1 FILLER_53_228 ();
 sg13g2_fill_1 FILLER_53_235 ();
 sg13g2_decap_4 FILLER_53_245 ();
 sg13g2_fill_1 FILLER_53_249 ();
 sg13g2_decap_8 FILLER_53_272 ();
 sg13g2_fill_2 FILLER_53_279 ();
 sg13g2_decap_8 FILLER_53_291 ();
 sg13g2_fill_1 FILLER_53_298 ();
 sg13g2_decap_8 FILLER_53_309 ();
 sg13g2_decap_8 FILLER_53_316 ();
 sg13g2_decap_8 FILLER_53_323 ();
 sg13g2_decap_8 FILLER_53_342 ();
 sg13g2_decap_8 FILLER_53_349 ();
 sg13g2_fill_2 FILLER_53_356 ();
 sg13g2_fill_1 FILLER_53_358 ();
 sg13g2_fill_2 FILLER_53_369 ();
 sg13g2_decap_4 FILLER_53_376 ();
 sg13g2_fill_1 FILLER_53_380 ();
 sg13g2_decap_4 FILLER_53_386 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_436 ();
 sg13g2_decap_4 FILLER_53_443 ();
 sg13g2_fill_2 FILLER_53_447 ();
 sg13g2_decap_8 FILLER_53_455 ();
 sg13g2_decap_8 FILLER_53_462 ();
 sg13g2_decap_8 FILLER_53_469 ();
 sg13g2_fill_1 FILLER_53_476 ();
 sg13g2_decap_8 FILLER_53_486 ();
 sg13g2_decap_8 FILLER_53_493 ();
 sg13g2_decap_4 FILLER_53_500 ();
 sg13g2_decap_4 FILLER_53_507 ();
 sg13g2_decap_8 FILLER_53_515 ();
 sg13g2_decap_8 FILLER_53_526 ();
 sg13g2_decap_4 FILLER_53_533 ();
 sg13g2_fill_1 FILLER_53_537 ();
 sg13g2_decap_8 FILLER_53_545 ();
 sg13g2_decap_8 FILLER_53_552 ();
 sg13g2_decap_4 FILLER_53_559 ();
 sg13g2_decap_4 FILLER_53_568 ();
 sg13g2_fill_2 FILLER_53_572 ();
 sg13g2_decap_4 FILLER_53_585 ();
 sg13g2_fill_2 FILLER_53_589 ();
 sg13g2_decap_8 FILLER_53_596 ();
 sg13g2_decap_8 FILLER_53_603 ();
 sg13g2_decap_8 FILLER_53_610 ();
 sg13g2_decap_4 FILLER_53_617 ();
 sg13g2_fill_2 FILLER_53_621 ();
 sg13g2_fill_2 FILLER_53_639 ();
 sg13g2_decap_8 FILLER_53_651 ();
 sg13g2_fill_2 FILLER_53_666 ();
 sg13g2_fill_1 FILLER_53_679 ();
 sg13g2_fill_1 FILLER_53_697 ();
 sg13g2_decap_8 FILLER_53_711 ();
 sg13g2_decap_8 FILLER_53_718 ();
 sg13g2_decap_8 FILLER_53_725 ();
 sg13g2_decap_8 FILLER_53_732 ();
 sg13g2_decap_4 FILLER_53_739 ();
 sg13g2_decap_8 FILLER_53_751 ();
 sg13g2_decap_8 FILLER_53_758 ();
 sg13g2_fill_2 FILLER_53_765 ();
 sg13g2_decap_8 FILLER_53_773 ();
 sg13g2_decap_8 FILLER_53_780 ();
 sg13g2_decap_8 FILLER_53_787 ();
 sg13g2_decap_8 FILLER_53_794 ();
 sg13g2_decap_4 FILLER_53_801 ();
 sg13g2_decap_8 FILLER_53_813 ();
 sg13g2_decap_8 FILLER_53_820 ();
 sg13g2_decap_8 FILLER_53_827 ();
 sg13g2_decap_8 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_841 ();
 sg13g2_decap_8 FILLER_53_848 ();
 sg13g2_decap_8 FILLER_53_855 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_4 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_46 ();
 sg13g2_decap_8 FILLER_54_53 ();
 sg13g2_decap_8 FILLER_54_60 ();
 sg13g2_decap_8 FILLER_54_83 ();
 sg13g2_decap_8 FILLER_54_90 ();
 sg13g2_fill_2 FILLER_54_97 ();
 sg13g2_fill_1 FILLER_54_99 ();
 sg13g2_fill_2 FILLER_54_126 ();
 sg13g2_fill_1 FILLER_54_128 ();
 sg13g2_fill_1 FILLER_54_137 ();
 sg13g2_fill_2 FILLER_54_145 ();
 sg13g2_decap_8 FILLER_54_166 ();
 sg13g2_fill_2 FILLER_54_173 ();
 sg13g2_decap_4 FILLER_54_199 ();
 sg13g2_fill_1 FILLER_54_203 ();
 sg13g2_decap_8 FILLER_54_215 ();
 sg13g2_fill_2 FILLER_54_222 ();
 sg13g2_fill_1 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_237 ();
 sg13g2_decap_4 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_248 ();
 sg13g2_decap_8 FILLER_54_262 ();
 sg13g2_decap_8 FILLER_54_269 ();
 sg13g2_decap_8 FILLER_54_276 ();
 sg13g2_decap_8 FILLER_54_283 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_decap_8 FILLER_54_304 ();
 sg13g2_decap_4 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_315 ();
 sg13g2_decap_8 FILLER_54_323 ();
 sg13g2_decap_4 FILLER_54_330 ();
 sg13g2_fill_1 FILLER_54_334 ();
 sg13g2_decap_8 FILLER_54_351 ();
 sg13g2_decap_4 FILLER_54_358 ();
 sg13g2_fill_1 FILLER_54_362 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_fill_2 FILLER_54_385 ();
 sg13g2_fill_1 FILLER_54_387 ();
 sg13g2_fill_1 FILLER_54_393 ();
 sg13g2_decap_8 FILLER_54_404 ();
 sg13g2_decap_8 FILLER_54_411 ();
 sg13g2_decap_8 FILLER_54_418 ();
 sg13g2_decap_8 FILLER_54_425 ();
 sg13g2_decap_8 FILLER_54_432 ();
 sg13g2_fill_1 FILLER_54_439 ();
 sg13g2_fill_1 FILLER_54_466 ();
 sg13g2_decap_4 FILLER_54_487 ();
 sg13g2_fill_2 FILLER_54_491 ();
 sg13g2_fill_1 FILLER_54_537 ();
 sg13g2_fill_2 FILLER_54_563 ();
 sg13g2_fill_1 FILLER_54_565 ();
 sg13g2_decap_8 FILLER_54_586 ();
 sg13g2_fill_2 FILLER_54_603 ();
 sg13g2_decap_4 FILLER_54_621 ();
 sg13g2_fill_1 FILLER_54_625 ();
 sg13g2_decap_8 FILLER_54_631 ();
 sg13g2_fill_2 FILLER_54_638 ();
 sg13g2_fill_1 FILLER_54_640 ();
 sg13g2_decap_4 FILLER_54_659 ();
 sg13g2_decap_4 FILLER_54_669 ();
 sg13g2_fill_2 FILLER_54_673 ();
 sg13g2_decap_4 FILLER_54_680 ();
 sg13g2_fill_2 FILLER_54_692 ();
 sg13g2_fill_1 FILLER_54_694 ();
 sg13g2_decap_8 FILLER_54_701 ();
 sg13g2_fill_2 FILLER_54_708 ();
 sg13g2_fill_1 FILLER_54_710 ();
 sg13g2_decap_4 FILLER_54_716 ();
 sg13g2_decap_8 FILLER_54_736 ();
 sg13g2_decap_4 FILLER_54_743 ();
 sg13g2_fill_1 FILLER_54_747 ();
 sg13g2_decap_8 FILLER_54_754 ();
 sg13g2_fill_1 FILLER_54_766 ();
 sg13g2_decap_8 FILLER_54_772 ();
 sg13g2_decap_8 FILLER_54_787 ();
 sg13g2_decap_8 FILLER_54_794 ();
 sg13g2_decap_8 FILLER_54_801 ();
 sg13g2_decap_8 FILLER_54_808 ();
 sg13g2_decap_8 FILLER_54_815 ();
 sg13g2_decap_8 FILLER_54_822 ();
 sg13g2_decap_8 FILLER_54_829 ();
 sg13g2_decap_8 FILLER_54_836 ();
 sg13g2_decap_8 FILLER_54_843 ();
 sg13g2_decap_8 FILLER_54_850 ();
 sg13g2_decap_4 FILLER_54_857 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_36 ();
 sg13g2_decap_8 FILLER_55_43 ();
 sg13g2_decap_8 FILLER_55_50 ();
 sg13g2_decap_8 FILLER_55_57 ();
 sg13g2_decap_8 FILLER_55_64 ();
 sg13g2_decap_8 FILLER_55_71 ();
 sg13g2_decap_8 FILLER_55_78 ();
 sg13g2_decap_8 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_92 ();
 sg13g2_decap_8 FILLER_55_107 ();
 sg13g2_decap_8 FILLER_55_114 ();
 sg13g2_decap_8 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_128 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_2 FILLER_55_153 ();
 sg13g2_fill_1 FILLER_55_155 ();
 sg13g2_fill_1 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_171 ();
 sg13g2_decap_8 FILLER_55_183 ();
 sg13g2_decap_8 FILLER_55_190 ();
 sg13g2_decap_8 FILLER_55_197 ();
 sg13g2_decap_4 FILLER_55_204 ();
 sg13g2_decap_8 FILLER_55_218 ();
 sg13g2_fill_1 FILLER_55_225 ();
 sg13g2_decap_8 FILLER_55_243 ();
 sg13g2_decap_8 FILLER_55_250 ();
 sg13g2_fill_2 FILLER_55_257 ();
 sg13g2_fill_1 FILLER_55_275 ();
 sg13g2_fill_2 FILLER_55_294 ();
 sg13g2_fill_1 FILLER_55_296 ();
 sg13g2_fill_1 FILLER_55_315 ();
 sg13g2_decap_8 FILLER_55_340 ();
 sg13g2_decap_4 FILLER_55_355 ();
 sg13g2_fill_2 FILLER_55_359 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_4 FILLER_55_378 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_decap_8 FILLER_55_388 ();
 sg13g2_decap_8 FILLER_55_395 ();
 sg13g2_decap_4 FILLER_55_402 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_2 FILLER_55_416 ();
 sg13g2_fill_1 FILLER_55_418 ();
 sg13g2_decap_8 FILLER_55_441 ();
 sg13g2_decap_8 FILLER_55_448 ();
 sg13g2_decap_8 FILLER_55_455 ();
 sg13g2_decap_8 FILLER_55_462 ();
 sg13g2_decap_8 FILLER_55_485 ();
 sg13g2_decap_4 FILLER_55_492 ();
 sg13g2_fill_2 FILLER_55_496 ();
 sg13g2_decap_8 FILLER_55_508 ();
 sg13g2_decap_8 FILLER_55_515 ();
 sg13g2_decap_4 FILLER_55_522 ();
 sg13g2_decap_8 FILLER_55_533 ();
 sg13g2_decap_4 FILLER_55_540 ();
 sg13g2_fill_2 FILLER_55_544 ();
 sg13g2_decap_8 FILLER_55_556 ();
 sg13g2_decap_4 FILLER_55_563 ();
 sg13g2_decap_8 FILLER_55_574 ();
 sg13g2_decap_8 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_588 ();
 sg13g2_decap_8 FILLER_55_595 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_decap_8 FILLER_55_609 ();
 sg13g2_fill_1 FILLER_55_616 ();
 sg13g2_fill_2 FILLER_55_642 ();
 sg13g2_fill_1 FILLER_55_644 ();
 sg13g2_decap_8 FILLER_55_659 ();
 sg13g2_decap_8 FILLER_55_666 ();
 sg13g2_fill_1 FILLER_55_684 ();
 sg13g2_decap_8 FILLER_55_692 ();
 sg13g2_decap_8 FILLER_55_704 ();
 sg13g2_fill_1 FILLER_55_711 ();
 sg13g2_decap_8 FILLER_55_724 ();
 sg13g2_fill_2 FILLER_55_731 ();
 sg13g2_fill_1 FILLER_55_733 ();
 sg13g2_decap_4 FILLER_55_747 ();
 sg13g2_fill_1 FILLER_55_751 ();
 sg13g2_fill_2 FILLER_55_760 ();
 sg13g2_fill_1 FILLER_55_762 ();
 sg13g2_decap_8 FILLER_55_771 ();
 sg13g2_decap_8 FILLER_55_778 ();
 sg13g2_decap_8 FILLER_55_785 ();
 sg13g2_decap_8 FILLER_55_792 ();
 sg13g2_decap_8 FILLER_55_799 ();
 sg13g2_decap_8 FILLER_55_806 ();
 sg13g2_decap_8 FILLER_55_813 ();
 sg13g2_decap_8 FILLER_55_820 ();
 sg13g2_decap_8 FILLER_55_827 ();
 sg13g2_decap_8 FILLER_55_834 ();
 sg13g2_decap_8 FILLER_55_841 ();
 sg13g2_decap_8 FILLER_55_848 ();
 sg13g2_decap_8 FILLER_55_855 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_4 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_82 ();
 sg13g2_decap_8 FILLER_56_89 ();
 sg13g2_decap_8 FILLER_56_96 ();
 sg13g2_decap_8 FILLER_56_111 ();
 sg13g2_decap_8 FILLER_56_118 ();
 sg13g2_fill_1 FILLER_56_125 ();
 sg13g2_decap_8 FILLER_56_134 ();
 sg13g2_fill_2 FILLER_56_141 ();
 sg13g2_fill_1 FILLER_56_143 ();
 sg13g2_decap_8 FILLER_56_149 ();
 sg13g2_decap_4 FILLER_56_156 ();
 sg13g2_decap_8 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_178 ();
 sg13g2_fill_1 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_185 ();
 sg13g2_decap_8 FILLER_56_193 ();
 sg13g2_decap_8 FILLER_56_200 ();
 sg13g2_decap_4 FILLER_56_207 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_fill_1 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_decap_4 FILLER_56_245 ();
 sg13g2_fill_1 FILLER_56_274 ();
 sg13g2_decap_4 FILLER_56_285 ();
 sg13g2_fill_1 FILLER_56_289 ();
 sg13g2_decap_4 FILLER_56_294 ();
 sg13g2_fill_1 FILLER_56_298 ();
 sg13g2_decap_8 FILLER_56_303 ();
 sg13g2_decap_8 FILLER_56_310 ();
 sg13g2_decap_8 FILLER_56_317 ();
 sg13g2_decap_8 FILLER_56_329 ();
 sg13g2_fill_2 FILLER_56_336 ();
 sg13g2_fill_1 FILLER_56_338 ();
 sg13g2_decap_8 FILLER_56_347 ();
 sg13g2_fill_2 FILLER_56_354 ();
 sg13g2_fill_1 FILLER_56_356 ();
 sg13g2_decap_8 FILLER_56_365 ();
 sg13g2_fill_2 FILLER_56_372 ();
 sg13g2_decap_4 FILLER_56_393 ();
 sg13g2_fill_1 FILLER_56_413 ();
 sg13g2_decap_8 FILLER_56_422 ();
 sg13g2_decap_8 FILLER_56_433 ();
 sg13g2_decap_4 FILLER_56_440 ();
 sg13g2_fill_1 FILLER_56_444 ();
 sg13g2_decap_8 FILLER_56_461 ();
 sg13g2_fill_1 FILLER_56_468 ();
 sg13g2_decap_4 FILLER_56_488 ();
 sg13g2_fill_1 FILLER_56_503 ();
 sg13g2_decap_8 FILLER_56_515 ();
 sg13g2_fill_2 FILLER_56_522 ();
 sg13g2_decap_4 FILLER_56_532 ();
 sg13g2_fill_1 FILLER_56_536 ();
 sg13g2_decap_8 FILLER_56_552 ();
 sg13g2_fill_2 FILLER_56_559 ();
 sg13g2_fill_1 FILLER_56_569 ();
 sg13g2_fill_2 FILLER_56_587 ();
 sg13g2_decap_8 FILLER_56_637 ();
 sg13g2_fill_2 FILLER_56_644 ();
 sg13g2_fill_1 FILLER_56_646 ();
 sg13g2_decap_4 FILLER_56_655 ();
 sg13g2_fill_1 FILLER_56_659 ();
 sg13g2_decap_8 FILLER_56_668 ();
 sg13g2_fill_1 FILLER_56_675 ();
 sg13g2_decap_4 FILLER_56_689 ();
 sg13g2_fill_1 FILLER_56_693 ();
 sg13g2_decap_4 FILLER_56_710 ();
 sg13g2_decap_8 FILLER_56_722 ();
 sg13g2_fill_1 FILLER_56_729 ();
 sg13g2_decap_8 FILLER_56_743 ();
 sg13g2_decap_8 FILLER_56_750 ();
 sg13g2_decap_8 FILLER_56_757 ();
 sg13g2_decap_8 FILLER_56_764 ();
 sg13g2_decap_8 FILLER_56_771 ();
 sg13g2_decap_8 FILLER_56_778 ();
 sg13g2_decap_8 FILLER_56_785 ();
 sg13g2_decap_8 FILLER_56_792 ();
 sg13g2_decap_8 FILLER_56_799 ();
 sg13g2_decap_8 FILLER_56_806 ();
 sg13g2_decap_8 FILLER_56_813 ();
 sg13g2_decap_8 FILLER_56_820 ();
 sg13g2_decap_8 FILLER_56_827 ();
 sg13g2_decap_8 FILLER_56_834 ();
 sg13g2_decap_8 FILLER_56_841 ();
 sg13g2_decap_8 FILLER_56_848 ();
 sg13g2_decap_8 FILLER_56_855 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_4 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_132 ();
 sg13g2_decap_8 FILLER_57_139 ();
 sg13g2_decap_8 FILLER_57_146 ();
 sg13g2_fill_1 FILLER_57_153 ();
 sg13g2_decap_4 FILLER_57_167 ();
 sg13g2_fill_1 FILLER_57_187 ();
 sg13g2_decap_4 FILLER_57_217 ();
 sg13g2_fill_1 FILLER_57_230 ();
 sg13g2_decap_8 FILLER_57_239 ();
 sg13g2_fill_2 FILLER_57_246 ();
 sg13g2_fill_1 FILLER_57_248 ();
 sg13g2_decap_8 FILLER_57_253 ();
 sg13g2_decap_8 FILLER_57_260 ();
 sg13g2_decap_8 FILLER_57_267 ();
 sg13g2_decap_4 FILLER_57_274 ();
 sg13g2_decap_8 FILLER_57_282 ();
 sg13g2_fill_1 FILLER_57_289 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_decap_8 FILLER_57_312 ();
 sg13g2_fill_2 FILLER_57_319 ();
 sg13g2_fill_2 FILLER_57_329 ();
 sg13g2_fill_2 FILLER_57_348 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_374 ();
 sg13g2_fill_2 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_396 ();
 sg13g2_decap_8 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_57_412 ();
 sg13g2_fill_2 FILLER_57_419 ();
 sg13g2_fill_1 FILLER_57_421 ();
 sg13g2_decap_4 FILLER_57_430 ();
 sg13g2_decap_4 FILLER_57_442 ();
 sg13g2_fill_2 FILLER_57_446 ();
 sg13g2_decap_8 FILLER_57_461 ();
 sg13g2_decap_8 FILLER_57_468 ();
 sg13g2_decap_8 FILLER_57_475 ();
 sg13g2_decap_8 FILLER_57_482 ();
 sg13g2_decap_8 FILLER_57_489 ();
 sg13g2_fill_1 FILLER_57_496 ();
 sg13g2_decap_4 FILLER_57_510 ();
 sg13g2_fill_2 FILLER_57_514 ();
 sg13g2_fill_1 FILLER_57_520 ();
 sg13g2_decap_8 FILLER_57_526 ();
 sg13g2_decap_8 FILLER_57_533 ();
 sg13g2_decap_8 FILLER_57_540 ();
 sg13g2_fill_1 FILLER_57_547 ();
 sg13g2_fill_2 FILLER_57_561 ();
 sg13g2_fill_1 FILLER_57_563 ();
 sg13g2_decap_8 FILLER_57_577 ();
 sg13g2_decap_8 FILLER_57_584 ();
 sg13g2_decap_8 FILLER_57_591 ();
 sg13g2_decap_4 FILLER_57_598 ();
 sg13g2_fill_2 FILLER_57_602 ();
 sg13g2_decap_4 FILLER_57_618 ();
 sg13g2_fill_2 FILLER_57_622 ();
 sg13g2_decap_8 FILLER_57_632 ();
 sg13g2_decap_8 FILLER_57_639 ();
 sg13g2_fill_2 FILLER_57_646 ();
 sg13g2_fill_2 FILLER_57_656 ();
 sg13g2_decap_8 FILLER_57_674 ();
 sg13g2_decap_4 FILLER_57_681 ();
 sg13g2_decap_4 FILLER_57_688 ();
 sg13g2_fill_2 FILLER_57_692 ();
 sg13g2_decap_8 FILLER_57_703 ();
 sg13g2_decap_8 FILLER_57_710 ();
 sg13g2_decap_8 FILLER_57_717 ();
 sg13g2_fill_2 FILLER_57_724 ();
 sg13g2_decap_8 FILLER_57_730 ();
 sg13g2_decap_8 FILLER_57_737 ();
 sg13g2_decap_8 FILLER_57_744 ();
 sg13g2_decap_8 FILLER_57_751 ();
 sg13g2_decap_8 FILLER_57_758 ();
 sg13g2_decap_8 FILLER_57_765 ();
 sg13g2_decap_8 FILLER_57_772 ();
 sg13g2_decap_8 FILLER_57_779 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_793 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_decap_8 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_decap_8 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_842 ();
 sg13g2_decap_8 FILLER_57_849 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_fill_2 FILLER_58_210 ();
 sg13g2_fill_1 FILLER_58_212 ();
 sg13g2_fill_2 FILLER_58_245 ();
 sg13g2_fill_2 FILLER_58_281 ();
 sg13g2_decap_8 FILLER_58_291 ();
 sg13g2_fill_2 FILLER_58_298 ();
 sg13g2_fill_1 FILLER_58_300 ();
 sg13g2_fill_1 FILLER_58_314 ();
 sg13g2_decap_8 FILLER_58_323 ();
 sg13g2_decap_8 FILLER_58_330 ();
 sg13g2_decap_8 FILLER_58_337 ();
 sg13g2_decap_8 FILLER_58_344 ();
 sg13g2_decap_8 FILLER_58_351 ();
 sg13g2_decap_8 FILLER_58_358 ();
 sg13g2_fill_1 FILLER_58_365 ();
 sg13g2_decap_8 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_386 ();
 sg13g2_decap_8 FILLER_58_403 ();
 sg13g2_fill_1 FILLER_58_410 ();
 sg13g2_decap_8 FILLER_58_419 ();
 sg13g2_decap_8 FILLER_58_426 ();
 sg13g2_decap_8 FILLER_58_433 ();
 sg13g2_decap_8 FILLER_58_440 ();
 sg13g2_decap_8 FILLER_58_447 ();
 sg13g2_decap_4 FILLER_58_454 ();
 sg13g2_decap_8 FILLER_58_466 ();
 sg13g2_decap_4 FILLER_58_473 ();
 sg13g2_fill_1 FILLER_58_477 ();
 sg13g2_fill_2 FILLER_58_499 ();
 sg13g2_fill_1 FILLER_58_501 ();
 sg13g2_decap_8 FILLER_58_506 ();
 sg13g2_decap_8 FILLER_58_513 ();
 sg13g2_fill_2 FILLER_58_520 ();
 sg13g2_fill_1 FILLER_58_522 ();
 sg13g2_decap_4 FILLER_58_537 ();
 sg13g2_fill_2 FILLER_58_541 ();
 sg13g2_decap_8 FILLER_58_551 ();
 sg13g2_decap_8 FILLER_58_558 ();
 sg13g2_fill_2 FILLER_58_565 ();
 sg13g2_fill_1 FILLER_58_567 ();
 sg13g2_decap_8 FILLER_58_584 ();
 sg13g2_decap_8 FILLER_58_591 ();
 sg13g2_fill_1 FILLER_58_598 ();
 sg13g2_fill_1 FILLER_58_621 ();
 sg13g2_decap_8 FILLER_58_638 ();
 sg13g2_decap_8 FILLER_58_661 ();
 sg13g2_decap_8 FILLER_58_668 ();
 sg13g2_decap_4 FILLER_58_675 ();
 sg13g2_decap_8 FILLER_58_705 ();
 sg13g2_fill_2 FILLER_58_712 ();
 sg13g2_fill_1 FILLER_58_714 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_decap_8 FILLER_58_748 ();
 sg13g2_fill_1 FILLER_58_755 ();
 sg13g2_decap_8 FILLER_58_773 ();
 sg13g2_fill_2 FILLER_58_780 ();
 sg13g2_decap_8 FILLER_58_786 ();
 sg13g2_decap_8 FILLER_58_793 ();
 sg13g2_decap_8 FILLER_58_800 ();
 sg13g2_decap_8 FILLER_58_807 ();
 sg13g2_decap_8 FILLER_58_814 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_4 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_230 ();
 sg13g2_decap_8 FILLER_59_237 ();
 sg13g2_decap_8 FILLER_59_244 ();
 sg13g2_decap_8 FILLER_59_251 ();
 sg13g2_decap_8 FILLER_59_258 ();
 sg13g2_decap_8 FILLER_59_265 ();
 sg13g2_decap_8 FILLER_59_272 ();
 sg13g2_decap_8 FILLER_59_279 ();
 sg13g2_decap_8 FILLER_59_286 ();
 sg13g2_decap_8 FILLER_59_293 ();
 sg13g2_decap_8 FILLER_59_300 ();
 sg13g2_decap_8 FILLER_59_307 ();
 sg13g2_fill_2 FILLER_59_314 ();
 sg13g2_decap_8 FILLER_59_320 ();
 sg13g2_decap_4 FILLER_59_327 ();
 sg13g2_fill_2 FILLER_59_331 ();
 sg13g2_decap_4 FILLER_59_357 ();
 sg13g2_fill_2 FILLER_59_366 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_4 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_423 ();
 sg13g2_fill_2 FILLER_59_430 ();
 sg13g2_fill_1 FILLER_59_432 ();
 sg13g2_decap_4 FILLER_59_449 ();
 sg13g2_fill_1 FILLER_59_453 ();
 sg13g2_fill_2 FILLER_59_470 ();
 sg13g2_decap_8 FILLER_59_481 ();
 sg13g2_decap_8 FILLER_59_488 ();
 sg13g2_fill_2 FILLER_59_495 ();
 sg13g2_decap_8 FILLER_59_513 ();
 sg13g2_decap_8 FILLER_59_520 ();
 sg13g2_decap_8 FILLER_59_527 ();
 sg13g2_decap_4 FILLER_59_534 ();
 sg13g2_decap_8 FILLER_59_551 ();
 sg13g2_decap_8 FILLER_59_558 ();
 sg13g2_decap_8 FILLER_59_565 ();
 sg13g2_fill_2 FILLER_59_572 ();
 sg13g2_decap_8 FILLER_59_590 ();
 sg13g2_fill_2 FILLER_59_597 ();
 sg13g2_decap_8 FILLER_59_612 ();
 sg13g2_decap_4 FILLER_59_619 ();
 sg13g2_fill_2 FILLER_59_623 ();
 sg13g2_decap_4 FILLER_59_633 ();
 sg13g2_fill_1 FILLER_59_637 ();
 sg13g2_decap_8 FILLER_59_643 ();
 sg13g2_decap_4 FILLER_59_650 ();
 sg13g2_decap_8 FILLER_59_664 ();
 sg13g2_decap_4 FILLER_59_671 ();
 sg13g2_fill_2 FILLER_59_675 ();
 sg13g2_fill_2 FILLER_59_696 ();
 sg13g2_fill_1 FILLER_59_698 ();
 sg13g2_decap_4 FILLER_59_704 ();
 sg13g2_fill_1 FILLER_59_708 ();
 sg13g2_fill_2 FILLER_59_731 ();
 sg13g2_decap_8 FILLER_59_738 ();
 sg13g2_fill_2 FILLER_59_745 ();
 sg13g2_fill_1 FILLER_59_747 ();
 sg13g2_fill_2 FILLER_59_756 ();
 sg13g2_decap_8 FILLER_59_798 ();
 sg13g2_decap_8 FILLER_59_805 ();
 sg13g2_decap_8 FILLER_59_812 ();
 sg13g2_decap_8 FILLER_59_819 ();
 sg13g2_decap_8 FILLER_59_826 ();
 sg13g2_decap_8 FILLER_59_833 ();
 sg13g2_decap_8 FILLER_59_840 ();
 sg13g2_decap_8 FILLER_59_847 ();
 sg13g2_decap_8 FILLER_59_854 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_4 FILLER_60_301 ();
 sg13g2_fill_2 FILLER_60_335 ();
 sg13g2_decap_8 FILLER_60_345 ();
 sg13g2_decap_4 FILLER_60_352 ();
 sg13g2_fill_2 FILLER_60_356 ();
 sg13g2_decap_8 FILLER_60_366 ();
 sg13g2_fill_2 FILLER_60_373 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_decap_8 FILLER_60_389 ();
 sg13g2_decap_8 FILLER_60_396 ();
 sg13g2_fill_2 FILLER_60_403 ();
 sg13g2_decap_4 FILLER_60_409 ();
 sg13g2_fill_2 FILLER_60_413 ();
 sg13g2_decap_8 FILLER_60_431 ();
 sg13g2_decap_4 FILLER_60_438 ();
 sg13g2_decap_8 FILLER_60_446 ();
 sg13g2_decap_8 FILLER_60_453 ();
 sg13g2_decap_4 FILLER_60_460 ();
 sg13g2_fill_2 FILLER_60_472 ();
 sg13g2_fill_1 FILLER_60_474 ();
 sg13g2_decap_8 FILLER_60_483 ();
 sg13g2_decap_4 FILLER_60_490 ();
 sg13g2_fill_1 FILLER_60_502 ();
 sg13g2_decap_8 FILLER_60_522 ();
 sg13g2_fill_2 FILLER_60_529 ();
 sg13g2_fill_1 FILLER_60_539 ();
 sg13g2_decap_8 FILLER_60_556 ();
 sg13g2_fill_2 FILLER_60_563 ();
 sg13g2_decap_8 FILLER_60_581 ();
 sg13g2_decap_4 FILLER_60_588 ();
 sg13g2_decap_8 FILLER_60_607 ();
 sg13g2_decap_8 FILLER_60_614 ();
 sg13g2_decap_4 FILLER_60_621 ();
 sg13g2_fill_2 FILLER_60_625 ();
 sg13g2_fill_1 FILLER_60_640 ();
 sg13g2_decap_4 FILLER_60_645 ();
 sg13g2_fill_1 FILLER_60_649 ();
 sg13g2_fill_2 FILLER_60_658 ();
 sg13g2_decap_8 FILLER_60_673 ();
 sg13g2_decap_4 FILLER_60_680 ();
 sg13g2_decap_4 FILLER_60_711 ();
 sg13g2_fill_1 FILLER_60_715 ();
 sg13g2_decap_8 FILLER_60_733 ();
 sg13g2_decap_8 FILLER_60_744 ();
 sg13g2_decap_8 FILLER_60_751 ();
 sg13g2_fill_2 FILLER_60_762 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_decap_8 FILLER_60_781 ();
 sg13g2_decap_8 FILLER_60_788 ();
 sg13g2_decap_4 FILLER_60_795 ();
 sg13g2_fill_2 FILLER_60_799 ();
 sg13g2_decap_8 FILLER_60_827 ();
 sg13g2_decap_8 FILLER_60_834 ();
 sg13g2_decap_8 FILLER_60_841 ();
 sg13g2_decap_8 FILLER_60_848 ();
 sg13g2_decap_8 FILLER_60_855 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_266 ();
 sg13g2_decap_8 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_fill_2 FILLER_61_294 ();
 sg13g2_fill_1 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_307 ();
 sg13g2_fill_1 FILLER_61_309 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_decap_4 FILLER_61_322 ();
 sg13g2_decap_8 FILLER_61_335 ();
 sg13g2_fill_2 FILLER_61_342 ();
 sg13g2_fill_1 FILLER_61_344 ();
 sg13g2_decap_8 FILLER_61_349 ();
 sg13g2_decap_8 FILLER_61_356 ();
 sg13g2_fill_2 FILLER_61_363 ();
 sg13g2_fill_1 FILLER_61_365 ();
 sg13g2_decap_4 FILLER_61_374 ();
 sg13g2_fill_1 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_396 ();
 sg13g2_decap_8 FILLER_61_403 ();
 sg13g2_fill_1 FILLER_61_410 ();
 sg13g2_decap_8 FILLER_61_419 ();
 sg13g2_decap_4 FILLER_61_426 ();
 sg13g2_fill_1 FILLER_61_430 ();
 sg13g2_fill_2 FILLER_61_463 ();
 sg13g2_decap_8 FILLER_61_473 ();
 sg13g2_decap_4 FILLER_61_480 ();
 sg13g2_fill_2 FILLER_61_484 ();
 sg13g2_fill_2 FILLER_61_489 ();
 sg13g2_decap_8 FILLER_61_495 ();
 sg13g2_fill_2 FILLER_61_502 ();
 sg13g2_fill_1 FILLER_61_504 ();
 sg13g2_decap_4 FILLER_61_513 ();
 sg13g2_fill_2 FILLER_61_525 ();
 sg13g2_fill_1 FILLER_61_527 ();
 sg13g2_fill_1 FILLER_61_533 ();
 sg13g2_decap_8 FILLER_61_538 ();
 sg13g2_decap_4 FILLER_61_545 ();
 sg13g2_fill_1 FILLER_61_549 ();
 sg13g2_decap_8 FILLER_61_559 ();
 sg13g2_fill_1 FILLER_61_566 ();
 sg13g2_decap_8 FILLER_61_583 ();
 sg13g2_fill_1 FILLER_61_590 ();
 sg13g2_decap_8 FILLER_61_615 ();
 sg13g2_fill_2 FILLER_61_622 ();
 sg13g2_decap_8 FILLER_61_644 ();
 sg13g2_decap_4 FILLER_61_651 ();
 sg13g2_decap_8 FILLER_61_665 ();
 sg13g2_fill_2 FILLER_61_672 ();
 sg13g2_fill_1 FILLER_61_674 ();
 sg13g2_fill_1 FILLER_61_680 ();
 sg13g2_decap_8 FILLER_61_690 ();
 sg13g2_decap_8 FILLER_61_697 ();
 sg13g2_decap_4 FILLER_61_714 ();
 sg13g2_decap_8 FILLER_61_722 ();
 sg13g2_decap_4 FILLER_61_729 ();
 sg13g2_fill_2 FILLER_61_733 ();
 sg13g2_decap_8 FILLER_61_739 ();
 sg13g2_decap_8 FILLER_61_746 ();
 sg13g2_decap_8 FILLER_61_753 ();
 sg13g2_decap_8 FILLER_61_773 ();
 sg13g2_fill_2 FILLER_61_780 ();
 sg13g2_fill_1 FILLER_61_782 ();
 sg13g2_fill_1 FILLER_61_806 ();
 sg13g2_decap_8 FILLER_61_820 ();
 sg13g2_decap_8 FILLER_61_827 ();
 sg13g2_decap_8 FILLER_61_834 ();
 sg13g2_decap_8 FILLER_61_841 ();
 sg13g2_decap_8 FILLER_61_848 ();
 sg13g2_decap_8 FILLER_61_855 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_decap_4 FILLER_62_280 ();
 sg13g2_fill_1 FILLER_62_284 ();
 sg13g2_fill_1 FILLER_62_301 ();
 sg13g2_fill_2 FILLER_62_316 ();
 sg13g2_fill_2 FILLER_62_331 ();
 sg13g2_fill_1 FILLER_62_333 ();
 sg13g2_decap_8 FILLER_62_360 ();
 sg13g2_fill_2 FILLER_62_367 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_1 FILLER_62_387 ();
 sg13g2_decap_4 FILLER_62_400 ();
 sg13g2_fill_2 FILLER_62_404 ();
 sg13g2_decap_4 FILLER_62_429 ();
 sg13g2_fill_2 FILLER_62_433 ();
 sg13g2_decap_8 FILLER_62_445 ();
 sg13g2_decap_8 FILLER_62_452 ();
 sg13g2_decap_4 FILLER_62_459 ();
 sg13g2_decap_4 FILLER_62_469 ();
 sg13g2_fill_2 FILLER_62_473 ();
 sg13g2_fill_2 FILLER_62_499 ();
 sg13g2_decap_8 FILLER_62_506 ();
 sg13g2_decap_8 FILLER_62_513 ();
 sg13g2_decap_4 FILLER_62_564 ();
 sg13g2_fill_2 FILLER_62_568 ();
 sg13g2_decap_4 FILLER_62_588 ();
 sg13g2_fill_2 FILLER_62_592 ();
 sg13g2_decap_4 FILLER_62_599 ();
 sg13g2_fill_1 FILLER_62_603 ();
 sg13g2_decap_8 FILLER_62_609 ();
 sg13g2_decap_8 FILLER_62_616 ();
 sg13g2_decap_8 FILLER_62_623 ();
 sg13g2_fill_2 FILLER_62_630 ();
 sg13g2_fill_1 FILLER_62_632 ();
 sg13g2_decap_8 FILLER_62_646 ();
 sg13g2_decap_8 FILLER_62_653 ();
 sg13g2_decap_4 FILLER_62_660 ();
 sg13g2_fill_2 FILLER_62_664 ();
 sg13g2_decap_8 FILLER_62_697 ();
 sg13g2_fill_1 FILLER_62_704 ();
 sg13g2_fill_1 FILLER_62_717 ();
 sg13g2_decap_8 FILLER_62_797 ();
 sg13g2_decap_8 FILLER_62_804 ();
 sg13g2_decap_8 FILLER_62_811 ();
 sg13g2_decap_8 FILLER_62_818 ();
 sg13g2_decap_8 FILLER_62_825 ();
 sg13g2_decap_8 FILLER_62_832 ();
 sg13g2_decap_8 FILLER_62_839 ();
 sg13g2_decap_8 FILLER_62_846 ();
 sg13g2_decap_8 FILLER_62_853 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_fill_1 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_309 ();
 sg13g2_decap_8 FILLER_63_316 ();
 sg13g2_decap_8 FILLER_63_323 ();
 sg13g2_decap_8 FILLER_63_330 ();
 sg13g2_decap_4 FILLER_63_337 ();
 sg13g2_fill_1 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_368 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_63_409 ();
 sg13g2_decap_8 FILLER_63_425 ();
 sg13g2_decap_8 FILLER_63_432 ();
 sg13g2_fill_2 FILLER_63_439 ();
 sg13g2_decap_8 FILLER_63_481 ();
 sg13g2_decap_8 FILLER_63_488 ();
 sg13g2_fill_2 FILLER_63_499 ();
 sg13g2_decap_4 FILLER_63_513 ();
 sg13g2_fill_1 FILLER_63_517 ();
 sg13g2_fill_2 FILLER_63_526 ();
 sg13g2_fill_1 FILLER_63_528 ();
 sg13g2_decap_4 FILLER_63_543 ();
 sg13g2_fill_2 FILLER_63_547 ();
 sg13g2_decap_8 FILLER_63_553 ();
 sg13g2_decap_8 FILLER_63_560 ();
 sg13g2_decap_8 FILLER_63_567 ();
 sg13g2_decap_8 FILLER_63_582 ();
 sg13g2_decap_8 FILLER_63_589 ();
 sg13g2_decap_4 FILLER_63_596 ();
 sg13g2_fill_2 FILLER_63_600 ();
 sg13g2_decap_8 FILLER_63_628 ();
 sg13g2_fill_1 FILLER_63_635 ();
 sg13g2_fill_1 FILLER_63_667 ();
 sg13g2_fill_2 FILLER_63_676 ();
 sg13g2_decap_4 FILLER_63_690 ();
 sg13g2_fill_2 FILLER_63_694 ();
 sg13g2_fill_2 FILLER_63_700 ();
 sg13g2_fill_1 FILLER_63_702 ();
 sg13g2_decap_8 FILLER_63_709 ();
 sg13g2_decap_8 FILLER_63_716 ();
 sg13g2_decap_8 FILLER_63_728 ();
 sg13g2_decap_8 FILLER_63_735 ();
 sg13g2_decap_4 FILLER_63_742 ();
 sg13g2_decap_4 FILLER_63_778 ();
 sg13g2_fill_2 FILLER_63_782 ();
 sg13g2_decap_4 FILLER_63_789 ();
 sg13g2_fill_1 FILLER_63_793 ();
 sg13g2_decap_8 FILLER_63_802 ();
 sg13g2_decap_8 FILLER_63_809 ();
 sg13g2_decap_8 FILLER_63_816 ();
 sg13g2_decap_8 FILLER_63_823 ();
 sg13g2_decap_8 FILLER_63_830 ();
 sg13g2_decap_8 FILLER_63_837 ();
 sg13g2_decap_8 FILLER_63_844 ();
 sg13g2_decap_8 FILLER_63_851 ();
 sg13g2_decap_4 FILLER_63_858 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_fill_2 FILLER_64_280 ();
 sg13g2_fill_1 FILLER_64_282 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_fill_2 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_fill_2 FILLER_64_350 ();
 sg13g2_fill_1 FILLER_64_352 ();
 sg13g2_decap_4 FILLER_64_357 ();
 sg13g2_decap_4 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_378 ();
 sg13g2_decap_8 FILLER_64_384 ();
 sg13g2_decap_4 FILLER_64_391 ();
 sg13g2_fill_1 FILLER_64_395 ();
 sg13g2_decap_8 FILLER_64_409 ();
 sg13g2_decap_8 FILLER_64_416 ();
 sg13g2_decap_8 FILLER_64_423 ();
 sg13g2_decap_4 FILLER_64_434 ();
 sg13g2_fill_2 FILLER_64_438 ();
 sg13g2_decap_8 FILLER_64_448 ();
 sg13g2_decap_8 FILLER_64_455 ();
 sg13g2_fill_2 FILLER_64_462 ();
 sg13g2_fill_1 FILLER_64_464 ();
 sg13g2_fill_2 FILLER_64_479 ();
 sg13g2_fill_1 FILLER_64_481 ();
 sg13g2_decap_4 FILLER_64_485 ();
 sg13g2_decap_8 FILLER_64_509 ();
 sg13g2_decap_4 FILLER_64_516 ();
 sg13g2_fill_1 FILLER_64_524 ();
 sg13g2_decap_8 FILLER_64_529 ();
 sg13g2_decap_8 FILLER_64_536 ();
 sg13g2_decap_8 FILLER_64_543 ();
 sg13g2_decap_4 FILLER_64_550 ();
 sg13g2_fill_2 FILLER_64_554 ();
 sg13g2_decap_8 FILLER_64_566 ();
 sg13g2_fill_1 FILLER_64_573 ();
 sg13g2_decap_8 FILLER_64_589 ();
 sg13g2_decap_4 FILLER_64_596 ();
 sg13g2_fill_1 FILLER_64_600 ();
 sg13g2_decap_4 FILLER_64_605 ();
 sg13g2_fill_2 FILLER_64_609 ();
 sg13g2_fill_2 FILLER_64_624 ();
 sg13g2_fill_1 FILLER_64_626 ();
 sg13g2_decap_8 FILLER_64_640 ();
 sg13g2_decap_8 FILLER_64_656 ();
 sg13g2_decap_8 FILLER_64_663 ();
 sg13g2_decap_8 FILLER_64_670 ();
 sg13g2_decap_4 FILLER_64_677 ();
 sg13g2_fill_2 FILLER_64_695 ();
 sg13g2_fill_1 FILLER_64_697 ();
 sg13g2_fill_2 FILLER_64_707 ();
 sg13g2_fill_2 FILLER_64_714 ();
 sg13g2_decap_8 FILLER_64_734 ();
 sg13g2_decap_4 FILLER_64_741 ();
 sg13g2_fill_2 FILLER_64_745 ();
 sg13g2_decap_8 FILLER_64_756 ();
 sg13g2_decap_4 FILLER_64_763 ();
 sg13g2_fill_2 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_809 ();
 sg13g2_fill_2 FILLER_64_816 ();
 sg13g2_decap_8 FILLER_64_822 ();
 sg13g2_decap_8 FILLER_64_829 ();
 sg13g2_decap_8 FILLER_64_836 ();
 sg13g2_decap_8 FILLER_64_843 ();
 sg13g2_decap_8 FILLER_64_850 ();
 sg13g2_decap_4 FILLER_64_857 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_fill_2 FILLER_65_238 ();
 sg13g2_fill_1 FILLER_65_240 ();
 sg13g2_decap_4 FILLER_65_267 ();
 sg13g2_fill_1 FILLER_65_271 ();
 sg13g2_decap_4 FILLER_65_305 ();
 sg13g2_fill_1 FILLER_65_309 ();
 sg13g2_decap_4 FILLER_65_315 ();
 sg13g2_fill_2 FILLER_65_319 ();
 sg13g2_fill_2 FILLER_65_328 ();
 sg13g2_fill_2 FILLER_65_333 ();
 sg13g2_fill_1 FILLER_65_335 ();
 sg13g2_decap_8 FILLER_65_345 ();
 sg13g2_decap_4 FILLER_65_386 ();
 sg13g2_fill_1 FILLER_65_390 ();
 sg13g2_fill_2 FILLER_65_409 ();
 sg13g2_fill_1 FILLER_65_419 ();
 sg13g2_decap_8 FILLER_65_476 ();
 sg13g2_decap_8 FILLER_65_483 ();
 sg13g2_decap_4 FILLER_65_490 ();
 sg13g2_fill_1 FILLER_65_494 ();
 sg13g2_fill_2 FILLER_65_499 ();
 sg13g2_fill_1 FILLER_65_501 ();
 sg13g2_decap_8 FILLER_65_510 ();
 sg13g2_fill_2 FILLER_65_517 ();
 sg13g2_fill_1 FILLER_65_529 ();
 sg13g2_decap_4 FILLER_65_572 ();
 sg13g2_fill_2 FILLER_65_576 ();
 sg13g2_decap_8 FILLER_65_586 ();
 sg13g2_fill_2 FILLER_65_593 ();
 sg13g2_fill_1 FILLER_65_595 ();
 sg13g2_fill_2 FILLER_65_622 ();
 sg13g2_fill_2 FILLER_65_678 ();
 sg13g2_decap_8 FILLER_65_711 ();
 sg13g2_decap_4 FILLER_65_718 ();
 sg13g2_fill_1 FILLER_65_722 ();
 sg13g2_decap_8 FILLER_65_728 ();
 sg13g2_fill_2 FILLER_65_735 ();
 sg13g2_decap_8 FILLER_65_764 ();
 sg13g2_fill_2 FILLER_65_771 ();
 sg13g2_fill_2 FILLER_65_783 ();
 sg13g2_fill_1 FILLER_65_785 ();
 sg13g2_decap_8 FILLER_65_789 ();
 sg13g2_decap_4 FILLER_65_796 ();
 sg13g2_fill_1 FILLER_65_800 ();
 sg13g2_fill_1 FILLER_65_806 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_65_847 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_4 FILLER_66_245 ();
 sg13g2_fill_2 FILLER_66_295 ();
 sg13g2_fill_1 FILLER_66_302 ();
 sg13g2_fill_2 FILLER_66_309 ();
 sg13g2_fill_1 FILLER_66_311 ();
 sg13g2_fill_2 FILLER_66_325 ();
 sg13g2_fill_1 FILLER_66_327 ();
 sg13g2_fill_2 FILLER_66_337 ();
 sg13g2_fill_1 FILLER_66_339 ();
 sg13g2_fill_2 FILLER_66_348 ();
 sg13g2_fill_1 FILLER_66_356 ();
 sg13g2_decap_8 FILLER_66_361 ();
 sg13g2_decap_8 FILLER_66_368 ();
 sg13g2_fill_2 FILLER_66_375 ();
 sg13g2_decap_4 FILLER_66_382 ();
 sg13g2_fill_2 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_423 ();
 sg13g2_fill_2 FILLER_66_430 ();
 sg13g2_fill_1 FILLER_66_432 ();
 sg13g2_fill_1 FILLER_66_447 ();
 sg13g2_decap_4 FILLER_66_521 ();
 sg13g2_fill_2 FILLER_66_534 ();
 sg13g2_fill_1 FILLER_66_536 ();
 sg13g2_decap_8 FILLER_66_545 ();
 sg13g2_decap_8 FILLER_66_552 ();
 sg13g2_decap_8 FILLER_66_559 ();
 sg13g2_decap_8 FILLER_66_566 ();
 sg13g2_decap_4 FILLER_66_573 ();
 sg13g2_fill_1 FILLER_66_577 ();
 sg13g2_decap_4 FILLER_66_590 ();
 sg13g2_fill_1 FILLER_66_594 ();
 sg13g2_decap_4 FILLER_66_600 ();
 sg13g2_decap_8 FILLER_66_617 ();
 sg13g2_fill_2 FILLER_66_624 ();
 sg13g2_fill_1 FILLER_66_626 ();
 sg13g2_fill_2 FILLER_66_645 ();
 sg13g2_decap_4 FILLER_66_675 ();
 sg13g2_decap_8 FILLER_66_685 ();
 sg13g2_decap_8 FILLER_66_692 ();
 sg13g2_fill_2 FILLER_66_699 ();
 sg13g2_decap_4 FILLER_66_711 ();
 sg13g2_decap_4 FILLER_66_741 ();
 sg13g2_fill_2 FILLER_66_745 ();
 sg13g2_decap_8 FILLER_66_754 ();
 sg13g2_decap_8 FILLER_66_761 ();
 sg13g2_fill_1 FILLER_66_768 ();
 sg13g2_decap_8 FILLER_66_787 ();
 sg13g2_fill_1 FILLER_66_794 ();
 sg13g2_decap_8 FILLER_66_799 ();
 sg13g2_decap_8 FILLER_66_806 ();
 sg13g2_decap_8 FILLER_66_813 ();
 sg13g2_decap_8 FILLER_66_820 ();
 sg13g2_decap_8 FILLER_66_827 ();
 sg13g2_decap_8 FILLER_66_834 ();
 sg13g2_decap_8 FILLER_66_841 ();
 sg13g2_decap_8 FILLER_66_848 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_fill_2 FILLER_67_245 ();
 sg13g2_fill_1 FILLER_67_247 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_266 ();
 sg13g2_decap_4 FILLER_67_281 ();
 sg13g2_fill_2 FILLER_67_299 ();
 sg13g2_decap_8 FILLER_67_320 ();
 sg13g2_decap_8 FILLER_67_327 ();
 sg13g2_decap_8 FILLER_67_334 ();
 sg13g2_decap_4 FILLER_67_341 ();
 sg13g2_fill_2 FILLER_67_345 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_403 ();
 sg13g2_fill_2 FILLER_67_410 ();
 sg13g2_fill_1 FILLER_67_412 ();
 sg13g2_decap_8 FILLER_67_444 ();
 sg13g2_decap_8 FILLER_67_451 ();
 sg13g2_decap_8 FILLER_67_458 ();
 sg13g2_decap_8 FILLER_67_465 ();
 sg13g2_decap_4 FILLER_67_472 ();
 sg13g2_fill_1 FILLER_67_476 ();
 sg13g2_decap_8 FILLER_67_481 ();
 sg13g2_decap_4 FILLER_67_488 ();
 sg13g2_fill_1 FILLER_67_492 ();
 sg13g2_decap_8 FILLER_67_497 ();
 sg13g2_fill_1 FILLER_67_504 ();
 sg13g2_fill_2 FILLER_67_510 ();
 sg13g2_fill_1 FILLER_67_512 ();
 sg13g2_decap_8 FILLER_67_518 ();
 sg13g2_decap_8 FILLER_67_525 ();
 sg13g2_decap_8 FILLER_67_547 ();
 sg13g2_fill_1 FILLER_67_554 ();
 sg13g2_decap_8 FILLER_67_592 ();
 sg13g2_fill_2 FILLER_67_599 ();
 sg13g2_fill_1 FILLER_67_601 ();
 sg13g2_decap_8 FILLER_67_607 ();
 sg13g2_fill_1 FILLER_67_614 ();
 sg13g2_decap_8 FILLER_67_628 ();
 sg13g2_decap_4 FILLER_67_635 ();
 sg13g2_fill_2 FILLER_67_639 ();
 sg13g2_decap_8 FILLER_67_673 ();
 sg13g2_fill_2 FILLER_67_680 ();
 sg13g2_fill_1 FILLER_67_682 ();
 sg13g2_decap_8 FILLER_67_696 ();
 sg13g2_fill_1 FILLER_67_703 ();
 sg13g2_decap_4 FILLER_67_746 ();
 sg13g2_fill_2 FILLER_67_750 ();
 sg13g2_decap_8 FILLER_67_775 ();
 sg13g2_fill_2 FILLER_67_782 ();
 sg13g2_decap_8 FILLER_67_810 ();
 sg13g2_decap_8 FILLER_67_817 ();
 sg13g2_decap_8 FILLER_67_824 ();
 sg13g2_decap_8 FILLER_67_831 ();
 sg13g2_decap_8 FILLER_67_838 ();
 sg13g2_decap_8 FILLER_67_845 ();
 sg13g2_decap_8 FILLER_67_852 ();
 sg13g2_fill_2 FILLER_67_859 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_4 FILLER_68_231 ();
 sg13g2_fill_1 FILLER_68_235 ();
 sg13g2_fill_2 FILLER_68_307 ();
 sg13g2_fill_1 FILLER_68_309 ();
 sg13g2_decap_8 FILLER_68_334 ();
 sg13g2_decap_4 FILLER_68_341 ();
 sg13g2_decap_8 FILLER_68_359 ();
 sg13g2_decap_4 FILLER_68_366 ();
 sg13g2_fill_2 FILLER_68_370 ();
 sg13g2_decap_8 FILLER_68_388 ();
 sg13g2_decap_8 FILLER_68_395 ();
 sg13g2_fill_1 FILLER_68_402 ();
 sg13g2_decap_8 FILLER_68_412 ();
 sg13g2_decap_4 FILLER_68_419 ();
 sg13g2_fill_1 FILLER_68_423 ();
 sg13g2_decap_8 FILLER_68_428 ();
 sg13g2_decap_8 FILLER_68_435 ();
 sg13g2_decap_8 FILLER_68_442 ();
 sg13g2_fill_2 FILLER_68_449 ();
 sg13g2_decap_8 FILLER_68_459 ();
 sg13g2_fill_1 FILLER_68_466 ();
 sg13g2_decap_8 FILLER_68_490 ();
 sg13g2_decap_4 FILLER_68_497 ();
 sg13g2_decap_8 FILLER_68_545 ();
 sg13g2_decap_4 FILLER_68_552 ();
 sg13g2_fill_2 FILLER_68_556 ();
 sg13g2_decap_8 FILLER_68_576 ();
 sg13g2_decap_8 FILLER_68_583 ();
 sg13g2_decap_4 FILLER_68_590 ();
 sg13g2_fill_2 FILLER_68_594 ();
 sg13g2_decap_8 FILLER_68_632 ();
 sg13g2_decap_4 FILLER_68_639 ();
 sg13g2_decap_4 FILLER_68_669 ();
 sg13g2_decap_8 FILLER_68_743 ();
 sg13g2_fill_2 FILLER_68_750 ();
 sg13g2_fill_1 FILLER_68_752 ();
 sg13g2_decap_8 FILLER_68_788 ();
 sg13g2_decap_8 FILLER_68_795 ();
 sg13g2_decap_8 FILLER_68_802 ();
 sg13g2_decap_8 FILLER_68_809 ();
 sg13g2_decap_8 FILLER_68_816 ();
 sg13g2_decap_8 FILLER_68_823 ();
 sg13g2_decap_8 FILLER_68_830 ();
 sg13g2_decap_8 FILLER_68_837 ();
 sg13g2_decap_8 FILLER_68_844 ();
 sg13g2_decap_8 FILLER_68_851 ();
 sg13g2_decap_4 FILLER_68_858 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_189 ();
 sg13g2_decap_8 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_4 FILLER_69_252 ();
 sg13g2_fill_2 FILLER_69_256 ();
 sg13g2_fill_1 FILLER_69_267 ();
 sg13g2_decap_8 FILLER_69_281 ();
 sg13g2_decap_8 FILLER_69_293 ();
 sg13g2_decap_8 FILLER_69_300 ();
 sg13g2_fill_2 FILLER_69_324 ();
 sg13g2_decap_8 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_4 FILLER_69_343 ();
 sg13g2_fill_1 FILLER_69_347 ();
 sg13g2_decap_4 FILLER_69_367 ();
 sg13g2_fill_2 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_fill_2 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_417 ();
 sg13g2_fill_1 FILLER_69_424 ();
 sg13g2_decap_8 FILLER_69_428 ();
 sg13g2_fill_2 FILLER_69_461 ();
 sg13g2_fill_1 FILLER_69_463 ();
 sg13g2_decap_8 FILLER_69_495 ();
 sg13g2_fill_2 FILLER_69_510 ();
 sg13g2_decap_8 FILLER_69_516 ();
 sg13g2_decap_4 FILLER_69_523 ();
 sg13g2_fill_1 FILLER_69_527 ();
 sg13g2_fill_2 FILLER_69_549 ();
 sg13g2_decap_4 FILLER_69_568 ();
 sg13g2_fill_1 FILLER_69_581 ();
 sg13g2_decap_4 FILLER_69_588 ();
 sg13g2_fill_2 FILLER_69_592 ();
 sg13g2_fill_1 FILLER_69_599 ();
 sg13g2_decap_8 FILLER_69_612 ();
 sg13g2_decap_4 FILLER_69_619 ();
 sg13g2_fill_2 FILLER_69_623 ();
 sg13g2_decap_4 FILLER_69_634 ();
 sg13g2_fill_2 FILLER_69_657 ();
 sg13g2_fill_1 FILLER_69_659 ();
 sg13g2_decap_8 FILLER_69_676 ();
 sg13g2_fill_2 FILLER_69_683 ();
 sg13g2_fill_2 FILLER_69_694 ();
 sg13g2_fill_1 FILLER_69_696 ();
 sg13g2_fill_2 FILLER_69_720 ();
 sg13g2_decap_8 FILLER_69_748 ();
 sg13g2_decap_8 FILLER_69_755 ();
 sg13g2_decap_8 FILLER_69_762 ();
 sg13g2_decap_8 FILLER_69_769 ();
 sg13g2_decap_8 FILLER_69_776 ();
 sg13g2_decap_8 FILLER_69_783 ();
 sg13g2_decap_8 FILLER_69_790 ();
 sg13g2_decap_8 FILLER_69_797 ();
 sg13g2_decap_8 FILLER_69_804 ();
 sg13g2_decap_8 FILLER_69_811 ();
 sg13g2_decap_8 FILLER_69_818 ();
 sg13g2_decap_8 FILLER_69_825 ();
 sg13g2_decap_8 FILLER_69_832 ();
 sg13g2_decap_8 FILLER_69_839 ();
 sg13g2_decap_8 FILLER_69_846 ();
 sg13g2_decap_8 FILLER_69_853 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_fill_1 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_303 ();
 sg13g2_fill_1 FILLER_70_305 ();
 sg13g2_fill_2 FILLER_70_342 ();
 sg13g2_fill_1 FILLER_70_344 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_fill_1 FILLER_70_357 ();
 sg13g2_decap_4 FILLER_70_374 ();
 sg13g2_fill_2 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_4 FILLER_70_399 ();
 sg13g2_decap_4 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_70_412 ();
 sg13g2_fill_1 FILLER_70_420 ();
 sg13g2_decap_4 FILLER_70_437 ();
 sg13g2_fill_2 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_456 ();
 sg13g2_decap_4 FILLER_70_463 ();
 sg13g2_decap_8 FILLER_70_479 ();
 sg13g2_fill_2 FILLER_70_486 ();
 sg13g2_fill_1 FILLER_70_488 ();
 sg13g2_decap_8 FILLER_70_493 ();
 sg13g2_fill_1 FILLER_70_500 ();
 sg13g2_decap_8 FILLER_70_513 ();
 sg13g2_decap_4 FILLER_70_520 ();
 sg13g2_fill_2 FILLER_70_524 ();
 sg13g2_decap_8 FILLER_70_530 ();
 sg13g2_fill_2 FILLER_70_537 ();
 sg13g2_fill_2 FILLER_70_544 ();
 sg13g2_decap_8 FILLER_70_554 ();
 sg13g2_decap_8 FILLER_70_561 ();
 sg13g2_decap_8 FILLER_70_568 ();
 sg13g2_fill_2 FILLER_70_575 ();
 sg13g2_fill_1 FILLER_70_577 ();
 sg13g2_fill_2 FILLER_70_598 ();
 sg13g2_decap_4 FILLER_70_610 ();
 sg13g2_fill_1 FILLER_70_614 ();
 sg13g2_decap_8 FILLER_70_641 ();
 sg13g2_decap_8 FILLER_70_648 ();
 sg13g2_decap_8 FILLER_70_694 ();
 sg13g2_fill_1 FILLER_70_701 ();
 sg13g2_decap_8 FILLER_70_728 ();
 sg13g2_decap_8 FILLER_70_735 ();
 sg13g2_decap_8 FILLER_70_742 ();
 sg13g2_decap_8 FILLER_70_749 ();
 sg13g2_decap_8 FILLER_70_756 ();
 sg13g2_decap_8 FILLER_70_763 ();
 sg13g2_decap_8 FILLER_70_770 ();
 sg13g2_decap_8 FILLER_70_777 ();
 sg13g2_decap_8 FILLER_70_784 ();
 sg13g2_decap_8 FILLER_70_791 ();
 sg13g2_decap_8 FILLER_70_798 ();
 sg13g2_decap_8 FILLER_70_805 ();
 sg13g2_decap_8 FILLER_70_812 ();
 sg13g2_decap_8 FILLER_70_819 ();
 sg13g2_decap_8 FILLER_70_826 ();
 sg13g2_decap_8 FILLER_70_833 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_4 FILLER_71_252 ();
 sg13g2_fill_1 FILLER_71_256 ();
 sg13g2_decap_8 FILLER_71_261 ();
 sg13g2_decap_8 FILLER_71_268 ();
 sg13g2_decap_8 FILLER_71_275 ();
 sg13g2_decap_4 FILLER_71_282 ();
 sg13g2_fill_1 FILLER_71_286 ();
 sg13g2_decap_8 FILLER_71_291 ();
 sg13g2_decap_8 FILLER_71_298 ();
 sg13g2_fill_1 FILLER_71_305 ();
 sg13g2_decap_8 FILLER_71_323 ();
 sg13g2_decap_8 FILLER_71_330 ();
 sg13g2_decap_4 FILLER_71_337 ();
 sg13g2_decap_4 FILLER_71_345 ();
 sg13g2_fill_2 FILLER_71_349 ();
 sg13g2_fill_2 FILLER_71_356 ();
 sg13g2_decap_4 FILLER_71_367 ();
 sg13g2_fill_1 FILLER_71_376 ();
 sg13g2_fill_2 FILLER_71_402 ();
 sg13g2_fill_2 FILLER_71_410 ();
 sg13g2_fill_2 FILLER_71_426 ();
 sg13g2_decap_8 FILLER_71_433 ();
 sg13g2_decap_8 FILLER_71_440 ();
 sg13g2_fill_1 FILLER_71_447 ();
 sg13g2_decap_8 FILLER_71_452 ();
 sg13g2_decap_8 FILLER_71_459 ();
 sg13g2_fill_2 FILLER_71_466 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_decap_4 FILLER_71_541 ();
 sg13g2_decap_4 FILLER_71_576 ();
 sg13g2_fill_1 FILLER_71_580 ();
 sg13g2_decap_8 FILLER_71_587 ();
 sg13g2_decap_8 FILLER_71_594 ();
 sg13g2_decap_8 FILLER_71_611 ();
 sg13g2_decap_8 FILLER_71_618 ();
 sg13g2_fill_2 FILLER_71_629 ();
 sg13g2_fill_1 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_663 ();
 sg13g2_fill_2 FILLER_71_678 ();
 sg13g2_decap_8 FILLER_71_693 ();
 sg13g2_decap_4 FILLER_71_700 ();
 sg13g2_decap_8 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_733 ();
 sg13g2_decap_8 FILLER_71_740 ();
 sg13g2_decap_8 FILLER_71_747 ();
 sg13g2_decap_8 FILLER_71_754 ();
 sg13g2_decap_8 FILLER_71_761 ();
 sg13g2_decap_8 FILLER_71_768 ();
 sg13g2_decap_8 FILLER_71_775 ();
 sg13g2_decap_8 FILLER_71_782 ();
 sg13g2_decap_8 FILLER_71_789 ();
 sg13g2_decap_8 FILLER_71_796 ();
 sg13g2_decap_8 FILLER_71_803 ();
 sg13g2_decap_8 FILLER_71_810 ();
 sg13g2_decap_8 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_824 ();
 sg13g2_decap_8 FILLER_71_831 ();
 sg13g2_decap_8 FILLER_71_838 ();
 sg13g2_decap_8 FILLER_71_845 ();
 sg13g2_decap_8 FILLER_71_852 ();
 sg13g2_fill_2 FILLER_71_859 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_decap_4 FILLER_72_326 ();
 sg13g2_decap_8 FILLER_72_356 ();
 sg13g2_decap_8 FILLER_72_376 ();
 sg13g2_decap_8 FILLER_72_383 ();
 sg13g2_fill_1 FILLER_72_390 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_fill_1 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_423 ();
 sg13g2_decap_8 FILLER_72_430 ();
 sg13g2_fill_1 FILLER_72_437 ();
 sg13g2_decap_8 FILLER_72_464 ();
 sg13g2_fill_2 FILLER_72_471 ();
 sg13g2_fill_1 FILLER_72_473 ();
 sg13g2_fill_2 FILLER_72_486 ();
 sg13g2_fill_1 FILLER_72_488 ();
 sg13g2_decap_8 FILLER_72_498 ();
 sg13g2_decap_8 FILLER_72_505 ();
 sg13g2_decap_8 FILLER_72_512 ();
 sg13g2_decap_8 FILLER_72_519 ();
 sg13g2_decap_8 FILLER_72_526 ();
 sg13g2_decap_8 FILLER_72_533 ();
 sg13g2_decap_4 FILLER_72_540 ();
 sg13g2_fill_1 FILLER_72_544 ();
 sg13g2_decap_4 FILLER_72_550 ();
 sg13g2_decap_8 FILLER_72_589 ();
 sg13g2_decap_4 FILLER_72_596 ();
 sg13g2_decap_4 FILLER_72_605 ();
 sg13g2_fill_2 FILLER_72_609 ();
 sg13g2_decap_8 FILLER_72_703 ();
 sg13g2_decap_8 FILLER_72_710 ();
 sg13g2_decap_8 FILLER_72_717 ();
 sg13g2_decap_8 FILLER_72_724 ();
 sg13g2_decap_8 FILLER_72_731 ();
 sg13g2_decap_8 FILLER_72_738 ();
 sg13g2_decap_8 FILLER_72_745 ();
 sg13g2_decap_8 FILLER_72_752 ();
 sg13g2_decap_8 FILLER_72_759 ();
 sg13g2_decap_8 FILLER_72_766 ();
 sg13g2_decap_8 FILLER_72_773 ();
 sg13g2_decap_8 FILLER_72_780 ();
 sg13g2_decap_8 FILLER_72_787 ();
 sg13g2_decap_8 FILLER_72_794 ();
 sg13g2_decap_8 FILLER_72_801 ();
 sg13g2_decap_8 FILLER_72_808 ();
 sg13g2_decap_8 FILLER_72_815 ();
 sg13g2_decap_8 FILLER_72_822 ();
 sg13g2_decap_8 FILLER_72_829 ();
 sg13g2_decap_8 FILLER_72_836 ();
 sg13g2_decap_8 FILLER_72_843 ();
 sg13g2_decap_8 FILLER_72_850 ();
 sg13g2_decap_4 FILLER_72_857 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_305 ();
 sg13g2_decap_8 FILLER_73_312 ();
 sg13g2_decap_4 FILLER_73_319 ();
 sg13g2_fill_2 FILLER_73_323 ();
 sg13g2_decap_4 FILLER_73_334 ();
 sg13g2_fill_1 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_356 ();
 sg13g2_fill_2 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_370 ();
 sg13g2_fill_2 FILLER_73_377 ();
 sg13g2_decap_8 FILLER_73_384 ();
 sg13g2_decap_4 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_441 ();
 sg13g2_fill_1 FILLER_73_452 ();
 sg13g2_decap_4 FILLER_73_458 ();
 sg13g2_decap_8 FILLER_73_466 ();
 sg13g2_decap_8 FILLER_73_473 ();
 sg13g2_decap_4 FILLER_73_480 ();
 sg13g2_decap_4 FILLER_73_536 ();
 sg13g2_decap_8 FILLER_73_556 ();
 sg13g2_fill_2 FILLER_73_572 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_4 FILLER_73_585 ();
 sg13g2_fill_1 FILLER_73_589 ();
 sg13g2_decap_8 FILLER_73_611 ();
 sg13g2_decap_4 FILLER_73_618 ();
 sg13g2_decap_8 FILLER_73_626 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_decap_8 FILLER_73_640 ();
 sg13g2_fill_1 FILLER_73_654 ();
 sg13g2_decap_4 FILLER_73_681 ();
 sg13g2_fill_1 FILLER_73_685 ();
 sg13g2_decap_8 FILLER_73_699 ();
 sg13g2_decap_8 FILLER_73_706 ();
 sg13g2_decap_8 FILLER_73_713 ();
 sg13g2_decap_8 FILLER_73_720 ();
 sg13g2_decap_8 FILLER_73_727 ();
 sg13g2_decap_8 FILLER_73_734 ();
 sg13g2_decap_8 FILLER_73_741 ();
 sg13g2_decap_8 FILLER_73_748 ();
 sg13g2_decap_8 FILLER_73_755 ();
 sg13g2_decap_8 FILLER_73_762 ();
 sg13g2_decap_8 FILLER_73_769 ();
 sg13g2_decap_8 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_decap_8 FILLER_73_790 ();
 sg13g2_decap_8 FILLER_73_797 ();
 sg13g2_decap_8 FILLER_73_804 ();
 sg13g2_decap_8 FILLER_73_811 ();
 sg13g2_decap_8 FILLER_73_818 ();
 sg13g2_decap_8 FILLER_73_825 ();
 sg13g2_decap_8 FILLER_73_832 ();
 sg13g2_decap_8 FILLER_73_839 ();
 sg13g2_decap_8 FILLER_73_846 ();
 sg13g2_decap_8 FILLER_73_853 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_fill_2 FILLER_74_308 ();
 sg13g2_fill_1 FILLER_74_310 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_fill_1 FILLER_74_354 ();
 sg13g2_fill_2 FILLER_74_381 ();
 sg13g2_fill_1 FILLER_74_383 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_fill_2 FILLER_74_403 ();
 sg13g2_fill_1 FILLER_74_405 ();
 sg13g2_decap_8 FILLER_74_410 ();
 sg13g2_fill_1 FILLER_74_417 ();
 sg13g2_fill_2 FILLER_74_449 ();
 sg13g2_decap_4 FILLER_74_477 ();
 sg13g2_fill_2 FILLER_74_481 ();
 sg13g2_decap_8 FILLER_74_501 ();
 sg13g2_fill_2 FILLER_74_508 ();
 sg13g2_fill_2 FILLER_74_514 ();
 sg13g2_fill_1 FILLER_74_516 ();
 sg13g2_decap_8 FILLER_74_529 ();
 sg13g2_decap_8 FILLER_74_536 ();
 sg13g2_decap_8 FILLER_74_547 ();
 sg13g2_fill_2 FILLER_74_554 ();
 sg13g2_fill_1 FILLER_74_556 ();
 sg13g2_decap_8 FILLER_74_610 ();
 sg13g2_fill_2 FILLER_74_617 ();
 sg13g2_decap_8 FILLER_74_624 ();
 sg13g2_decap_4 FILLER_74_631 ();
 sg13g2_fill_1 FILLER_74_635 ();
 sg13g2_decap_4 FILLER_74_653 ();
 sg13g2_decap_8 FILLER_74_670 ();
 sg13g2_decap_8 FILLER_74_677 ();
 sg13g2_decap_8 FILLER_74_684 ();
 sg13g2_decap_8 FILLER_74_691 ();
 sg13g2_decap_8 FILLER_74_698 ();
 sg13g2_decap_8 FILLER_74_705 ();
 sg13g2_decap_8 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_719 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_740 ();
 sg13g2_decap_8 FILLER_74_747 ();
 sg13g2_decap_8 FILLER_74_754 ();
 sg13g2_decap_8 FILLER_74_761 ();
 sg13g2_decap_8 FILLER_74_768 ();
 sg13g2_decap_8 FILLER_74_775 ();
 sg13g2_decap_8 FILLER_74_782 ();
 sg13g2_decap_8 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_796 ();
 sg13g2_decap_8 FILLER_74_803 ();
 sg13g2_decap_8 FILLER_74_810 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_8 FILLER_74_824 ();
 sg13g2_decap_8 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_4 FILLER_75_315 ();
 sg13g2_fill_2 FILLER_75_319 ();
 sg13g2_decap_8 FILLER_75_325 ();
 sg13g2_decap_8 FILLER_75_332 ();
 sg13g2_decap_8 FILLER_75_339 ();
 sg13g2_decap_8 FILLER_75_346 ();
 sg13g2_decap_8 FILLER_75_353 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_fill_2 FILLER_75_374 ();
 sg13g2_fill_1 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_decap_4 FILLER_75_402 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_416 ();
 sg13g2_decap_8 FILLER_75_423 ();
 sg13g2_decap_8 FILLER_75_430 ();
 sg13g2_decap_8 FILLER_75_437 ();
 sg13g2_fill_1 FILLER_75_453 ();
 sg13g2_fill_2 FILLER_75_468 ();
 sg13g2_decap_8 FILLER_75_495 ();
 sg13g2_fill_1 FILLER_75_502 ();
 sg13g2_fill_2 FILLER_75_513 ();
 sg13g2_decap_8 FILLER_75_531 ();
 sg13g2_decap_8 FILLER_75_538 ();
 sg13g2_decap_8 FILLER_75_568 ();
 sg13g2_decap_8 FILLER_75_575 ();
 sg13g2_decap_4 FILLER_75_582 ();
 sg13g2_fill_1 FILLER_75_586 ();
 sg13g2_decap_4 FILLER_75_605 ();
 sg13g2_fill_2 FILLER_75_609 ();
 sg13g2_fill_2 FILLER_75_645 ();
 sg13g2_fill_1 FILLER_75_647 ();
 sg13g2_decap_8 FILLER_75_674 ();
 sg13g2_decap_8 FILLER_75_681 ();
 sg13g2_decap_8 FILLER_75_688 ();
 sg13g2_decap_8 FILLER_75_695 ();
 sg13g2_decap_8 FILLER_75_702 ();
 sg13g2_decap_8 FILLER_75_709 ();
 sg13g2_decap_8 FILLER_75_716 ();
 sg13g2_decap_8 FILLER_75_723 ();
 sg13g2_decap_8 FILLER_75_730 ();
 sg13g2_decap_8 FILLER_75_737 ();
 sg13g2_decap_8 FILLER_75_744 ();
 sg13g2_decap_8 FILLER_75_751 ();
 sg13g2_decap_8 FILLER_75_758 ();
 sg13g2_decap_8 FILLER_75_765 ();
 sg13g2_decap_8 FILLER_75_772 ();
 sg13g2_decap_8 FILLER_75_779 ();
 sg13g2_decap_8 FILLER_75_786 ();
 sg13g2_decap_8 FILLER_75_793 ();
 sg13g2_decap_8 FILLER_75_800 ();
 sg13g2_decap_8 FILLER_75_807 ();
 sg13g2_decap_8 FILLER_75_814 ();
 sg13g2_decap_8 FILLER_75_821 ();
 sg13g2_decap_8 FILLER_75_828 ();
 sg13g2_decap_8 FILLER_75_835 ();
 sg13g2_decap_8 FILLER_75_842 ();
 sg13g2_decap_8 FILLER_75_849 ();
 sg13g2_decap_4 FILLER_75_856 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_fill_2 FILLER_76_385 ();
 sg13g2_decap_4 FILLER_76_413 ();
 sg13g2_fill_1 FILLER_76_417 ();
 sg13g2_fill_2 FILLER_76_484 ();
 sg13g2_decap_8 FILLER_76_505 ();
 sg13g2_decap_8 FILLER_76_512 ();
 sg13g2_decap_8 FILLER_76_519 ();
 sg13g2_decap_8 FILLER_76_526 ();
 sg13g2_decap_8 FILLER_76_533 ();
 sg13g2_fill_1 FILLER_76_540 ();
 sg13g2_fill_2 FILLER_76_554 ();
 sg13g2_fill_1 FILLER_76_556 ();
 sg13g2_decap_8 FILLER_76_573 ();
 sg13g2_decap_8 FILLER_76_580 ();
 sg13g2_fill_2 FILLER_76_587 ();
 sg13g2_fill_1 FILLER_76_589 ();
 sg13g2_fill_1 FILLER_76_600 ();
 sg13g2_decap_4 FILLER_76_611 ();
 sg13g2_fill_1 FILLER_76_615 ();
 sg13g2_fill_2 FILLER_76_625 ();
 sg13g2_decap_8 FILLER_76_640 ();
 sg13g2_fill_1 FILLER_76_647 ();
 sg13g2_decap_8 FILLER_76_657 ();
 sg13g2_decap_8 FILLER_76_664 ();
 sg13g2_decap_8 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_678 ();
 sg13g2_decap_8 FILLER_76_685 ();
 sg13g2_decap_8 FILLER_76_692 ();
 sg13g2_decap_8 FILLER_76_699 ();
 sg13g2_decap_8 FILLER_76_706 ();
 sg13g2_decap_8 FILLER_76_713 ();
 sg13g2_decap_8 FILLER_76_720 ();
 sg13g2_decap_8 FILLER_76_727 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_decap_8 FILLER_76_741 ();
 sg13g2_decap_8 FILLER_76_748 ();
 sg13g2_decap_8 FILLER_76_755 ();
 sg13g2_decap_8 FILLER_76_762 ();
 sg13g2_decap_8 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_776 ();
 sg13g2_decap_8 FILLER_76_783 ();
 sg13g2_decap_8 FILLER_76_790 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_804 ();
 sg13g2_decap_8 FILLER_76_811 ();
 sg13g2_decap_8 FILLER_76_818 ();
 sg13g2_decap_8 FILLER_76_825 ();
 sg13g2_decap_8 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_839 ();
 sg13g2_decap_8 FILLER_76_846 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_fill_1 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_437 ();
 sg13g2_fill_1 FILLER_77_472 ();
 sg13g2_fill_2 FILLER_77_482 ();
 sg13g2_fill_2 FILLER_77_493 ();
 sg13g2_decap_8 FILLER_77_503 ();
 sg13g2_fill_2 FILLER_77_510 ();
 sg13g2_fill_2 FILLER_77_524 ();
 sg13g2_decap_8 FILLER_77_534 ();
 sg13g2_decap_8 FILLER_77_541 ();
 sg13g2_decap_8 FILLER_77_548 ();
 sg13g2_fill_2 FILLER_77_555 ();
 sg13g2_decap_4 FILLER_77_565 ();
 sg13g2_fill_2 FILLER_77_569 ();
 sg13g2_fill_1 FILLER_77_595 ();
 sg13g2_fill_2 FILLER_77_637 ();
 sg13g2_fill_1 FILLER_77_639 ();
 sg13g2_decap_8 FILLER_77_671 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_decap_8 FILLER_77_685 ();
 sg13g2_decap_8 FILLER_77_692 ();
 sg13g2_decap_8 FILLER_77_699 ();
 sg13g2_decap_8 FILLER_77_706 ();
 sg13g2_decap_8 FILLER_77_713 ();
 sg13g2_decap_8 FILLER_77_720 ();
 sg13g2_decap_8 FILLER_77_727 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_decap_8 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_776 ();
 sg13g2_decap_8 FILLER_77_783 ();
 sg13g2_decap_8 FILLER_77_790 ();
 sg13g2_decap_8 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_decap_8 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_832 ();
 sg13g2_decap_8 FILLER_77_839 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_fill_1 FILLER_78_448 ();
 sg13g2_fill_2 FILLER_78_475 ();
 sg13g2_decap_8 FILLER_78_515 ();
 sg13g2_decap_8 FILLER_78_522 ();
 sg13g2_fill_1 FILLER_78_529 ();
 sg13g2_decap_8 FILLER_78_554 ();
 sg13g2_decap_8 FILLER_78_561 ();
 sg13g2_decap_8 FILLER_78_568 ();
 sg13g2_decap_8 FILLER_78_575 ();
 sg13g2_decap_8 FILLER_78_582 ();
 sg13g2_decap_8 FILLER_78_589 ();
 sg13g2_decap_8 FILLER_78_596 ();
 sg13g2_decap_8 FILLER_78_603 ();
 sg13g2_decap_8 FILLER_78_632 ();
 sg13g2_decap_8 FILLER_78_639 ();
 sg13g2_decap_4 FILLER_78_646 ();
 sg13g2_decap_8 FILLER_78_654 ();
 sg13g2_decap_8 FILLER_78_661 ();
 sg13g2_decap_8 FILLER_78_668 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_fill_2 FILLER_78_682 ();
 sg13g2_fill_1 FILLER_78_684 ();
 sg13g2_decap_8 FILLER_78_690 ();
 sg13g2_decap_8 FILLER_78_697 ();
 sg13g2_decap_8 FILLER_78_704 ();
 sg13g2_decap_8 FILLER_78_711 ();
 sg13g2_decap_8 FILLER_78_718 ();
 sg13g2_decap_8 FILLER_78_725 ();
 sg13g2_decap_8 FILLER_78_732 ();
 sg13g2_decap_8 FILLER_78_739 ();
 sg13g2_decap_8 FILLER_78_746 ();
 sg13g2_decap_8 FILLER_78_753 ();
 sg13g2_decap_8 FILLER_78_760 ();
 sg13g2_decap_8 FILLER_78_767 ();
 sg13g2_decap_8 FILLER_78_774 ();
 sg13g2_decap_8 FILLER_78_781 ();
 sg13g2_decap_8 FILLER_78_788 ();
 sg13g2_decap_8 FILLER_78_795 ();
 sg13g2_decap_8 FILLER_78_802 ();
 sg13g2_decap_8 FILLER_78_809 ();
 sg13g2_decap_8 FILLER_78_816 ();
 sg13g2_decap_8 FILLER_78_823 ();
 sg13g2_decap_8 FILLER_78_830 ();
 sg13g2_decap_8 FILLER_78_837 ();
 sg13g2_decap_8 FILLER_78_844 ();
 sg13g2_decap_8 FILLER_78_851 ();
 sg13g2_decap_4 FILLER_78_858 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_4 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_461 ();
 sg13g2_decap_4 FILLER_79_468 ();
 sg13g2_decap_8 FILLER_79_475 ();
 sg13g2_fill_2 FILLER_79_482 ();
 sg13g2_fill_2 FILLER_79_510 ();
 sg13g2_fill_1 FILLER_79_512 ();
 sg13g2_fill_1 FILLER_79_539 ();
 sg13g2_fill_2 FILLER_79_544 ();
 sg13g2_decap_8 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_631 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_667 ();
 sg13g2_decap_8 FILLER_79_674 ();
 sg13g2_decap_8 FILLER_79_681 ();
 sg13g2_decap_8 FILLER_79_688 ();
 sg13g2_decap_8 FILLER_79_695 ();
 sg13g2_decap_8 FILLER_79_702 ();
 sg13g2_decap_8 FILLER_79_709 ();
 sg13g2_decap_8 FILLER_79_716 ();
 sg13g2_decap_8 FILLER_79_723 ();
 sg13g2_decap_8 FILLER_79_730 ();
 sg13g2_decap_8 FILLER_79_737 ();
 sg13g2_decap_8 FILLER_79_744 ();
 sg13g2_decap_8 FILLER_79_751 ();
 sg13g2_decap_8 FILLER_79_758 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_decap_8 FILLER_79_772 ();
 sg13g2_decap_8 FILLER_79_779 ();
 sg13g2_decap_8 FILLER_79_786 ();
 sg13g2_decap_8 FILLER_79_793 ();
 sg13g2_decap_8 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_807 ();
 sg13g2_decap_8 FILLER_79_814 ();
 sg13g2_decap_8 FILLER_79_821 ();
 sg13g2_decap_8 FILLER_79_828 ();
 sg13g2_decap_8 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_decap_8 FILLER_79_849 ();
 sg13g2_decap_4 FILLER_79_856 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_355 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_4 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_451 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_fill_2 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_499 ();
 sg13g2_decap_8 FILLER_80_506 ();
 sg13g2_decap_8 FILLER_80_513 ();
 sg13g2_decap_4 FILLER_80_520 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_decap_4 FILLER_80_574 ();
 sg13g2_decap_8 FILLER_80_582 ();
 sg13g2_decap_8 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_fill_1 FILLER_80_603 ();
 sg13g2_fill_2 FILLER_80_608 ();
 sg13g2_fill_1 FILLER_80_610 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_decap_8 FILLER_80_851 ();
 sg13g2_decap_4 FILLER_80_858 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule
