module tt_um_algofoogle_ro_worker (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire \ca[0] ;
 wire \ca[10] ;
 wire \ca[11] ;
 wire \ca[12] ;
 wire \ca[13] ;
 wire \ca[14] ;
 wire \ca[15] ;
 wire \ca[1] ;
 wire \ca[2] ;
 wire \ca[3] ;
 wire \ca[4] ;
 wire \ca[5] ;
 wire \ca[6] ;
 wire \ca[7] ;
 wire \ca[8] ;
 wire \ca[9] ;
 wire \cb[0] ;
 wire \cb[10] ;
 wire \cb[11] ;
 wire \cb[12] ;
 wire \cb[13] ;
 wire \cb[14] ;
 wire \cb[15] ;
 wire \cb[1] ;
 wire \cb[2] ;
 wire \cb[3] ;
 wire \cb[4] ;
 wire \cb[5] ;
 wire \cb[6] ;
 wire \cb[7] ;
 wire \cb[8] ;
 wire \cb[9] ;
 wire \clock_div[0] ;
 wire \clock_div[1] ;
 wire \clock_div[2] ;
 wire \clock_div[3] ;
 wire \da[0] ;
 wire \da[10] ;
 wire \da[11] ;
 wire \da[12] ;
 wire \da[13] ;
 wire \da[14] ;
 wire \da[15] ;
 wire \da[1] ;
 wire \da[2] ;
 wire \da[3] ;
 wire \da[4] ;
 wire \da[5] ;
 wire \da[6] ;
 wire \da[7] ;
 wire \da[8] ;
 wire \da[9] ;
 wire \db[0] ;
 wire \db[10] ;
 wire \db[11] ;
 wire \db[12] ;
 wire \db[13] ;
 wire \db[14] ;
 wire \db[15] ;
 wire \db[1] ;
 wire \db[2] ;
 wire \db[3] ;
 wire \db[4] ;
 wire \db[5] ;
 wire \db[6] ;
 wire \db[7] ;
 wire \db[8] ;
 wire \db[9] ;
 wire done;
 wire internal_clock;
 wire internal_clock_unbuffered;
 wire \myring.inv_in[0] ;
 wire \myring.inv_in[1] ;
 wire \myring.inv_in[2] ;
 wire \myring.inv_in[3] ;
 wire \myring.inv_in[4] ;
 wire \myring.inv_in[5] ;
 wire \myring.inv_in[6] ;
 wire \myring.inv_in[7] ;
 wire \myring.inv_in[8] ;
 wire \myring.inv_out[8] ;
 wire reset;
 wire \resetsync.buff[0] ;
 wire \resetsync.in ;
 wire run;
 wire \shift_counter[0] ;
 wire \shift_counter[1] ;
 wire \shiftedge.buff[0] ;
 wire \shiftedge.buff[1] ;
 wire \shiftedge.buff[2] ;
 wire \shiftedge.buff[3] ;
 wire \stopedge.buff[0] ;
 wire \stopedge.buff[1] ;
 wire \stopedge.buff[2] ;
 wire \stopedge.buff[3] ;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net172;
 wire net173;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;

 sg13g2_inv_1 _0615_ (.Y(_0084_),
    .A(_0002_));
 sg13g2_inv_1 _0616_ (.Y(_0085_),
    .A(\cb[15] ));
 sg13g2_inv_1 _0617_ (.Y(_0086_),
    .A(\cb[14] ));
 sg13g2_inv_1 _0618_ (.Y(_0087_),
    .A(\cb[13] ));
 sg13g2_inv_1 _0619_ (.Y(_0088_),
    .A(\cb[12] ));
 sg13g2_inv_1 _0620_ (.Y(_0089_),
    .A(\cb[10] ));
 sg13g2_inv_1 _0621_ (.Y(_0090_),
    .A(\cb[9] ));
 sg13g2_inv_1 _0622_ (.Y(_0091_),
    .A(\cb[7] ));
 sg13g2_inv_1 _0623_ (.Y(_0092_),
    .A(\cb[4] ));
 sg13g2_inv_1 _0624_ (.Y(_0093_),
    .A(\cb[2] ));
 sg13g2_inv_1 _0625_ (.Y(_0094_),
    .A(\cb[1] ));
 sg13g2_inv_1 _0626_ (.Y(_0095_),
    .A(\cb[0] ));
 sg13g2_inv_1 _0627_ (.Y(_0096_),
    .A(\ca[13] ));
 sg13g2_inv_1 _0628_ (.Y(_0097_),
    .A(\ca[12] ));
 sg13g2_inv_1 _0629_ (.Y(_0098_),
    .A(\ca[10] ));
 sg13g2_inv_1 _0630_ (.Y(_0099_),
    .A(\ca[8] ));
 sg13g2_inv_1 _0631_ (.Y(_0100_),
    .A(\ca[7] ));
 sg13g2_inv_1 _0632_ (.Y(_0101_),
    .A(\db[15] ));
 sg13g2_inv_2 _0633_ (.Y(_0102_),
    .A(\db[7] ));
 sg13g2_inv_1 _0634_ (.Y(_0103_),
    .A(\db[6] ));
 sg13g2_inv_1 _0635_ (.Y(_0104_),
    .A(\db[13] ));
 sg13g2_inv_1 _0636_ (.Y(_0105_),
    .A(\db[5] ));
 sg13g2_inv_1 _0637_ (.Y(_0106_),
    .A(\db[12] ));
 sg13g2_inv_1 _0638_ (.Y(_0107_),
    .A(\db[4] ));
 sg13g2_inv_1 _0639_ (.Y(_0108_),
    .A(\db[3] ));
 sg13g2_inv_1 _0640_ (.Y(_0109_),
    .A(\db[2] ));
 sg13g2_inv_1 _0641_ (.Y(_0110_),
    .A(\db[9] ));
 sg13g2_inv_1 _0642_ (.Y(_0111_),
    .A(\db[1] ));
 sg13g2_inv_1 _0643_ (.Y(_0112_),
    .A(\db[0] ));
 sg13g2_inv_1 _0644_ (.Y(_0113_),
    .A(\da[7] ));
 sg13g2_inv_1 _0645_ (.Y(_0114_),
    .A(\da[6] ));
 sg13g2_inv_1 _0646_ (.Y(_0115_),
    .A(\da[5] ));
 sg13g2_inv_1 _0647_ (.Y(_0116_),
    .A(\da[4] ));
 sg13g2_inv_1 _0648_ (.Y(_0117_),
    .A(\da[3] ));
 sg13g2_inv_1 _0649_ (.Y(_0118_),
    .A(\da[2] ));
 sg13g2_inv_1 _0650_ (.Y(_0119_),
    .A(\da[1] ));
 sg13g2_inv_1 _0651_ (.Y(_0120_),
    .A(\da[0] ));
 sg13g2_inv_1 _0652_ (.Y(_0121_),
    .A(net56));
 sg13g2_inv_1 _0653_ (.Y(_0122_),
    .A(\shiftedge.buff[3] ));
 sg13g2_inv_1 _0654_ (.Y(\resetsync.in ),
    .A(net3));
 sg13g2_inv_1 _0655_ (.Y(_0123_),
    .A(net54));
 sg13g2_and3_1 _0656_ (.X(\myring.inv_in[0] ),
    .A(net2),
    .B(net13),
    .C(\myring.inv_out[8] ));
 sg13g2_nand2b_1 _0657_ (.Y(_0124_),
    .B(net1),
    .A_N(net13));
 sg13g2_nand2b_1 _0658_ (.Y(internal_clock_unbuffered),
    .B(_0124_),
    .A_N(\myring.inv_in[0] ));
 sg13g2_nor2b_1 _0659_ (.A(net51),
    .B_N(_0003_),
    .Y(_0004_));
 sg13g2_nor2_1 _0660_ (.A(\clock_div[0] ),
    .B(\clock_div[1] ),
    .Y(_0125_));
 sg13g2_and2_1 _0661_ (.A(\clock_div[0] ),
    .B(\clock_div[1] ),
    .X(_0126_));
 sg13g2_nor3_1 _0662_ (.A(net51),
    .B(_0125_),
    .C(_0126_),
    .Y(_0005_));
 sg13g2_nor2_1 _0663_ (.A(\clock_div[2] ),
    .B(_0126_),
    .Y(_0127_));
 sg13g2_and2_1 _0664_ (.A(\clock_div[2] ),
    .B(_0126_),
    .X(_0128_));
 sg13g2_nor3_1 _0665_ (.A(net51),
    .B(_0127_),
    .C(_0128_),
    .Y(_0006_));
 sg13g2_and2_1 _0666_ (.A(\clock_div[3] ),
    .B(_0128_),
    .X(_0129_));
 sg13g2_nor2_1 _0667_ (.A(\clock_div[3] ),
    .B(_0128_),
    .Y(_0130_));
 sg13g2_nor3_1 _0668_ (.A(net51),
    .B(_0129_),
    .C(_0130_),
    .Y(_0007_));
 sg13g2_nor2b_1 _0669_ (.A(\stopedge.buff[3] ),
    .B_N(\stopedge.buff[1] ),
    .Y(_0131_));
 sg13g2_and4_1 _0670_ (.A(net57),
    .B(net77),
    .C(\stopedge.buff[2] ),
    .D(_0131_),
    .X(_0132_));
 sg13g2_nand2b_1 _0671_ (.Y(_0133_),
    .B(\db[8] ),
    .A_N(\cb[8] ));
 sg13g2_xnor2_1 _0672_ (.Y(_0134_),
    .A(\cb[5] ),
    .B(\db[5] ));
 sg13g2_nand2b_1 _0673_ (.Y(_0135_),
    .B(\db[6] ),
    .A_N(\cb[6] ));
 sg13g2_nand2_1 _0674_ (.Y(_0136_),
    .A(\cb[2] ),
    .B(_0109_));
 sg13g2_nor2b_1 _0675_ (.A(\db[8] ),
    .B_N(\cb[8] ),
    .Y(_0137_));
 sg13g2_nand2b_1 _0676_ (.Y(_0138_),
    .B(\cb[14] ),
    .A_N(\db[14] ));
 sg13g2_nand2b_1 _0677_ (.Y(_0139_),
    .B(\cb[10] ),
    .A_N(\db[10] ));
 sg13g2_a22oi_1 _0678_ (.Y(_0140_),
    .B1(\db[7] ),
    .B2(_0091_),
    .A2(_0101_),
    .A1(\cb[15] ));
 sg13g2_a22oi_1 _0679_ (.Y(_0141_),
    .B1(_0106_),
    .B2(\cb[12] ),
    .A2(_0102_),
    .A1(\cb[7] ));
 sg13g2_a22oi_1 _0680_ (.Y(_0142_),
    .B1(\db[1] ),
    .B2(_0094_),
    .A2(\db[9] ),
    .A1(_0090_));
 sg13g2_a22oi_1 _0681_ (.Y(_0143_),
    .B1(\db[13] ),
    .B2(_0087_),
    .A2(\db[14] ),
    .A1(_0086_));
 sg13g2_and4_1 _0682_ (.A(_0140_),
    .B(_0141_),
    .C(_0142_),
    .D(_0143_),
    .X(_0144_));
 sg13g2_a22oi_1 _0683_ (.Y(_0145_),
    .B1(\db[0] ),
    .B2(_0095_),
    .A2(_0107_),
    .A1(\cb[4] ));
 sg13g2_nand4_1 _0684_ (.B(_0136_),
    .C(_0144_),
    .A(_0135_),
    .Y(_0146_),
    .D(_0145_));
 sg13g2_a22oi_1 _0685_ (.Y(_0147_),
    .B1(_0111_),
    .B2(\cb[1] ),
    .A2(\db[15] ),
    .A1(_0085_));
 sg13g2_nand3_1 _0686_ (.B(_0139_),
    .C(_0147_),
    .A(_0133_),
    .Y(_0148_));
 sg13g2_a22oi_1 _0687_ (.Y(_0149_),
    .B1(_0110_),
    .B2(\cb[9] ),
    .A2(\db[12] ),
    .A1(_0088_));
 sg13g2_a22oi_1 _0688_ (.Y(_0150_),
    .B1(\db[2] ),
    .B2(_0093_),
    .A2(\db[4] ),
    .A1(_0092_));
 sg13g2_xnor2_1 _0689_ (.Y(_0151_),
    .A(\cb[11] ),
    .B(\db[11] ));
 sg13g2_nand4_1 _0690_ (.B(_0149_),
    .C(_0150_),
    .A(_0138_),
    .Y(_0152_),
    .D(_0151_));
 sg13g2_a22oi_1 _0691_ (.Y(_0153_),
    .B1(_0112_),
    .B2(\cb[0] ),
    .A2(\db[10] ),
    .A1(_0089_));
 sg13g2_a22oi_1 _0692_ (.Y(_0154_),
    .B1(_0104_),
    .B2(\cb[13] ),
    .A2(_0103_),
    .A1(\cb[6] ));
 sg13g2_xnor2_1 _0693_ (.Y(_0155_),
    .A(\cb[3] ),
    .B(\db[3] ));
 sg13g2_nand2_1 _0694_ (.Y(_0156_),
    .A(_0134_),
    .B(_0155_));
 sg13g2_nor4_1 _0695_ (.A(_0121_),
    .B(net76),
    .C(_0137_),
    .D(_0156_),
    .Y(_0157_));
 sg13g2_nand3_1 _0696_ (.B(_0154_),
    .C(_0157_),
    .A(_0153_),
    .Y(_0158_));
 sg13g2_nor4_2 _0697_ (.A(_0146_),
    .B(_0148_),
    .C(_0152_),
    .Y(_0159_),
    .D(_0158_));
 sg13g2_a21oi_2 _0698_ (.B1(_0159_),
    .Y(_0160_),
    .A2(_0132_),
    .A1(\stopedge.buff[0] ));
 sg13g2_and4_2 _0699_ (.A(\shiftedge.buff[1] ),
    .B(\shiftedge.buff[0] ),
    .C(_0122_),
    .D(\shiftedge.buff[2] ),
    .X(_0161_));
 sg13g2_nand4_1 _0700_ (.B(\shiftedge.buff[0] ),
    .C(_0122_),
    .A(\shiftedge.buff[1] ),
    .Y(_0162_),
    .D(\shiftedge.buff[2] ));
 sg13g2_nand2_1 _0701_ (.Y(_0163_),
    .A(done),
    .B(net24));
 sg13g2_a21oi_1 _0702_ (.A1(_0160_),
    .A2(_0163_),
    .Y(_0008_),
    .B1(net51));
 sg13g2_and2_2 _0703_ (.A(\shift_counter[1] ),
    .B(\shift_counter[0] ),
    .X(_0164_));
 sg13g2_nand2_1 _0704_ (.Y(_0165_),
    .A(\shift_counter[1] ),
    .B(\shift_counter[0] ));
 sg13g2_a22oi_1 _0705_ (.Y(_0166_),
    .B1(net30),
    .B2(net40),
    .A2(_0160_),
    .A1(net57));
 sg13g2_nor2_1 _0706_ (.A(net51),
    .B(_0166_),
    .Y(_0009_));
 sg13g2_o21ai_1 _0707_ (.B1(net41),
    .Y(_0167_),
    .A1(\db[8] ),
    .A2(net24));
 sg13g2_a21oi_1 _0708_ (.A1(_0120_),
    .A2(net24),
    .Y(_0010_),
    .B1(_0167_));
 sg13g2_o21ai_1 _0709_ (.B1(net44),
    .Y(_0168_),
    .A1(\da[1] ),
    .A2(net29));
 sg13g2_a21oi_1 _0710_ (.A1(_0110_),
    .A2(net31),
    .Y(_0011_),
    .B1(_0168_));
 sg13g2_o21ai_1 _0711_ (.B1(net45),
    .Y(_0169_),
    .A1(\db[10] ),
    .A2(net25));
 sg13g2_a21oi_1 _0712_ (.A1(_0118_),
    .A2(net25),
    .Y(_0012_),
    .B1(_0169_));
 sg13g2_o21ai_1 _0713_ (.B1(net45),
    .Y(_0170_),
    .A1(\db[11] ),
    .A2(net25));
 sg13g2_a21oi_1 _0714_ (.A1(_0117_),
    .A2(net25),
    .Y(_0013_),
    .B1(_0170_));
 sg13g2_o21ai_1 _0715_ (.B1(net45),
    .Y(_0171_),
    .A1(\db[12] ),
    .A2(net25));
 sg13g2_a21oi_1 _0716_ (.A1(_0116_),
    .A2(net28),
    .Y(_0014_),
    .B1(_0171_));
 sg13g2_o21ai_1 _0717_ (.B1(net46),
    .Y(_0172_),
    .A1(\db[13] ),
    .A2(net26));
 sg13g2_a21oi_1 _0718_ (.A1(_0115_),
    .A2(net26),
    .Y(_0015_),
    .B1(_0172_));
 sg13g2_o21ai_1 _0719_ (.B1(net47),
    .Y(_0173_),
    .A1(\db[14] ),
    .A2(net27));
 sg13g2_a21oi_1 _0720_ (.A1(_0114_),
    .A2(net27),
    .Y(_0016_),
    .B1(_0173_));
 sg13g2_o21ai_1 _0721_ (.B1(net43),
    .Y(_0174_),
    .A1(\db[15] ),
    .A2(_0162_));
 sg13g2_a21oi_1 _0722_ (.A1(_0113_),
    .A2(net24),
    .Y(_0017_),
    .B1(_0174_));
 sg13g2_o21ai_1 _0723_ (.B1(net44),
    .Y(_0175_),
    .A1(\da[8] ),
    .A2(net31));
 sg13g2_a21oi_1 _0724_ (.A1(_0120_),
    .A2(net31),
    .Y(_0018_),
    .B1(_0175_));
 sg13g2_o21ai_1 _0725_ (.B1(net44),
    .Y(_0176_),
    .A1(\da[9] ),
    .A2(net31));
 sg13g2_a21oi_1 _0726_ (.A1(_0119_),
    .A2(net31),
    .Y(_0019_),
    .B1(_0176_));
 sg13g2_o21ai_1 _0727_ (.B1(net45),
    .Y(_0177_),
    .A1(\da[10] ),
    .A2(net32));
 sg13g2_a21oi_1 _0728_ (.A1(_0118_),
    .A2(net32),
    .Y(_0020_),
    .B1(_0177_));
 sg13g2_o21ai_1 _0729_ (.B1(net44),
    .Y(_0178_),
    .A1(\da[11] ),
    .A2(net32));
 sg13g2_a21oi_1 _0730_ (.A1(_0117_),
    .A2(net32),
    .Y(_0021_),
    .B1(_0178_));
 sg13g2_o21ai_1 _0731_ (.B1(net46),
    .Y(_0179_),
    .A1(\da[12] ),
    .A2(net34));
 sg13g2_a21oi_1 _0732_ (.A1(_0116_),
    .A2(net34),
    .Y(_0022_),
    .B1(_0179_));
 sg13g2_o21ai_1 _0733_ (.B1(net46),
    .Y(_0180_),
    .A1(\da[13] ),
    .A2(net34));
 sg13g2_a21oi_1 _0734_ (.A1(_0115_),
    .A2(net33),
    .Y(_0023_),
    .B1(_0180_));
 sg13g2_o21ai_1 _0735_ (.B1(net47),
    .Y(_0181_),
    .A1(\da[14] ),
    .A2(net33));
 sg13g2_a21oi_1 _0736_ (.A1(_0114_),
    .A2(net33),
    .Y(_0024_),
    .B1(_0181_));
 sg13g2_o21ai_1 _0737_ (.B1(net43),
    .Y(_0182_),
    .A1(\da[15] ),
    .A2(net30));
 sg13g2_a21oi_1 _0738_ (.A1(_0113_),
    .A2(net30),
    .Y(_0025_),
    .B1(_0182_));
 sg13g2_o21ai_1 _0739_ (.B1(net47),
    .Y(_0183_),
    .A1(net4),
    .A2(net26));
 sg13g2_a21oi_1 _0740_ (.A1(_0112_),
    .A2(net28),
    .Y(_0026_),
    .B1(_0183_));
 sg13g2_o21ai_1 _0741_ (.B1(net46),
    .Y(_0184_),
    .A1(net5),
    .A2(net26));
 sg13g2_a21oi_1 _0742_ (.A1(_0111_),
    .A2(net24),
    .Y(_0027_),
    .B1(_0184_));
 sg13g2_o21ai_1 _0743_ (.B1(net46),
    .Y(_0185_),
    .A1(net6),
    .A2(net26));
 sg13g2_a21oi_1 _0744_ (.A1(_0109_),
    .A2(net25),
    .Y(_0028_),
    .B1(_0185_));
 sg13g2_o21ai_1 _0745_ (.B1(net46),
    .Y(_0186_),
    .A1(net7),
    .A2(net26));
 sg13g2_a21oi_1 _0746_ (.A1(_0108_),
    .A2(net25),
    .Y(_0029_),
    .B1(_0186_));
 sg13g2_o21ai_1 _0747_ (.B1(net46),
    .Y(_0187_),
    .A1(net8),
    .A2(net26));
 sg13g2_a21oi_1 _0748_ (.A1(_0107_),
    .A2(net25),
    .Y(_0030_),
    .B1(_0187_));
 sg13g2_o21ai_1 _0749_ (.B1(net46),
    .Y(_0188_),
    .A1(net9),
    .A2(net26));
 sg13g2_a21oi_1 _0750_ (.A1(_0105_),
    .A2(net27),
    .Y(_0031_),
    .B1(_0188_));
 sg13g2_o21ai_1 _0751_ (.B1(net47),
    .Y(_0189_),
    .A1(net10),
    .A2(net27));
 sg13g2_a21oi_1 _0752_ (.A1(_0103_),
    .A2(net27),
    .Y(_0032_),
    .B1(_0189_));
 sg13g2_o21ai_1 _0753_ (.B1(net47),
    .Y(_0190_),
    .A1(net11),
    .A2(net27));
 sg13g2_a21oi_1 _0754_ (.A1(_0102_),
    .A2(net27),
    .Y(_0033_),
    .B1(_0190_));
 sg13g2_o21ai_1 _0755_ (.B1(net44),
    .Y(_0191_),
    .A1(\db[8] ),
    .A2(net32));
 sg13g2_a21oi_1 _0756_ (.A1(_0112_),
    .A2(net31),
    .Y(_0034_),
    .B1(_0191_));
 sg13g2_o21ai_1 _0757_ (.B1(net41),
    .Y(_0192_),
    .A1(\db[9] ),
    .A2(net29));
 sg13g2_a21oi_1 _0758_ (.A1(_0111_),
    .A2(net29),
    .Y(_0035_),
    .B1(_0192_));
 sg13g2_o21ai_1 _0759_ (.B1(net44),
    .Y(_0193_),
    .A1(\db[10] ),
    .A2(net31));
 sg13g2_a21oi_1 _0760_ (.A1(_0109_),
    .A2(net31),
    .Y(_0036_),
    .B1(_0193_));
 sg13g2_o21ai_1 _0761_ (.B1(net44),
    .Y(_0194_),
    .A1(\db[11] ),
    .A2(net32));
 sg13g2_a21oi_1 _0762_ (.A1(_0108_),
    .A2(net32),
    .Y(_0037_),
    .B1(_0194_));
 sg13g2_o21ai_1 _0763_ (.B1(net44),
    .Y(_0195_),
    .A1(\db[12] ),
    .A2(net33));
 sg13g2_a21oi_1 _0764_ (.A1(_0107_),
    .A2(net33),
    .Y(_0038_),
    .B1(_0195_));
 sg13g2_o21ai_1 _0765_ (.B1(net47),
    .Y(_0196_),
    .A1(\db[13] ),
    .A2(net33));
 sg13g2_a21oi_1 _0766_ (.A1(_0105_),
    .A2(net33),
    .Y(_0039_),
    .B1(_0196_));
 sg13g2_o21ai_1 _0767_ (.B1(net43),
    .Y(_0197_),
    .A1(\db[14] ),
    .A2(net30));
 sg13g2_a21oi_1 _0768_ (.A1(_0103_),
    .A2(net33),
    .Y(_0040_),
    .B1(_0197_));
 sg13g2_o21ai_1 _0769_ (.B1(net42),
    .Y(_0198_),
    .A1(\db[15] ),
    .A2(net30));
 sg13g2_a21oi_1 _0770_ (.A1(_0102_),
    .A2(net30),
    .Y(_0041_),
    .B1(_0198_));
 sg13g2_nand2_1 _0771_ (.Y(_0199_),
    .A(\db[0] ),
    .B(net76));
 sg13g2_xnor2_1 _0772_ (.Y(_0200_),
    .A(_0120_),
    .B(_0199_));
 sg13g2_nor2_1 _0773_ (.A(net57),
    .B(net24),
    .Y(_0201_));
 sg13g2_nand2_1 _0774_ (.Y(_0202_),
    .A(net49),
    .B(net29));
 sg13g2_o21ai_1 _0775_ (.B1(net23),
    .Y(_0203_),
    .A1(\cb[8] ),
    .A2(net40));
 sg13g2_a21oi_1 _0776_ (.A1(net40),
    .A2(_0200_),
    .Y(_0204_),
    .B1(_0203_));
 sg13g2_nor2_2 _0777_ (.A(net57),
    .B(net29),
    .Y(_0205_));
 sg13g2_nand2_1 _0778_ (.Y(_0206_),
    .A(net49),
    .B(net24));
 sg13g2_a221oi_1 _0779_ (.B2(\ca[0] ),
    .C1(_0204_),
    .B1(_0205_),
    .A1(net55),
    .Y(_0207_),
    .A2(_0000_));
 sg13g2_nor2_1 _0780_ (.A(net50),
    .B(_0207_),
    .Y(_0042_));
 sg13g2_nand2_1 _0781_ (.Y(_0208_),
    .A(\db[0] ),
    .B(\da[0] ));
 sg13g2_nand2_1 _0782_ (.Y(_0209_),
    .A(\db[1] ),
    .B(\da[1] ));
 sg13g2_xnor2_1 _0783_ (.Y(_0210_),
    .A(\db[1] ),
    .B(\da[1] ));
 sg13g2_nand3_1 _0784_ (.B(\ca[0] ),
    .C(net56),
    .A(\ca[1] ),
    .Y(_0211_));
 sg13g2_nand2_1 _0785_ (.Y(_0212_),
    .A(net43),
    .B(_0211_));
 sg13g2_a21oi_1 _0786_ (.A1(\ca[0] ),
    .A2(net56),
    .Y(_0213_),
    .B1(\ca[1] ));
 sg13g2_nor2_2 _0787_ (.A(net40),
    .B(net19),
    .Y(_0214_));
 sg13g2_a21oi_1 _0788_ (.A1(\cb[9] ),
    .A2(net37),
    .Y(_0215_),
    .B1(net20));
 sg13g2_xnor2_1 _0789_ (.Y(_0216_),
    .A(_0208_),
    .B(_0210_));
 sg13g2_o21ai_1 _0790_ (.B1(net38),
    .Y(_0217_),
    .A1(\da[1] ),
    .A2(net76));
 sg13g2_a21o_1 _0791_ (.A2(_0216_),
    .A1(net76),
    .B1(_0217_),
    .X(_0218_));
 sg13g2_a221oi_1 _0792_ (.B2(_0218_),
    .C1(_0212_),
    .B1(_0215_),
    .A1(net20),
    .Y(_0043_),
    .A2(_0213_));
 sg13g2_nor3_1 _0793_ (.A(\cb[10] ),
    .B(net40),
    .C(net20),
    .Y(_0219_));
 sg13g2_nand3_1 _0794_ (.B(\ca[1] ),
    .C(\ca[0] ),
    .A(\ca[2] ),
    .Y(_0220_));
 sg13g2_a21o_1 _0795_ (.A2(\ca[0] ),
    .A1(\ca[1] ),
    .B1(\ca[2] ),
    .X(_0221_));
 sg13g2_a21oi_1 _0796_ (.A1(_0220_),
    .A2(_0221_),
    .Y(_0222_),
    .B1(net49));
 sg13g2_o21ai_1 _0797_ (.B1(net41),
    .Y(_0223_),
    .A1(\ca[2] ),
    .A2(net17));
 sg13g2_o21ai_1 _0798_ (.B1(_0209_),
    .Y(_0224_),
    .A1(_0208_),
    .A2(_0210_));
 sg13g2_nand2_1 _0799_ (.Y(_0225_),
    .A(\db[2] ),
    .B(\da[2] ));
 sg13g2_xnor2_1 _0800_ (.Y(_0226_),
    .A(\db[2] ),
    .B(\da[2] ));
 sg13g2_nand2b_1 _0801_ (.Y(_0227_),
    .B(_0224_),
    .A_N(_0226_));
 sg13g2_nand2b_1 _0802_ (.Y(_0228_),
    .B(_0226_),
    .A_N(_0224_));
 sg13g2_nand3_1 _0803_ (.B(_0227_),
    .C(_0228_),
    .A(net74),
    .Y(_0229_));
 sg13g2_o21ai_1 _0804_ (.B1(_0229_),
    .Y(_0230_),
    .A1(_0118_),
    .A2(net74));
 sg13g2_nor3_1 _0805_ (.A(net35),
    .B(net20),
    .C(_0230_),
    .Y(_0231_));
 sg13g2_nor4_1 _0806_ (.A(_0219_),
    .B(_0222_),
    .C(_0223_),
    .D(_0231_),
    .Y(_0044_));
 sg13g2_nor2_1 _0807_ (.A(\db[3] ),
    .B(\da[3] ),
    .Y(_0232_));
 sg13g2_nand2_1 _0808_ (.Y(_0233_),
    .A(\db[3] ),
    .B(\da[3] ));
 sg13g2_xnor2_1 _0809_ (.Y(_0234_),
    .A(\db[3] ),
    .B(\da[3] ));
 sg13g2_nand2_1 _0810_ (.Y(_0235_),
    .A(_0225_),
    .B(_0227_));
 sg13g2_xor2_1 _0811_ (.B(_0235_),
    .A(_0234_),
    .X(_0236_));
 sg13g2_o21ai_1 _0812_ (.B1(net38),
    .Y(_0237_),
    .A1(\da[3] ),
    .A2(net74));
 sg13g2_a21o_1 _0813_ (.A2(_0236_),
    .A1(net74),
    .B1(_0237_),
    .X(_0238_));
 sg13g2_a21oi_1 _0814_ (.A1(\cb[11] ),
    .A2(net35),
    .Y(_0239_),
    .B1(net20));
 sg13g2_o21ai_1 _0815_ (.B1(net41),
    .Y(_0240_),
    .A1(\ca[3] ),
    .A2(net17));
 sg13g2_and4_2 _0816_ (.A(\ca[3] ),
    .B(\ca[2] ),
    .C(\ca[1] ),
    .D(\ca[0] ),
    .X(_0241_));
 sg13g2_xor2_1 _0817_ (.B(_0220_),
    .A(\ca[3] ),
    .X(_0242_));
 sg13g2_a221oi_1 _0818_ (.B2(net55),
    .C1(_0240_),
    .B1(_0242_),
    .A1(_0238_),
    .Y(_0045_),
    .A2(_0239_));
 sg13g2_nor2_1 _0819_ (.A(_0226_),
    .B(_0234_),
    .Y(_0243_));
 sg13g2_o21ai_1 _0820_ (.B1(_0233_),
    .Y(_0244_),
    .A1(_0225_),
    .A2(_0232_));
 sg13g2_a21oi_1 _0821_ (.A1(_0224_),
    .A2(_0243_),
    .Y(_0245_),
    .B1(_0244_));
 sg13g2_a21o_1 _0822_ (.A2(_0243_),
    .A1(_0224_),
    .B1(_0244_),
    .X(_0246_));
 sg13g2_nand2_1 _0823_ (.Y(_0247_),
    .A(\db[4] ),
    .B(\da[4] ));
 sg13g2_xor2_1 _0824_ (.B(\da[4] ),
    .A(\db[4] ),
    .X(_0248_));
 sg13g2_nand2_1 _0825_ (.Y(_0249_),
    .A(_0246_),
    .B(_0248_));
 sg13g2_xnor2_1 _0826_ (.Y(_0250_),
    .A(_0246_),
    .B(_0248_));
 sg13g2_o21ai_1 _0827_ (.B1(net38),
    .Y(_0251_),
    .A1(\da[4] ),
    .A2(net75));
 sg13g2_a21o_1 _0828_ (.A2(_0250_),
    .A1(net75),
    .B1(_0251_),
    .X(_0252_));
 sg13g2_a21oi_1 _0829_ (.A1(\cb[12] ),
    .A2(net36),
    .Y(_0253_),
    .B1(net21));
 sg13g2_o21ai_1 _0830_ (.B1(net43),
    .Y(_0254_),
    .A1(\ca[4] ),
    .A2(net18));
 sg13g2_xnor2_1 _0831_ (.Y(_0255_),
    .A(\ca[4] ),
    .B(_0241_));
 sg13g2_a221oi_1 _0832_ (.B2(net56),
    .C1(_0254_),
    .B1(_0255_),
    .A1(_0252_),
    .Y(_0046_),
    .A2(_0253_));
 sg13g2_nor2_1 _0833_ (.A(\db[5] ),
    .B(\da[5] ),
    .Y(_0256_));
 sg13g2_and2_1 _0834_ (.A(_0247_),
    .B(_0249_),
    .X(_0257_));
 sg13g2_nand2_1 _0835_ (.Y(_0258_),
    .A(\db[5] ),
    .B(\da[5] ));
 sg13g2_nor2b_1 _0836_ (.A(_0256_),
    .B_N(_0258_),
    .Y(_0259_));
 sg13g2_xor2_1 _0837_ (.B(_0259_),
    .A(_0257_),
    .X(_0260_));
 sg13g2_o21ai_1 _0838_ (.B1(net39),
    .Y(_0261_),
    .A1(\da[5] ),
    .A2(net77));
 sg13g2_a21oi_1 _0839_ (.A1(net78),
    .A2(_0260_),
    .Y(_0262_),
    .B1(_0261_));
 sg13g2_a21oi_1 _0840_ (.A1(\cb[13] ),
    .A2(net37),
    .Y(_0263_),
    .B1(_0262_));
 sg13g2_nand3_1 _0841_ (.B(\ca[4] ),
    .C(_0241_),
    .A(\ca[5] ),
    .Y(_0264_));
 sg13g2_a21o_1 _0842_ (.A2(_0241_),
    .A1(\ca[4] ),
    .B1(\ca[5] ),
    .X(_0265_));
 sg13g2_nand2_1 _0843_ (.Y(_0266_),
    .A(_0264_),
    .B(_0265_));
 sg13g2_o21ai_1 _0844_ (.B1(net42),
    .Y(_0267_),
    .A1(\ca[5] ),
    .A2(net18));
 sg13g2_a221oi_1 _0845_ (.B2(net58),
    .C1(_0267_),
    .B1(_0266_),
    .A1(_0201_),
    .Y(_0047_),
    .A2(_0263_));
 sg13g2_nor2_1 _0846_ (.A(\db[6] ),
    .B(\da[6] ),
    .Y(_0268_));
 sg13g2_nand2_1 _0847_ (.Y(_0269_),
    .A(\db[6] ),
    .B(\da[6] ));
 sg13g2_xor2_1 _0848_ (.B(\da[6] ),
    .A(\db[6] ),
    .X(_0270_));
 sg13g2_a21oi_1 _0849_ (.A1(_0247_),
    .A2(_0258_),
    .Y(_0271_),
    .B1(_0256_));
 sg13g2_a21o_1 _0850_ (.A2(_0258_),
    .A1(_0257_),
    .B1(_0256_),
    .X(_0272_));
 sg13g2_xor2_1 _0851_ (.B(_0272_),
    .A(_0270_),
    .X(_0273_));
 sg13g2_o21ai_1 _0852_ (.B1(net39),
    .Y(_0274_),
    .A1(\da[6] ),
    .A2(net78));
 sg13g2_a21o_1 _0853_ (.A2(_0273_),
    .A1(net78),
    .B1(_0274_),
    .X(_0275_));
 sg13g2_a21oi_1 _0854_ (.A1(\cb[14] ),
    .A2(net36),
    .Y(_0276_),
    .B1(net21));
 sg13g2_o21ai_1 _0855_ (.B1(net42),
    .Y(_0277_),
    .A1(\ca[6] ),
    .A2(net18));
 sg13g2_nand4_1 _0856_ (.B(\ca[5] ),
    .C(\ca[4] ),
    .A(\ca[6] ),
    .Y(_0278_),
    .D(_0241_));
 sg13g2_xor2_1 _0857_ (.B(_0264_),
    .A(\ca[6] ),
    .X(_0279_));
 sg13g2_a221oi_1 _0858_ (.B2(net58),
    .C1(_0277_),
    .B1(_0279_),
    .A1(_0275_),
    .Y(_0048_),
    .A2(_0276_));
 sg13g2_xor2_1 _0859_ (.B(\da[7] ),
    .A(\db[7] ),
    .X(_0280_));
 sg13g2_o21ai_1 _0860_ (.B1(_0269_),
    .Y(_0281_),
    .A1(_0268_),
    .A2(_0272_));
 sg13g2_xnor2_1 _0861_ (.Y(_0282_),
    .A(_0280_),
    .B(_0281_));
 sg13g2_o21ai_1 _0862_ (.B1(net39),
    .Y(_0283_),
    .A1(\da[7] ),
    .A2(net77));
 sg13g2_a21oi_1 _0863_ (.A1(net77),
    .A2(_0282_),
    .Y(_0284_),
    .B1(_0283_));
 sg13g2_a21oi_1 _0864_ (.A1(\cb[15] ),
    .A2(net36),
    .Y(_0285_),
    .B1(_0284_));
 sg13g2_nor2_1 _0865_ (.A(_0100_),
    .B(_0278_),
    .Y(_0286_));
 sg13g2_xnor2_1 _0866_ (.Y(_0287_),
    .A(_0100_),
    .B(_0278_));
 sg13g2_o21ai_1 _0867_ (.B1(net42),
    .Y(_0288_),
    .A1(\ca[7] ),
    .A2(net18));
 sg13g2_a221oi_1 _0868_ (.B2(net56),
    .C1(_0288_),
    .B1(_0287_),
    .A1(net23),
    .Y(_0049_),
    .A2(_0285_));
 sg13g2_and2_1 _0869_ (.A(_0270_),
    .B(_0280_),
    .X(_0289_));
 sg13g2_nand3_1 _0870_ (.B(_0259_),
    .C(_0289_),
    .A(_0248_),
    .Y(_0290_));
 sg13g2_a22oi_1 _0871_ (.Y(_0291_),
    .B1(\da[6] ),
    .B2(\db[6] ),
    .A2(\da[7] ),
    .A1(\db[7] ));
 sg13g2_a21oi_1 _0872_ (.A1(_0102_),
    .A2(_0113_),
    .Y(_0292_),
    .B1(_0291_));
 sg13g2_a21oi_1 _0873_ (.A1(_0271_),
    .A2(_0289_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_o21ai_1 _0874_ (.B1(_0293_),
    .Y(_0294_),
    .A1(_0245_),
    .A2(_0290_));
 sg13g2_nand2_1 _0875_ (.Y(_0295_),
    .A(\db[8] ),
    .B(\da[8] ));
 sg13g2_xor2_1 _0876_ (.B(\da[8] ),
    .A(\db[8] ),
    .X(_0296_));
 sg13g2_nand2_1 _0877_ (.Y(_0297_),
    .A(_0294_),
    .B(_0296_));
 sg13g2_xnor2_1 _0878_ (.Y(_0298_),
    .A(_0294_),
    .B(_0296_));
 sg13g2_o21ai_1 _0879_ (.B1(net38),
    .Y(_0299_),
    .A1(\da[8] ),
    .A2(net76));
 sg13g2_a21o_1 _0880_ (.A2(_0298_),
    .A1(net74),
    .B1(_0299_),
    .X(_0300_));
 sg13g2_a21oi_1 _0881_ (.A1(\ca[0] ),
    .A2(net37),
    .Y(_0301_),
    .B1(net20));
 sg13g2_o21ai_1 _0882_ (.B1(net41),
    .Y(_0302_),
    .A1(\ca[8] ),
    .A2(net17));
 sg13g2_nor3_2 _0883_ (.A(_0099_),
    .B(_0100_),
    .C(_0278_),
    .Y(_0303_));
 sg13g2_xnor2_1 _0884_ (.Y(_0304_),
    .A(\ca[8] ),
    .B(_0286_));
 sg13g2_a221oi_1 _0885_ (.B2(net56),
    .C1(_0302_),
    .B1(_0304_),
    .A1(_0300_),
    .Y(_0050_),
    .A2(_0301_));
 sg13g2_nand2_1 _0886_ (.Y(_0305_),
    .A(_0295_),
    .B(_0297_));
 sg13g2_nor2_1 _0887_ (.A(\db[9] ),
    .B(\da[9] ),
    .Y(_0306_));
 sg13g2_or2_1 _0888_ (.X(_0307_),
    .B(\da[9] ),
    .A(\db[9] ));
 sg13g2_nand2_1 _0889_ (.Y(_0308_),
    .A(\db[9] ),
    .B(\da[9] ));
 sg13g2_nand2_1 _0890_ (.Y(_0309_),
    .A(_0307_),
    .B(_0308_));
 sg13g2_xor2_1 _0891_ (.B(_0309_),
    .A(_0305_),
    .X(_0310_));
 sg13g2_o21ai_1 _0892_ (.B1(net38),
    .Y(_0311_),
    .A1(\da[9] ),
    .A2(net74));
 sg13g2_a21oi_1 _0893_ (.A1(net74),
    .A2(_0310_),
    .Y(_0312_),
    .B1(_0311_));
 sg13g2_a21o_1 _0894_ (.A2(net35),
    .A1(\ca[1] ),
    .B1(_0312_),
    .X(_0313_));
 sg13g2_nand2_1 _0895_ (.Y(_0314_),
    .A(\ca[9] ),
    .B(_0303_));
 sg13g2_nand2_1 _0896_ (.Y(_0315_),
    .A(net55),
    .B(_0314_));
 sg13g2_a21oi_1 _0897_ (.A1(net55),
    .A2(_0303_),
    .Y(_0316_),
    .B1(\ca[9] ));
 sg13g2_a21oi_1 _0898_ (.A1(net17),
    .A2(_0315_),
    .Y(_0317_),
    .B1(_0316_));
 sg13g2_a21oi_1 _0899_ (.A1(net23),
    .A2(_0313_),
    .Y(_0318_),
    .B1(_0317_));
 sg13g2_nor2_1 _0900_ (.A(net53),
    .B(_0318_),
    .Y(_0051_));
 sg13g2_and2_1 _0901_ (.A(\db[10] ),
    .B(\da[10] ),
    .X(_0319_));
 sg13g2_xor2_1 _0902_ (.B(\da[10] ),
    .A(\db[10] ),
    .X(_0320_));
 sg13g2_o21ai_1 _0903_ (.B1(_0308_),
    .Y(_0321_),
    .A1(_0295_),
    .A2(_0306_));
 sg13g2_nand3_1 _0904_ (.B(_0296_),
    .C(_0307_),
    .A(_0294_),
    .Y(_0322_));
 sg13g2_nand2b_1 _0905_ (.Y(_0323_),
    .B(_0322_),
    .A_N(_0321_));
 sg13g2_xnor2_1 _0906_ (.Y(_0324_),
    .A(_0320_),
    .B(_0323_));
 sg13g2_o21ai_1 _0907_ (.B1(net38),
    .Y(_0325_),
    .A1(\da[10] ),
    .A2(net74));
 sg13g2_a21oi_1 _0908_ (.A1(net75),
    .A2(_0324_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_a21oi_1 _0909_ (.A1(\ca[2] ),
    .A2(net35),
    .Y(_0327_),
    .B1(net20));
 sg13g2_nor2b_1 _0910_ (.A(_0326_),
    .B_N(_0327_),
    .Y(_0328_));
 sg13g2_nor3_1 _0911_ (.A(_0098_),
    .B(net49),
    .C(_0314_),
    .Y(_0329_));
 sg13g2_a21oi_1 _0912_ (.A1(net17),
    .A2(_0315_),
    .Y(_0330_),
    .B1(\ca[10] ));
 sg13g2_nor4_1 _0913_ (.A(net54),
    .B(_0328_),
    .C(_0329_),
    .D(_0330_),
    .Y(_0052_));
 sg13g2_nand2_1 _0914_ (.Y(_0331_),
    .A(\db[11] ),
    .B(\da[11] ));
 sg13g2_xor2_1 _0915_ (.B(\da[11] ),
    .A(\db[11] ),
    .X(_0332_));
 sg13g2_a21oi_1 _0916_ (.A1(_0320_),
    .A2(_0323_),
    .Y(_0333_),
    .B1(_0319_));
 sg13g2_xor2_1 _0917_ (.B(_0333_),
    .A(_0332_),
    .X(_0334_));
 sg13g2_o21ai_1 _0918_ (.B1(net38),
    .Y(_0335_),
    .A1(\da[11] ),
    .A2(net75));
 sg13g2_a21oi_2 _0919_ (.B1(_0335_),
    .Y(_0336_),
    .A2(_0334_),
    .A1(net75));
 sg13g2_a21oi_1 _0920_ (.A1(\ca[3] ),
    .A2(net35),
    .Y(_0337_),
    .B1(net20));
 sg13g2_nor2b_1 _0921_ (.A(_0336_),
    .B_N(_0337_),
    .Y(_0338_));
 sg13g2_nor3_1 _0922_ (.A(\ca[11] ),
    .B(net23),
    .C(_0329_),
    .Y(_0339_));
 sg13g2_and2_1 _0923_ (.A(\ca[11] ),
    .B(_0329_),
    .X(_0340_));
 sg13g2_nor4_1 _0924_ (.A(net53),
    .B(_0338_),
    .C(_0339_),
    .D(_0340_),
    .Y(_0053_));
 sg13g2_and2_1 _0925_ (.A(_0320_),
    .B(_0332_),
    .X(_0341_));
 sg13g2_and4_1 _0926_ (.A(_0296_),
    .B(_0307_),
    .C(_0308_),
    .D(_0341_),
    .X(_0342_));
 sg13g2_nand2_1 _0927_ (.Y(_0343_),
    .A(_0321_),
    .B(_0341_));
 sg13g2_o21ai_1 _0928_ (.B1(_0319_),
    .Y(_0344_),
    .A1(\db[11] ),
    .A2(\da[11] ));
 sg13g2_nand3_1 _0929_ (.B(_0343_),
    .C(_0344_),
    .A(_0331_),
    .Y(_0345_));
 sg13g2_a21o_2 _0930_ (.A2(_0342_),
    .A1(_0294_),
    .B1(_0345_),
    .X(_0346_));
 sg13g2_and2_1 _0931_ (.A(\db[12] ),
    .B(\da[12] ),
    .X(_0347_));
 sg13g2_or2_1 _0932_ (.X(_0348_),
    .B(\da[12] ),
    .A(\db[12] ));
 sg13g2_nand2b_1 _0933_ (.Y(_0349_),
    .B(_0348_),
    .A_N(_0347_));
 sg13g2_xor2_1 _0934_ (.B(_0349_),
    .A(_0346_),
    .X(_0350_));
 sg13g2_o21ai_1 _0935_ (.B1(net39),
    .Y(_0351_),
    .A1(\da[12] ),
    .A2(net78));
 sg13g2_a21o_1 _0936_ (.A2(_0350_),
    .A1(net78),
    .B1(_0351_),
    .X(_0352_));
 sg13g2_a21oi_1 _0937_ (.A1(\ca[4] ),
    .A2(net36),
    .Y(_0353_),
    .B1(net21));
 sg13g2_o21ai_1 _0938_ (.B1(net42),
    .Y(_0354_),
    .A1(\ca[12] ),
    .A2(net18));
 sg13g2_nand4_1 _0939_ (.B(\ca[10] ),
    .C(\ca[9] ),
    .A(\ca[11] ),
    .Y(_0355_),
    .D(_0303_));
 sg13g2_or2_1 _0940_ (.X(_0356_),
    .B(_0355_),
    .A(_0097_));
 sg13g2_xnor2_1 _0941_ (.Y(_0357_),
    .A(_0097_),
    .B(_0355_));
 sg13g2_a221oi_1 _0942_ (.B2(net58),
    .C1(_0354_),
    .B1(_0357_),
    .A1(_0352_),
    .Y(_0054_),
    .A2(_0353_));
 sg13g2_or2_1 _0943_ (.X(_0358_),
    .B(\da[13] ),
    .A(\db[13] ));
 sg13g2_and2_1 _0944_ (.A(\db[13] ),
    .B(\da[13] ),
    .X(_0359_));
 sg13g2_xnor2_1 _0945_ (.Y(_0360_),
    .A(\db[13] ),
    .B(\da[13] ));
 sg13g2_a21oi_1 _0946_ (.A1(_0346_),
    .A2(_0348_),
    .Y(_0361_),
    .B1(_0347_));
 sg13g2_xnor2_1 _0947_ (.Y(_0362_),
    .A(_0360_),
    .B(_0361_));
 sg13g2_o21ai_1 _0948_ (.B1(net39),
    .Y(_0363_),
    .A1(\da[13] ),
    .A2(net78));
 sg13g2_a21oi_1 _0949_ (.A1(net78),
    .A2(_0362_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_a21oi_1 _0950_ (.A1(\ca[5] ),
    .A2(net36),
    .Y(_0365_),
    .B1(_0364_));
 sg13g2_nor2_1 _0951_ (.A(_0096_),
    .B(_0356_),
    .Y(_0366_));
 sg13g2_xnor2_1 _0952_ (.Y(_0367_),
    .A(_0096_),
    .B(_0356_));
 sg13g2_o21ai_1 _0953_ (.B1(net42),
    .Y(_0368_),
    .A1(\ca[13] ),
    .A2(net18));
 sg13g2_a221oi_1 _0954_ (.B2(net57),
    .C1(_0368_),
    .B1(_0367_),
    .A1(net23),
    .Y(_0055_),
    .A2(_0365_));
 sg13g2_nand2_1 _0955_ (.Y(_0369_),
    .A(\db[14] ),
    .B(\da[14] ));
 sg13g2_xnor2_1 _0956_ (.Y(_0370_),
    .A(\db[14] ),
    .B(\da[14] ));
 sg13g2_nor2_1 _0957_ (.A(_0349_),
    .B(_0360_),
    .Y(_0371_));
 sg13g2_a221oi_1 _0958_ (.B2(_0346_),
    .C1(_0359_),
    .B1(_0371_),
    .A1(_0347_),
    .Y(_0372_),
    .A2(_0358_));
 sg13g2_xnor2_1 _0959_ (.Y(_0373_),
    .A(_0370_),
    .B(_0372_));
 sg13g2_o21ai_1 _0960_ (.B1(net39),
    .Y(_0374_),
    .A1(\da[14] ),
    .A2(net77));
 sg13g2_a21o_1 _0961_ (.A2(_0373_),
    .A1(net77),
    .B1(_0374_),
    .X(_0375_));
 sg13g2_a21oi_1 _0962_ (.A1(\ca[6] ),
    .A2(net36),
    .Y(_0376_),
    .B1(net21));
 sg13g2_o21ai_1 _0963_ (.B1(net42),
    .Y(_0377_),
    .A1(\ca[14] ),
    .A2(net18));
 sg13g2_nand2_1 _0964_ (.Y(_0378_),
    .A(\ca[14] ),
    .B(_0366_));
 sg13g2_xnor2_1 _0965_ (.Y(_0379_),
    .A(\ca[14] ),
    .B(_0366_));
 sg13g2_a221oi_1 _0966_ (.B2(net58),
    .C1(_0377_),
    .B1(_0379_),
    .A1(_0375_),
    .Y(_0056_),
    .A2(_0376_));
 sg13g2_o21ai_1 _0967_ (.B1(_0369_),
    .Y(_0380_),
    .A1(_0370_),
    .A2(_0372_));
 sg13g2_xor2_1 _0968_ (.B(\da[15] ),
    .A(\db[15] ),
    .X(_0381_));
 sg13g2_xnor2_1 _0969_ (.Y(_0382_),
    .A(_0380_),
    .B(_0381_));
 sg13g2_o21ai_1 _0970_ (.B1(net38),
    .Y(_0383_),
    .A1(\da[15] ),
    .A2(net77));
 sg13g2_a21oi_1 _0971_ (.A1(net77),
    .A2(_0382_),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_o21ai_1 _0972_ (.B1(net49),
    .Y(_0385_),
    .A1(_0100_),
    .A2(net40));
 sg13g2_xor2_1 _0973_ (.B(_0378_),
    .A(\ca[15] ),
    .X(_0386_));
 sg13g2_a21oi_1 _0974_ (.A1(net57),
    .A2(_0386_),
    .Y(_0387_),
    .B1(_0205_));
 sg13g2_o21ai_1 _0975_ (.B1(_0387_),
    .Y(_0388_),
    .A1(_0384_),
    .A2(_0385_));
 sg13g2_nand2_1 _0976_ (.Y(_0389_),
    .A(\ca[15] ),
    .B(_0205_));
 sg13g2_a21oi_1 _0977_ (.A1(_0388_),
    .A2(_0389_),
    .Y(_0057_),
    .B1(net51));
 sg13g2_nand2_1 _0978_ (.Y(_0390_),
    .A(\cb[0] ),
    .B(_0205_));
 sg13g2_a22oi_1 _0979_ (.Y(_0391_),
    .B1(_0214_),
    .B2(\ca[8] ),
    .A2(_0001_),
    .A1(net56));
 sg13g2_a21oi_1 _0980_ (.A1(_0390_),
    .A2(_0391_),
    .Y(_0058_),
    .B1(net53));
 sg13g2_nand2_1 _0981_ (.Y(_0392_),
    .A(\cb[1] ),
    .B(\cb[0] ));
 sg13g2_a21o_1 _0982_ (.A2(_0392_),
    .A1(net55),
    .B1(_0205_),
    .X(_0393_));
 sg13g2_nand3_1 _0983_ (.B(net55),
    .C(_0392_),
    .A(\cb[0] ),
    .Y(_0394_));
 sg13g2_nand2_1 _0984_ (.Y(_0395_),
    .A(\ca[9] ),
    .B(net49));
 sg13g2_o21ai_1 _0985_ (.B1(_0394_),
    .Y(_0396_),
    .A1(net40),
    .A2(_0395_));
 sg13g2_a22oi_1 _0986_ (.Y(_0397_),
    .B1(_0396_),
    .B2(net17),
    .A2(_0393_),
    .A1(\cb[1] ));
 sg13g2_nor2_1 _0987_ (.A(net50),
    .B(_0397_),
    .Y(_0059_));
 sg13g2_and2_1 _0988_ (.A(_0093_),
    .B(_0393_),
    .X(_0398_));
 sg13g2_a21oi_1 _0989_ (.A1(\ca[10] ),
    .A2(net36),
    .Y(_0399_),
    .B1(net21));
 sg13g2_nor3_2 _0990_ (.A(_0093_),
    .B(net49),
    .C(_0392_),
    .Y(_0400_));
 sg13g2_nor4_1 _0991_ (.A(net52),
    .B(_0398_),
    .C(_0399_),
    .D(_0400_),
    .Y(_0060_));
 sg13g2_and2_1 _0992_ (.A(\cb[3] ),
    .B(_0400_),
    .X(_0401_));
 sg13g2_xor2_1 _0993_ (.B(_0400_),
    .A(\cb[3] ),
    .X(_0402_));
 sg13g2_a22oi_1 _0994_ (.Y(_0403_),
    .B1(_0402_),
    .B2(net19),
    .A2(net16),
    .A1(\ca[11] ));
 sg13g2_nor2_1 _0995_ (.A(net50),
    .B(_0403_),
    .Y(_0061_));
 sg13g2_nand4_1 _0996_ (.B(\cb[2] ),
    .C(\cb[1] ),
    .A(\cb[3] ),
    .Y(_0404_),
    .D(\cb[0] ));
 sg13g2_nand2b_1 _0997_ (.Y(_0405_),
    .B(_0404_),
    .A_N(\cb[4] ));
 sg13g2_a21oi_1 _0998_ (.A1(\cb[4] ),
    .A2(_0401_),
    .Y(_0406_),
    .B1(net23));
 sg13g2_nor3_1 _0999_ (.A(_0097_),
    .B(net57),
    .C(net40),
    .Y(_0407_));
 sg13g2_a21oi_1 _1000_ (.A1(_0405_),
    .A2(_0406_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_o21ai_1 _1001_ (.B1(net42),
    .Y(_0409_),
    .A1(\cb[4] ),
    .A2(net18));
 sg13g2_nor2_1 _1002_ (.A(_0408_),
    .B(_0409_),
    .Y(_0062_));
 sg13g2_nor2b_1 _1003_ (.A(\cb[5] ),
    .B_N(_0406_),
    .Y(_0410_));
 sg13g2_and3_1 _1004_ (.X(_0411_),
    .A(\cb[5] ),
    .B(\cb[4] ),
    .C(_0401_));
 sg13g2_a21oi_1 _1005_ (.A1(\ca[13] ),
    .A2(net36),
    .Y(_0412_),
    .B1(net19));
 sg13g2_nor4_1 _1006_ (.A(net52),
    .B(_0410_),
    .C(_0411_),
    .D(_0412_),
    .Y(_0063_));
 sg13g2_or2_1 _1007_ (.X(_0413_),
    .B(_0411_),
    .A(\cb[6] ));
 sg13g2_and2_1 _1008_ (.A(\cb[6] ),
    .B(_0411_),
    .X(_0414_));
 sg13g2_a22oi_1 _1009_ (.Y(_0415_),
    .B1(_0413_),
    .B2(net19),
    .A2(net16),
    .A1(\ca[14] ));
 sg13g2_nor3_1 _1010_ (.A(net52),
    .B(_0414_),
    .C(_0415_),
    .Y(_0064_));
 sg13g2_nand3b_1 _1011_ (.B(\cb[7] ),
    .C(net19),
    .Y(_0416_),
    .A_N(_0414_));
 sg13g2_a22oi_1 _1012_ (.Y(_0417_),
    .B1(_0414_),
    .B2(_0091_),
    .A2(net16),
    .A1(\ca[15] ));
 sg13g2_a21oi_1 _1013_ (.A1(_0416_),
    .A2(_0417_),
    .Y(_0065_),
    .B1(net51));
 sg13g2_nand4_1 _1014_ (.B(\cb[6] ),
    .C(\cb[5] ),
    .A(\cb[7] ),
    .Y(_0418_),
    .D(\cb[4] ));
 sg13g2_nor2_1 _1015_ (.A(_0404_),
    .B(_0418_),
    .Y(_0419_));
 sg13g2_and2_1 _1016_ (.A(\cb[8] ),
    .B(_0419_),
    .X(_0420_));
 sg13g2_a21oi_1 _1017_ (.A1(net55),
    .A2(_0420_),
    .Y(_0421_),
    .B1(net23));
 sg13g2_o21ai_1 _1018_ (.B1(_0421_),
    .Y(_0422_),
    .A1(\cb[8] ),
    .A2(_0419_));
 sg13g2_nand3_1 _1019_ (.B(_0121_),
    .C(net35),
    .A(\cb[0] ),
    .Y(_0423_));
 sg13g2_o21ai_1 _1020_ (.B1(net41),
    .Y(_0424_),
    .A1(\cb[8] ),
    .A2(net17));
 sg13g2_a21oi_1 _1021_ (.A1(_0422_),
    .A2(_0423_),
    .Y(_0066_),
    .B1(_0424_));
 sg13g2_and3_2 _1022_ (.X(_0425_),
    .A(\cb[9] ),
    .B(net55),
    .C(_0420_));
 sg13g2_o21ai_1 _1023_ (.B1(net19),
    .Y(_0426_),
    .A1(\cb[9] ),
    .A2(_0420_));
 sg13g2_nand3_1 _1024_ (.B(net49),
    .C(net35),
    .A(\cb[1] ),
    .Y(_0427_));
 sg13g2_o21ai_1 _1025_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0425_),
    .A2(_0426_));
 sg13g2_o21ai_1 _1026_ (.B1(_0428_),
    .Y(_0429_),
    .A1(\cb[9] ),
    .A2(net17));
 sg13g2_nor2_1 _1027_ (.A(net50),
    .B(_0429_),
    .Y(_0067_));
 sg13g2_a21oi_1 _1028_ (.A1(\cb[10] ),
    .A2(net19),
    .Y(_0430_),
    .B1(_0425_));
 sg13g2_a21oi_1 _1029_ (.A1(\cb[10] ),
    .A2(_0425_),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_a21oi_1 _1030_ (.A1(\cb[2] ),
    .A2(net16),
    .Y(_0432_),
    .B1(_0431_));
 sg13g2_nor2_1 _1031_ (.A(net50),
    .B(_0432_),
    .Y(_0068_));
 sg13g2_a22oi_1 _1032_ (.Y(_0433_),
    .B1(_0425_),
    .B2(\cb[10] ),
    .A2(net19),
    .A1(\cb[11] ));
 sg13g2_inv_1 _1033_ (.Y(_0434_),
    .A(_0433_));
 sg13g2_nand3_1 _1034_ (.B(\cb[10] ),
    .C(_0425_),
    .A(\cb[11] ),
    .Y(_0435_));
 sg13g2_and3_1 _1035_ (.X(_0436_),
    .A(\cb[11] ),
    .B(\cb[10] ),
    .C(\cb[9] ));
 sg13g2_a22oi_1 _1036_ (.Y(_0437_),
    .B1(_0434_),
    .B2(_0435_),
    .A2(net16),
    .A1(\cb[3] ));
 sg13g2_nor2_1 _1037_ (.A(net50),
    .B(_0437_),
    .Y(_0069_));
 sg13g2_o21ai_1 _1038_ (.B1(_0435_),
    .Y(_0438_),
    .A1(_0088_),
    .A2(net23));
 sg13g2_or2_1 _1039_ (.X(_0439_),
    .B(_0435_),
    .A(_0088_));
 sg13g2_a22oi_1 _1040_ (.Y(_0440_),
    .B1(_0438_),
    .B2(_0439_),
    .A2(net16),
    .A1(\cb[4] ));
 sg13g2_nor2_1 _1041_ (.A(net50),
    .B(_0440_),
    .Y(_0070_));
 sg13g2_nand3_1 _1042_ (.B(net22),
    .C(_0439_),
    .A(\cb[13] ),
    .Y(_0441_));
 sg13g2_nor2_1 _1043_ (.A(\cb[13] ),
    .B(_0439_),
    .Y(_0442_));
 sg13g2_a21oi_1 _1044_ (.A1(\cb[5] ),
    .A2(net16),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_a21oi_1 _1045_ (.A1(_0441_),
    .A2(_0443_),
    .Y(_0071_),
    .B1(net50));
 sg13g2_nand4_1 _1046_ (.B(\cb[12] ),
    .C(_0420_),
    .A(\cb[13] ),
    .Y(_0444_),
    .D(_0436_));
 sg13g2_a22oi_1 _1047_ (.Y(_0445_),
    .B1(_0214_),
    .B2(\cb[6] ),
    .A2(_0205_),
    .A1(\cb[14] ));
 sg13g2_nand2_1 _1048_ (.Y(_0446_),
    .A(_0086_),
    .B(_0444_));
 sg13g2_or2_1 _1049_ (.X(_0447_),
    .B(_0444_),
    .A(_0086_));
 sg13g2_nand3_1 _1050_ (.B(_0446_),
    .C(_0447_),
    .A(net58),
    .Y(_0448_));
 sg13g2_a21oi_1 _1051_ (.A1(_0445_),
    .A2(_0448_),
    .Y(_0072_),
    .B1(net53));
 sg13g2_xnor2_1 _1052_ (.Y(_0449_),
    .A(\cb[15] ),
    .B(_0447_));
 sg13g2_nand2_1 _1053_ (.Y(_0450_),
    .A(net58),
    .B(_0449_));
 sg13g2_a22oi_1 _1054_ (.Y(_0451_),
    .B1(net16),
    .B2(\cb[7] ),
    .A2(_0205_),
    .A1(\cb[15] ));
 sg13g2_a21oi_1 _1055_ (.A1(_0450_),
    .A2(_0451_),
    .Y(_0073_),
    .B1(net53));
 sg13g2_o21ai_1 _1056_ (.B1(net41),
    .Y(_0452_),
    .A1(\shift_counter[0] ),
    .A2(net29));
 sg13g2_a21oi_1 _1057_ (.A1(_0084_),
    .A2(net29),
    .Y(_0074_),
    .B1(_0452_));
 sg13g2_a21oi_1 _1058_ (.A1(\shift_counter[0] ),
    .A2(net29),
    .Y(_0453_),
    .B1(\shift_counter[1] ));
 sg13g2_o21ai_1 _1059_ (.B1(net41),
    .Y(_0454_),
    .A1(net24),
    .A2(net35));
 sg13g2_nor2_1 _1060_ (.A(_0453_),
    .B(_0454_),
    .Y(_0075_));
 sg13g2_and2_1 _1061_ (.A(net54),
    .B(net15),
    .X(_0076_));
 sg13g2_and2_1 _1062_ (.A(\stopedge.buff[0] ),
    .B(net53),
    .X(_0077_));
 sg13g2_and2_1 _1063_ (.A(\stopedge.buff[1] ),
    .B(net53),
    .X(_0078_));
 sg13g2_and2_1 _1064_ (.A(\stopedge.buff[2] ),
    .B(reset),
    .X(_0079_));
 sg13g2_and2_1 _1065_ (.A(net54),
    .B(net12),
    .X(_0080_));
 sg13g2_and2_1 _1066_ (.A(\shiftedge.buff[0] ),
    .B(net54),
    .X(_0081_));
 sg13g2_and2_1 _1067_ (.A(\shiftedge.buff[1] ),
    .B(net54),
    .X(_0082_));
 sg13g2_and2_1 _1068_ (.A(\shiftedge.buff[2] ),
    .B(net54),
    .X(_0083_));
 sg13g2_dfrbp_1 _1069_ (.CLK(net63),
    .RESET_B(net165),
    .D(_0004_),
    .Q_N(_0003_),
    .Q(\clock_div[0] ));
 sg13g2_dfrbp_1 _1070_ (.CLK(net63),
    .RESET_B(net92),
    .D(_0005_),
    .Q_N(_0530_),
    .Q(\clock_div[1] ));
 sg13g2_dfrbp_1 _1071_ (.CLK(net62),
    .RESET_B(net91),
    .D(_0006_),
    .Q_N(_0529_),
    .Q(\clock_div[2] ));
 sg13g2_dfrbp_1 _1072_ (.CLK(net62),
    .RESET_B(net90),
    .D(_0007_),
    .Q_N(_0528_),
    .Q(\clock_div[3] ));
 sg13g2_dfrbp_1 _1073_ (.CLK(net62),
    .RESET_B(net89),
    .D(_0008_),
    .Q_N(_0527_),
    .Q(done));
 sg13g2_dfrbp_1 _1074_ (.CLK(net64),
    .RESET_B(net169),
    .D(_0009_),
    .Q_N(_0526_),
    .Q(run));
 sg13g2_dfrbp_1 _1075_ (.CLK(net67),
    .RESET_B(net167),
    .D(_0010_),
    .Q_N(_0525_),
    .Q(\da[0] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(net67),
    .RESET_B(net163),
    .D(_0011_),
    .Q_N(_0524_),
    .Q(\da[1] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(net69),
    .RESET_B(net161),
    .D(_0012_),
    .Q_N(_0523_),
    .Q(\da[2] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(net69),
    .RESET_B(net159),
    .D(_0013_),
    .Q_N(_0522_),
    .Q(\da[3] ));
 sg13g2_dfrbp_1 _1079_ (.CLK(net68),
    .RESET_B(net157),
    .D(_0014_),
    .Q_N(_0521_),
    .Q(\da[4] ));
 sg13g2_dfrbp_1 _1080_ (.CLK(net71),
    .RESET_B(net155),
    .D(_0015_),
    .Q_N(_0520_),
    .Q(\da[5] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(net71),
    .RESET_B(net153),
    .D(_0016_),
    .Q_N(_0519_),
    .Q(\da[6] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(net70),
    .RESET_B(net151),
    .D(_0017_),
    .Q_N(_0518_),
    .Q(\da[7] ));
 sg13g2_dfrbp_1 _1083_ (.CLK(net67),
    .RESET_B(net149),
    .D(_0018_),
    .Q_N(_0517_),
    .Q(\da[8] ));
 sg13g2_dfrbp_1 _1084_ (.CLK(net67),
    .RESET_B(net147),
    .D(_0019_),
    .Q_N(_0516_),
    .Q(\da[9] ));
 sg13g2_dfrbp_1 _1085_ (.CLK(net68),
    .RESET_B(net145),
    .D(_0020_),
    .Q_N(_0515_),
    .Q(\da[10] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(net68),
    .RESET_B(net143),
    .D(_0021_),
    .Q_N(_0514_),
    .Q(\da[11] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(net71),
    .RESET_B(net141),
    .D(_0022_),
    .Q_N(_0513_),
    .Q(\da[12] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(net71),
    .RESET_B(net139),
    .D(_0023_),
    .Q_N(_0512_),
    .Q(\da[13] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(net70),
    .RESET_B(net137),
    .D(_0024_),
    .Q_N(_0511_),
    .Q(\da[14] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(net64),
    .RESET_B(net135),
    .D(_0025_),
    .Q_N(_0510_),
    .Q(\da[15] ));
 sg13g2_dfrbp_1 _1091_ (.CLK(net67),
    .RESET_B(net133),
    .D(_0026_),
    .Q_N(_0509_),
    .Q(\db[0] ));
 sg13g2_dfrbp_1 _1092_ (.CLK(net67),
    .RESET_B(net131),
    .D(_0027_),
    .Q_N(_0508_),
    .Q(\db[1] ));
 sg13g2_dfrbp_1 _1093_ (.CLK(net68),
    .RESET_B(net129),
    .D(_0028_),
    .Q_N(_0507_),
    .Q(\db[2] ));
 sg13g2_dfrbp_1 _1094_ (.CLK(net68),
    .RESET_B(net127),
    .D(_0029_),
    .Q_N(_0506_),
    .Q(\db[3] ));
 sg13g2_dfrbp_1 _1095_ (.CLK(net71),
    .RESET_B(net125),
    .D(_0030_),
    .Q_N(_0505_),
    .Q(\db[4] ));
 sg13g2_dfrbp_1 _1096_ (.CLK(net72),
    .RESET_B(net123),
    .D(_0031_),
    .Q_N(_0504_),
    .Q(\db[5] ));
 sg13g2_dfrbp_1 _1097_ (.CLK(net73),
    .RESET_B(net121),
    .D(_0032_),
    .Q_N(_0503_),
    .Q(\db[6] ));
 sg13g2_dfrbp_1 _1098_ (.CLK(net70),
    .RESET_B(net119),
    .D(_0033_),
    .Q_N(_0502_),
    .Q(\db[7] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(net69),
    .RESET_B(net117),
    .D(_0034_),
    .Q_N(_0501_),
    .Q(\db[8] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(net67),
    .RESET_B(net115),
    .D(_0035_),
    .Q_N(_0500_),
    .Q(\db[9] ));
 sg13g2_dfrbp_1 _1101_ (.CLK(net68),
    .RESET_B(net113),
    .D(_0036_),
    .Q_N(_0499_),
    .Q(\db[10] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(net68),
    .RESET_B(net111),
    .D(_0037_),
    .Q_N(_0498_),
    .Q(\db[11] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(net68),
    .RESET_B(net109),
    .D(_0038_),
    .Q_N(_0497_),
    .Q(\db[12] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(net72),
    .RESET_B(net107),
    .D(_0039_),
    .Q_N(_0496_),
    .Q(\db[13] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(net70),
    .RESET_B(net105),
    .D(_0040_),
    .Q_N(_0495_),
    .Q(\db[14] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(net70),
    .RESET_B(net103),
    .D(_0041_),
    .Q_N(_0494_),
    .Q(\db[15] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(net60),
    .RESET_B(net101),
    .D(_0042_),
    .Q_N(_0000_),
    .Q(\ca[0] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(net66),
    .RESET_B(net99),
    .D(_0043_),
    .Q_N(_0493_),
    .Q(\ca[1] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(net66),
    .RESET_B(net97),
    .D(_0044_),
    .Q_N(_0492_),
    .Q(\ca[2] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(net61),
    .RESET_B(net95),
    .D(_0045_),
    .Q_N(_0491_),
    .Q(\ca[3] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(net66),
    .RESET_B(net93),
    .D(_0046_),
    .Q_N(_0490_),
    .Q(\ca[4] ));
 sg13g2_dfrbp_1 _1112_ (.CLK(net64),
    .RESET_B(net168),
    .D(_0047_),
    .Q_N(_0489_),
    .Q(\ca[5] ));
 sg13g2_dfrbp_1 _1113_ (.CLK(net65),
    .RESET_B(net162),
    .D(_0048_),
    .Q_N(_0488_),
    .Q(\ca[6] ));
 sg13g2_dfrbp_1 _1114_ (.CLK(net64),
    .RESET_B(net158),
    .D(_0049_),
    .Q_N(_0487_),
    .Q(\ca[7] ));
 sg13g2_dfrbp_1 _1115_ (.CLK(net67),
    .RESET_B(net154),
    .D(_0050_),
    .Q_N(_0486_),
    .Q(\ca[8] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(net61),
    .RESET_B(net150),
    .D(_0051_),
    .Q_N(_0485_),
    .Q(\ca[9] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(net61),
    .RESET_B(net146),
    .D(_0052_),
    .Q_N(_0484_),
    .Q(\ca[10] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(net60),
    .RESET_B(net142),
    .D(_0053_),
    .Q_N(_0483_),
    .Q(\ca[11] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(net64),
    .RESET_B(net138),
    .D(_0054_),
    .Q_N(_0482_),
    .Q(\ca[12] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(net63),
    .RESET_B(net134),
    .D(_0055_),
    .Q_N(_0481_),
    .Q(\ca[13] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(net64),
    .RESET_B(net130),
    .D(_0056_),
    .Q_N(_0480_),
    .Q(\ca[14] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(net63),
    .RESET_B(net126),
    .D(_0057_),
    .Q_N(_0479_),
    .Q(\ca[15] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(net61),
    .RESET_B(net122),
    .D(_0058_),
    .Q_N(_0001_),
    .Q(\cb[0] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(net60),
    .RESET_B(net118),
    .D(_0059_),
    .Q_N(_0478_),
    .Q(\cb[1] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(net60),
    .RESET_B(net114),
    .D(_0060_),
    .Q_N(_0477_),
    .Q(\cb[2] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(net60),
    .RESET_B(net110),
    .D(_0061_),
    .Q_N(_0476_),
    .Q(\cb[3] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(net62),
    .RESET_B(net106),
    .D(_0062_),
    .Q_N(_0475_),
    .Q(\cb[4] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(net62),
    .RESET_B(net102),
    .D(_0063_),
    .Q_N(_0474_),
    .Q(\cb[5] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(net62),
    .RESET_B(net98),
    .D(_0064_),
    .Q_N(_0473_),
    .Q(\cb[6] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(net63),
    .RESET_B(net94),
    .D(_0065_),
    .Q_N(_0472_),
    .Q(\cb[7] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(net61),
    .RESET_B(net164),
    .D(_0066_),
    .Q_N(_0471_),
    .Q(\cb[8] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(net60),
    .RESET_B(net156),
    .D(_0067_),
    .Q_N(_0470_),
    .Q(\cb[9] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(net61),
    .RESET_B(net148),
    .D(_0068_),
    .Q_N(_0469_),
    .Q(\cb[10] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(net61),
    .RESET_B(net140),
    .D(_0069_),
    .Q_N(_0468_),
    .Q(\cb[11] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(net62),
    .RESET_B(net132),
    .D(_0070_),
    .Q_N(_0467_),
    .Q(\cb[12] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(net62),
    .RESET_B(net124),
    .D(_0071_),
    .Q_N(_0466_),
    .Q(\cb[13] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(net70),
    .RESET_B(net116),
    .D(_0072_),
    .Q_N(_0465_),
    .Q(\cb[14] ));
 sg13g2_dfrbp_1 _1138_ (.CLK(net70),
    .RESET_B(net108),
    .D(_0073_),
    .Q_N(_0464_),
    .Q(\cb[15] ));
 sg13g2_dfrbp_1 _1139_ (.CLK(net60),
    .RESET_B(net100),
    .D(_0074_),
    .Q_N(_0002_),
    .Q(\shift_counter[0] ));
 sg13g2_dfrbp_1 _1140_ (.CLK(net60),
    .RESET_B(net170),
    .D(_0075_),
    .Q_N(_0463_),
    .Q(\shift_counter[1] ));
 sg13g2_dfrbp_1 _1141_ (.CLK(net70),
    .RESET_B(net152),
    .D(_0076_),
    .Q_N(_0462_),
    .Q(\stopedge.buff[0] ));
 sg13g2_dfrbp_1 _1142_ (.CLK(net64),
    .RESET_B(net144),
    .D(_0077_),
    .Q_N(_0461_),
    .Q(\stopedge.buff[1] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(net64),
    .RESET_B(net136),
    .D(_0078_),
    .Q_N(_0460_),
    .Q(\stopedge.buff[2] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(net73),
    .RESET_B(net166),
    .D(_0079_),
    .Q_N(_0531_),
    .Q(\stopedge.buff[3] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(net71),
    .RESET_B(net160),
    .D(\resetsync.in ),
    .Q_N(_0532_),
    .Q(\resetsync.buff[0] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(net71),
    .RESET_B(net128),
    .D(\resetsync.buff[0] ),
    .Q_N(_0459_),
    .Q(reset));
 sg13g2_dfrbp_1 _1147_ (.CLK(net72),
    .RESET_B(net120),
    .D(_0080_),
    .Q_N(_0458_),
    .Q(\shiftedge.buff[0] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(net72),
    .RESET_B(net112),
    .D(_0081_),
    .Q_N(_0457_),
    .Q(\shiftedge.buff[1] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(net72),
    .RESET_B(net104),
    .D(_0082_),
    .Q_N(_0456_),
    .Q(\shiftedge.buff[2] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(net71),
    .RESET_B(net96),
    .D(_0083_),
    .Q_N(_0455_),
    .Q(\shiftedge.buff[3] ));
 sg13g2_tiehi _1072__90 (.L_HI(net90));
 sg13g2_tiehi _1071__91 (.L_HI(net91));
 sg13g2_tiehi _1070__92 (.L_HI(net92));
 sg13g2_tiehi _1111__93 (.L_HI(net93));
 sg13g2_tiehi _1130__94 (.L_HI(net94));
 sg13g2_tiehi _1110__95 (.L_HI(net95));
 sg13g2_tiehi _1150__96 (.L_HI(net96));
 sg13g2_tiehi _1109__97 (.L_HI(net97));
 sg13g2_tiehi _1129__98 (.L_HI(net98));
 sg13g2_tiehi _1108__99 (.L_HI(net99));
 sg13g2_tiehi _1139__100 (.L_HI(net100));
 sg13g2_tiehi _1107__101 (.L_HI(net101));
 sg13g2_tiehi _1128__102 (.L_HI(net102));
 sg13g2_tiehi _1106__103 (.L_HI(net103));
 sg13g2_tiehi _1149__104 (.L_HI(net104));
 sg13g2_tiehi _1105__105 (.L_HI(net105));
 sg13g2_tiehi _1127__106 (.L_HI(net106));
 sg13g2_tiehi _1104__107 (.L_HI(net107));
 sg13g2_tiehi _1138__108 (.L_HI(net108));
 sg13g2_tiehi _1103__109 (.L_HI(net109));
 sg13g2_tiehi _1126__110 (.L_HI(net110));
 sg13g2_tiehi _1102__111 (.L_HI(net111));
 sg13g2_tiehi _1148__112 (.L_HI(net112));
 sg13g2_tiehi _1101__113 (.L_HI(net113));
 sg13g2_tiehi _1125__114 (.L_HI(net114));
 sg13g2_tiehi _1100__115 (.L_HI(net115));
 sg13g2_tiehi _1137__116 (.L_HI(net116));
 sg13g2_tiehi _1099__117 (.L_HI(net117));
 sg13g2_tiehi _1124__118 (.L_HI(net118));
 sg13g2_tiehi _1098__119 (.L_HI(net119));
 sg13g2_tiehi _1147__120 (.L_HI(net120));
 sg13g2_tiehi _1097__121 (.L_HI(net121));
 sg13g2_tiehi _1123__122 (.L_HI(net122));
 sg13g2_tiehi _1096__123 (.L_HI(net123));
 sg13g2_tiehi _1136__124 (.L_HI(net124));
 sg13g2_tiehi _1095__125 (.L_HI(net125));
 sg13g2_tiehi _1122__126 (.L_HI(net126));
 sg13g2_tiehi _1094__127 (.L_HI(net127));
 sg13g2_tiehi _1146__128 (.L_HI(net128));
 sg13g2_tiehi _1093__129 (.L_HI(net129));
 sg13g2_tiehi _1121__130 (.L_HI(net130));
 sg13g2_tiehi _1092__131 (.L_HI(net131));
 sg13g2_tiehi _1135__132 (.L_HI(net132));
 sg13g2_tiehi _1091__133 (.L_HI(net133));
 sg13g2_tiehi _1120__134 (.L_HI(net134));
 sg13g2_tiehi _1090__135 (.L_HI(net135));
 sg13g2_tiehi _1143__136 (.L_HI(net136));
 sg13g2_tiehi _1089__137 (.L_HI(net137));
 sg13g2_tiehi _1119__138 (.L_HI(net138));
 sg13g2_tiehi _1088__139 (.L_HI(net139));
 sg13g2_tiehi _1134__140 (.L_HI(net140));
 sg13g2_tiehi _1087__141 (.L_HI(net141));
 sg13g2_tiehi _1118__142 (.L_HI(net142));
 sg13g2_tiehi _1086__143 (.L_HI(net143));
 sg13g2_tiehi _1142__144 (.L_HI(net144));
 sg13g2_tiehi _1085__145 (.L_HI(net145));
 sg13g2_tiehi _1117__146 (.L_HI(net146));
 sg13g2_tiehi _1084__147 (.L_HI(net147));
 sg13g2_tiehi _1133__148 (.L_HI(net148));
 sg13g2_tiehi _1083__149 (.L_HI(net149));
 sg13g2_tiehi _1116__150 (.L_HI(net150));
 sg13g2_tiehi _1082__151 (.L_HI(net151));
 sg13g2_tiehi _1141__152 (.L_HI(net152));
 sg13g2_tiehi _1081__153 (.L_HI(net153));
 sg13g2_tiehi _1115__154 (.L_HI(net154));
 sg13g2_tiehi _1080__155 (.L_HI(net155));
 sg13g2_tiehi _1132__156 (.L_HI(net156));
 sg13g2_tiehi _1079__157 (.L_HI(net157));
 sg13g2_tiehi _1114__158 (.L_HI(net158));
 sg13g2_tiehi _1078__159 (.L_HI(net159));
 sg13g2_tiehi _1145__160 (.L_HI(net160));
 sg13g2_tiehi _1077__161 (.L_HI(net161));
 sg13g2_tiehi _1113__162 (.L_HI(net162));
 sg13g2_tiehi _1076__163 (.L_HI(net163));
 sg13g2_tiehi _1131__164 (.L_HI(net164));
 sg13g2_tiehi _1069__165 (.L_HI(net165));
 sg13g2_tiehi _1144__166 (.L_HI(net166));
 sg13g2_tiehi _1075__167 (.L_HI(net167));
 sg13g2_tiehi _1112__168 (.L_HI(net168));
 sg13g2_tiehi _1074__169 (.L_HI(net169));
 sg13g2_tiehi _1140__170 (.L_HI(net170));
 sg13g2_tiehi tt_um_algofoogle_ro_worker_171 (.L_HI(net171));
 sg13g2_tiehi tt_um_algofoogle_ro_worker_172 (.L_HI(net172));
 sg13g2_tiehi tt_um_algofoogle_ro_worker_173 (.L_HI(net173));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo tt_um_algofoogle_ro_worker_80 (.L_LO(net80));
 sg13g2_tielo tt_um_algofoogle_ro_worker_81 (.L_LO(net81));
 sg13g2_tielo tt_um_algofoogle_ro_worker_82 (.L_LO(net82));
 sg13g2_tielo tt_um_algofoogle_ro_worker_83 (.L_LO(net83));
 sg13g2_tielo tt_um_algofoogle_ro_worker_84 (.L_LO(net84));
 sg13g2_tielo tt_um_algofoogle_ro_worker_85 (.L_LO(net85));
 sg13g2_tielo tt_um_algofoogle_ro_worker_86 (.L_LO(net86));
 sg13g2_tielo tt_um_algofoogle_ro_worker_87 (.L_LO(net87));
 sg13g2_tielo tt_um_algofoogle_ro_worker_88 (.L_LO(net88));
 sg13g2_tiehi _1073__89 (.L_HI(net89));
 sg13g2_buf_1 _1246_ (.A(net57),
    .X(uio_out[5]));
 sg13g2_buf_1 _1247_ (.A(done),
    .X(uio_out[6]));
 sg13g2_buf_1 _1248_ (.A(\clock_div[3] ),
    .X(uio_out[7]));
 sg13g2_buf_1 _1249_ (.A(\ca[8] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1250_ (.A(\ca[9] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1251_ (.A(\ca[10] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _1252_ (.A(\ca[11] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1253_ (.A(\ca[12] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _1254_ (.A(\ca[13] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _1255_ (.A(\ca[14] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _1256_ (.A(\ca[15] ),
    .X(uo_out[7]));
 sg13g2_buf_8 intclkbuff (.A(internal_clock_unbuffered),
    .X(internal_clock));
 sg13g2_inv_1 \myring.inv_array[0]/inverter  (.Y(\myring.inv_in[1] ),
    .A(\myring.inv_in[0] ));
 sg13g2_inv_1 \myring.inv_array[1]/inverter  (.Y(\myring.inv_in[2] ),
    .A(\myring.inv_in[1] ));
 sg13g2_inv_1 \myring.inv_array[2]/inverter  (.Y(\myring.inv_in[3] ),
    .A(\myring.inv_in[2] ));
 sg13g2_inv_1 \myring.inv_array[3]/inverter  (.Y(\myring.inv_in[4] ),
    .A(\myring.inv_in[3] ));
 sg13g2_inv_1 \myring.inv_array[4]/inverter  (.Y(\myring.inv_in[5] ),
    .A(\myring.inv_in[4] ));
 sg13g2_inv_1 \myring.inv_array[5]/inverter  (.Y(\myring.inv_in[6] ),
    .A(\myring.inv_in[5] ));
 sg13g2_inv_1 \myring.inv_array[6]/inverter  (.Y(\myring.inv_in[7] ),
    .A(\myring.inv_in[6] ));
 sg13g2_inv_1 \myring.inv_array[7]/inverter  (.Y(\myring.inv_in[8] ),
    .A(\myring.inv_in[7] ));
 sg13g2_inv_1 \myring.inv_array[8]/inverter  (.Y(\myring.inv_out[8] ),
    .A(\myring.inv_in[8] ));
 sg13g2_buf_1 input1 (.A(clk),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ena),
    .X(net2));
 sg13g2_buf_1 input3 (.A(rst_n),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[0]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[1]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[2]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[3]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[4]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[5]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(ui_in[6]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(ui_in[7]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[0]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[1]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[2]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[3]),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0214_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0206_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0206_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(net22),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(net22),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(net22),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0202_),
    .X(net22));
 sg13g2_buf_4 fanout23 (.X(net23),
    .A(_0201_));
 sg13g2_buf_4 fanout24 (.X(net24),
    .A(_0162_));
 sg13g2_buf_2 fanout25 (.A(net28),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(net27),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(net28),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0162_),
    .X(net28));
 sg13g2_buf_4 fanout29 (.X(net29),
    .A(_0161_));
 sg13g2_buf_2 fanout30 (.A(_0161_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(net34),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(net34),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0161_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(net37),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(net37),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0165_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_0164_));
 sg13g2_buf_2 fanout39 (.A(_0164_),
    .X(net39));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(_0164_));
 sg13g2_buf_2 fanout41 (.A(net43),
    .X(net41));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net43));
 sg13g2_buf_2 fanout43 (.A(net48),
    .X(net43));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(net48));
 sg13g2_buf_1 fanout45 (.A(net48),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0123_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0121_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(net52),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(net52),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(net53),
    .X(net52));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(net54));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(reset));
 sg13g2_buf_2 fanout55 (.A(net59),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(net59),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(net59),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(net59),
    .X(net58));
 sg13g2_buf_1 fanout59 (.A(run),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(net61),
    .X(net60));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net66));
 sg13g2_buf_2 fanout62 (.A(net65),
    .X(net62));
 sg13g2_buf_1 fanout63 (.A(net65),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(net65),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(internal_clock),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(net69),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(net69),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(internal_clock),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(net73),
    .X(net70));
 sg13g2_buf_4 fanout71 (.X(net71),
    .A(net73));
 sg13g2_buf_2 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(internal_clock),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(net75),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net14),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(net14),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(net14),
    .X(net78));
 sg13g2_tielo tt_um_algofoogle_ro_worker_79 (.L_LO(net79));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_4 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_decap_4 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_4 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_4 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_fill_2 FILLER_15_160 ();
 sg13g2_fill_1 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_decap_4 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_120 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_4 FILLER_16_132 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_decap_8 FILLER_16_178 ();
 sg13g2_decap_4 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_201 ();
 sg13g2_decap_4 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_4 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_246 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_260 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_4 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_4 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_fill_2 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_decap_4 FILLER_17_171 ();
 sg13g2_decap_8 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_228 ();
 sg13g2_decap_4 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_decap_8 FILLER_17_267 ();
 sg13g2_fill_2 FILLER_17_274 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_317 ();
 sg13g2_decap_4 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_decap_4 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_315 ();
 sg13g2_decap_4 FILLER_18_329 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_4 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_fill_2 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_101 ();
 sg13g2_decap_8 FILLER_19_107 ();
 sg13g2_fill_2 FILLER_19_114 ();
 sg13g2_decap_4 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_205 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_238 ();
 sg13g2_fill_2 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_decap_4 FILLER_19_290 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_4 FILLER_19_389 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_decap_4 FILLER_20_122 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_decap_4 FILLER_20_152 ();
 sg13g2_decap_4 FILLER_20_167 ();
 sg13g2_decap_8 FILLER_20_177 ();
 sg13g2_decap_4 FILLER_20_184 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_2 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_4 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_decap_4 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_decap_4 FILLER_20_356 ();
 sg13g2_fill_2 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_fill_1 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_90 ();
 sg13g2_decap_8 FILLER_21_97 ();
 sg13g2_decap_4 FILLER_21_104 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_decap_4 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_decap_8 FILLER_21_288 ();
 sg13g2_decap_4 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_decap_4 FILLER_21_342 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_decap_4 FILLER_21_378 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_2 FILLER_22_72 ();
 sg13g2_fill_1 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_79 ();
 sg13g2_decap_4 FILLER_22_86 ();
 sg13g2_decap_4 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_fill_2 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_decap_4 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_172 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_237 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_4 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_353 ();
 sg13g2_decap_4 FILLER_22_360 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_fill_2 FILLER_22_375 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_decap_4 FILLER_22_388 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_46 ();
 sg13g2_decap_4 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_106 ();
 sg13g2_decap_8 FILLER_23_113 ();
 sg13g2_decap_4 FILLER_23_120 ();
 sg13g2_decap_4 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_156 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_decap_4 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_decap_4 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_265 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_fill_1 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_decap_4 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_decap_4 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_4 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_60 ();
 sg13g2_fill_2 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_fill_2 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_fill_2 FILLER_24_149 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_191 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_decap_8 FILLER_24_215 ();
 sg13g2_decap_4 FILLER_24_222 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_decap_4 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_fill_2 FILLER_24_267 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_decap_4 FILLER_24_327 ();
 sg13g2_fill_2 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_fill_1 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_decap_4 FILLER_24_384 ();
 sg13g2_fill_1 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_96 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_decap_8 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_4 FILLER_25_163 ();
 sg13g2_decap_4 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_245 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_decap_4 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_decap_4 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_85 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_decap_4 FILLER_26_103 ();
 sg13g2_decap_4 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_136 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_decap_4 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_8 FILLER_26_230 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_4 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_decap_4 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_312 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_4 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_71 ();
 sg13g2_fill_2 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_103 ();
 sg13g2_decap_8 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_decap_4 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_216 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_4 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_4 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_299 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_4 FILLER_27_337 ();
 sg13g2_fill_2 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_374 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_fill_2 FILLER_28_82 ();
 sg13g2_decap_4 FILLER_28_94 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_decap_4 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_232 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_decap_4 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_301 ();
 sg13g2_decap_4 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_71 ();
 sg13g2_fill_2 FILLER_29_78 ();
 sg13g2_fill_2 FILLER_29_106 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_121 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_decap_4 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_4 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_184 ();
 sg13g2_fill_2 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_197 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_289 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_321 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_decap_4 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_4 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_fill_2 FILLER_30_89 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_109 ();
 sg13g2_decap_8 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_decap_4 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_208 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_decap_4 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_254 ();
 sg13g2_decap_8 FILLER_30_284 ();
 sg13g2_decap_4 FILLER_30_291 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_319 ();
 sg13g2_decap_4 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_decap_4 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_94 ();
 sg13g2_decap_8 FILLER_31_101 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_110 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_decap_4 FILLER_31_163 ();
 sg13g2_decap_4 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_decap_8 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_decap_4 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_270 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_fill_2 FILLER_31_292 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_decap_8 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_fill_2 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_decap_4 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_decap_4 FILLER_32_90 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_decap_4 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_decap_4 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_157 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_decap_4 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_decap_4 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_decap_4 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_255 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_decap_4 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_321 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_decap_4 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_4 FILLER_32_386 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_39 ();
 sg13g2_decap_8 FILLER_33_71 ();
 sg13g2_decap_4 FILLER_33_78 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_fill_2 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_decap_8 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_124 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_174 ();
 sg13g2_decap_4 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_decap_4 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_fill_1 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_55 ();
 sg13g2_fill_2 FILLER_34_96 ();
 sg13g2_fill_1 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_4 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_decap_4 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_decap_8 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_decap_4 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_280 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_290 ();
 sg13g2_decap_8 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_decap_4 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_85 ();
 sg13g2_decap_8 FILLER_35_92 ();
 sg13g2_decap_8 FILLER_35_99 ();
 sg13g2_decap_4 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_decap_8 FILLER_35_116 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_decap_4 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_209 ();
 sg13g2_fill_2 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_decap_4 FILLER_35_310 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_4 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_4 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_decap_8 FILLER_36_120 ();
 sg13g2_decap_4 FILLER_36_127 ();
 sg13g2_decap_8 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_4 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_decap_4 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_decap_4 FILLER_36_386 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_decap_8 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_decap_8 FILLER_37_101 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_fill_1 FILLER_37_166 ();
 sg13g2_fill_1 FILLER_37_315 ();
 sg13g2_decap_4 FILLER_37_345 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_162 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net79;
 assign uio_oe[1] = net80;
 assign uio_oe[2] = net81;
 assign uio_oe[3] = net82;
 assign uio_oe[4] = net83;
 assign uio_oe[5] = net171;
 assign uio_oe[6] = net172;
 assign uio_oe[7] = net173;
 assign uio_out[0] = net84;
 assign uio_out[1] = net85;
 assign uio_out[2] = net86;
 assign uio_out[3] = net87;
 assign uio_out[4] = net88;
endmodule
