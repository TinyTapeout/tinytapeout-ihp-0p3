module tt_um_zerotoasic_logo_screensaver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire clknet_0_clk;
 wire \color_index[0] ;
 wire \color_index[1] ;
 wire \color_index[2] ;
 wire dir_x;
 wire dir_y;
 wire \gamepad.decoder.data_reg[0] ;
 wire \gamepad.decoder.data_reg[10] ;
 wire \gamepad.decoder.data_reg[11] ;
 wire \gamepad.decoder.data_reg[1] ;
 wire \gamepad.decoder.data_reg[2] ;
 wire \gamepad.decoder.data_reg[3] ;
 wire \gamepad.decoder.data_reg[4] ;
 wire \gamepad.decoder.data_reg[5] ;
 wire \gamepad.decoder.data_reg[6] ;
 wire \gamepad.decoder.data_reg[7] ;
 wire \gamepad.decoder.data_reg[8] ;
 wire \gamepad.decoder.data_reg[9] ;
 wire \gamepad.driver.pmod_clk_prev ;
 wire \gamepad.driver.pmod_clk_sync[0] ;
 wire \gamepad.driver.pmod_clk_sync[1] ;
 wire \gamepad.driver.pmod_data_sync[0] ;
 wire \gamepad.driver.pmod_data_sync[1] ;
 wire \gamepad.driver.pmod_latch_prev ;
 wire \gamepad.driver.pmod_latch_sync[0] ;
 wire \gamepad.driver.pmod_latch_sync[1] ;
 wire \gamepad.driver.shift_reg[0] ;
 wire \gamepad.driver.shift_reg[10] ;
 wire \gamepad.driver.shift_reg[11] ;
 wire \gamepad.driver.shift_reg[1] ;
 wire \gamepad.driver.shift_reg[2] ;
 wire \gamepad.driver.shift_reg[3] ;
 wire \gamepad.driver.shift_reg[4] ;
 wire \gamepad.driver.shift_reg[5] ;
 wire \gamepad.driver.shift_reg[6] ;
 wire \gamepad.driver.shift_reg[7] ;
 wire \gamepad.driver.shift_reg[8] ;
 wire \gamepad.driver.shift_reg[9] ;
 wire gamepad_start_prev;
 wire hsync;
 wire \logo_left[0] ;
 wire \logo_left[1] ;
 wire \logo_left[2] ;
 wire \logo_left[3] ;
 wire \logo_left[4] ;
 wire \logo_left[5] ;
 wire \logo_left[6] ;
 wire \logo_left[7] ;
 wire \logo_left[8] ;
 wire \logo_left[9] ;
 wire \logo_top[0] ;
 wire \logo_top[1] ;
 wire \logo_top[2] ;
 wire \logo_top[3] ;
 wire \logo_top[4] ;
 wire \logo_top[5] ;
 wire \logo_top[6] ;
 wire \logo_top[7] ;
 wire \logo_top[8] ;
 wire \logo_top[9] ;
 wire manual_mode;
 wire \palette_inst.rrggbb[0] ;
 wire \palette_inst.rrggbb[1] ;
 wire \palette_inst.rrggbb[2] ;
 wire \palette_inst.rrggbb[3] ;
 wire \palette_inst.rrggbb[4] ;
 wire \palette_inst.rrggbb[5] ;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \prev_y[0] ;
 wire \prev_y[1] ;
 wire \prev_y[2] ;
 wire \prev_y[3] ;
 wire \prev_y[4] ;
 wire \prev_y[5] ;
 wire \prev_y[6] ;
 wire \prev_y[7] ;
 wire \prev_y[8] ;
 wire \prev_y[9] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire \vga_sync_gen.vsync ;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;

 sg13g2_inv_1 _1708_ (.Y(_0744_),
    .A(net186));
 sg13g2_inv_1 _1709_ (.Y(_0745_),
    .A(net196));
 sg13g2_inv_1 _1710_ (.Y(_0746_),
    .A(net204));
 sg13g2_inv_1 _1711_ (.Y(_0747_),
    .A(net207));
 sg13g2_inv_1 _1712_ (.Y(_0748_),
    .A(net192));
 sg13g2_inv_1 _1713_ (.Y(_0749_),
    .A(net188));
 sg13g2_inv_1 _1714_ (.Y(_0750_),
    .A(net214));
 sg13g2_inv_1 _1715_ (.Y(_0751_),
    .A(net180));
 sg13g2_inv_1 _1716_ (.Y(_0752_),
    .A(net200));
 sg13g2_inv_1 _1717_ (.Y(_0753_),
    .A(net206));
 sg13g2_inv_1 _1718_ (.Y(_0754_),
    .A(net202));
 sg13g2_inv_1 _1719_ (.Y(_0755_),
    .A(\gamepad.driver.pmod_data_sync[1] ));
 sg13g2_inv_1 _1720_ (.Y(_0756_),
    .A(net784));
 sg13g2_inv_2 _1721_ (.Y(_0757_),
    .A(net789));
 sg13g2_inv_2 _1722_ (.Y(_0758_),
    .A(net268));
 sg13g2_inv_1 _1723_ (.Y(_0759_),
    .A(\logo_top[8] ));
 sg13g2_inv_1 _1724_ (.Y(_0760_),
    .A(net269));
 sg13g2_inv_1 _1725_ (.Y(_0761_),
    .A(\logo_top[3] ));
 sg13g2_inv_1 _1726_ (.Y(_0762_),
    .A(net242));
 sg13g2_inv_1 _1727_ (.Y(_0763_),
    .A(net138));
 sg13g2_inv_1 _1728_ (.Y(_0764_),
    .A(net798));
 sg13g2_inv_1 _1729_ (.Y(_0765_),
    .A(\logo_left[4] ));
 sg13g2_inv_1 _1730_ (.Y(_0766_),
    .A(net133));
 sg13g2_inv_1 _1731_ (.Y(_0767_),
    .A(net178));
 sg13g2_inv_1 _1732_ (.Y(_0768_),
    .A(\pix_y[0] ));
 sg13g2_inv_1 _1733_ (.Y(_0769_),
    .A(\pix_y[1] ));
 sg13g2_inv_2 _1734_ (.Y(_0770_),
    .A(\pix_y[2] ));
 sg13g2_inv_2 _1735_ (.Y(_0771_),
    .A(\pix_y[5] ));
 sg13g2_inv_2 _1736_ (.Y(_0772_),
    .A(net260));
 sg13g2_inv_2 _1737_ (.Y(_0773_),
    .A(net810));
 sg13g2_inv_2 _1738_ (.Y(_0774_),
    .A(net261));
 sg13g2_inv_2 _1739_ (.Y(_0775_),
    .A(net231));
 sg13g2_inv_1 _1740_ (.Y(_0776_),
    .A(\prev_y[0] ));
 sg13g2_inv_1 _1741_ (.Y(_0777_),
    .A(\prev_y[6] ));
 sg13g2_inv_1 _1742_ (.Y(_0778_),
    .A(\prev_y[8] ));
 sg13g2_inv_1 _1743_ (.Y(_0779_),
    .A(net159));
 sg13g2_inv_1 _1744_ (.Y(_0780_),
    .A(net150));
 sg13g2_inv_1 _1745_ (.Y(_0781_),
    .A(net142));
 sg13g2_inv_1 _1746_ (.Y(_0782_),
    .A(net140));
 sg13g2_inv_1 _1747_ (.Y(_0783_),
    .A(net148));
 sg13g2_inv_1 _1748_ (.Y(_0784_),
    .A(net210));
 sg13g2_inv_1 _1749_ (.Y(_0785_),
    .A(net198));
 sg13g2_inv_1 _1750_ (.Y(_0786_),
    .A(net194));
 sg13g2_inv_1 _1751_ (.Y(_0787_),
    .A(net209));
 sg13g2_inv_1 _1752_ (.Y(_0788_),
    .A(net161));
 sg13g2_inv_1 _1753_ (.Y(_0789_),
    .A(net182));
 sg13g2_inv_1 _1754_ (.Y(_0790_),
    .A(net144));
 sg13g2_inv_1 _1755_ (.Y(_0791_),
    .A(net154));
 sg13g2_inv_1 _1756_ (.Y(_0792_),
    .A(_0010_));
 sg13g2_inv_1 _1757_ (.Y(_0793_),
    .A(_0014_));
 sg13g2_inv_1 _1758_ (.Y(_0794_),
    .A(net127));
 sg13g2_nand2_1 _1759_ (.Y(_0795_),
    .A(\pix_y[5] ),
    .B(\pix_y[6] ));
 sg13g2_nand3_1 _1760_ (.B(\pix_y[6] ),
    .C(net231),
    .A(\pix_y[5] ),
    .Y(_0796_));
 sg13g2_or2_1 _1761_ (.X(_0797_),
    .B(_0796_),
    .A(_0774_));
 sg13g2_inv_1 _1762_ (.Y(_0798_),
    .A(_0797_));
 sg13g2_nor2_1 _1763_ (.A(net230),
    .B(_0797_),
    .Y(_0799_));
 sg13g2_nor3_1 _1764_ (.A(_0769_),
    .B(\pix_y[2] ),
    .C(\pix_y[4] ),
    .Y(_0800_));
 sg13g2_and3_1 _1765_ (.X(_0006_),
    .A(net783),
    .B(_0799_),
    .C(_0800_));
 sg13g2_and2_1 _1766_ (.A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .X(_0801_));
 sg13g2_and2_1 _1767_ (.A(net217),
    .B(_0801_),
    .X(_0802_));
 sg13g2_nor3_1 _1768_ (.A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .C(net217),
    .Y(_0803_));
 sg13g2_nand2_1 _1769_ (.Y(_0804_),
    .A(\pix_x[7] ),
    .B(net224));
 sg13g2_nor4_1 _1770_ (.A(\pix_x[8] ),
    .B(_0802_),
    .C(_0803_),
    .D(net225),
    .Y(_0005_));
 sg13g2_xor2_1 _1771_ (.B(\prev_y[7] ),
    .A(\pix_y[7] ),
    .X(_0805_));
 sg13g2_xnor2_1 _1772_ (.Y(_0806_),
    .A(\pix_y[9] ),
    .B(\prev_y[9] ));
 sg13g2_nor2_1 _1773_ (.A(_0771_),
    .B(\prev_y[5] ),
    .Y(_0807_));
 sg13g2_nor2_1 _1774_ (.A(_0769_),
    .B(\prev_y[1] ),
    .Y(_0808_));
 sg13g2_nand2_1 _1775_ (.Y(_0809_),
    .A(_0772_),
    .B(\prev_y[6] ));
 sg13g2_xnor2_1 _1776_ (.Y(_0810_),
    .A(\pix_y[4] ),
    .B(\prev_y[4] ));
 sg13g2_a22oi_1 _1777_ (.Y(_0811_),
    .B1(\prev_y[2] ),
    .B2(_0770_),
    .A2(\prev_y[0] ),
    .A1(_0768_));
 sg13g2_a22oi_1 _1778_ (.Y(_0812_),
    .B1(\prev_y[8] ),
    .B2(_0774_),
    .A2(\prev_y[5] ),
    .A1(_0771_));
 sg13g2_xnor2_1 _1779_ (.Y(_0813_),
    .A(net783),
    .B(\prev_y[3] ));
 sg13g2_o21ai_1 _1780_ (.B1(_0809_),
    .Y(_0814_),
    .A1(_0770_),
    .A2(\prev_y[2] ));
 sg13g2_a221oi_1 _1781_ (.B2(\pix_y[8] ),
    .C1(_0805_),
    .B1(_0778_),
    .A1(\pix_y[6] ),
    .Y(_0815_),
    .A2(_0777_));
 sg13g2_a22oi_1 _1782_ (.Y(_0816_),
    .B1(\prev_y[1] ),
    .B2(_0769_),
    .A2(_0776_),
    .A1(\pix_y[0] ));
 sg13g2_nand4_1 _1783_ (.B(_0812_),
    .C(_0813_),
    .A(_0810_),
    .Y(_0817_),
    .D(_0816_));
 sg13g2_nor4_1 _1784_ (.A(_0807_),
    .B(_0808_),
    .C(_0814_),
    .D(_0817_),
    .Y(_0818_));
 sg13g2_nand4_1 _1785_ (.B(_0811_),
    .C(_0815_),
    .A(_0806_),
    .Y(_0819_),
    .D(_0818_));
 sg13g2_nor4_1 _1786_ (.A(\pix_y[0] ),
    .B(\pix_y[1] ),
    .C(\pix_y[4] ),
    .D(\pix_y[5] ),
    .Y(_0820_));
 sg13g2_nand4_1 _1787_ (.B(_0774_),
    .C(_0775_),
    .A(_0772_),
    .Y(_0821_),
    .D(_0820_));
 sg13g2_nor4_1 _1788_ (.A(\pix_y[2] ),
    .B(net782),
    .C(\pix_y[9] ),
    .D(_0821_),
    .Y(_0822_));
 sg13g2_and2_2 _1789_ (.A(_0819_),
    .B(_0822_),
    .X(_0823_));
 sg13g2_inv_1 _1790_ (.Y(_0824_),
    .A(_0823_));
 sg13g2_nand2_1 _1791_ (.Y(_0825_),
    .A(net780),
    .B(_0823_));
 sg13g2_nand2_2 _1792_ (.Y(_0826_),
    .A(\logo_top[1] ),
    .B(\logo_top[0] ));
 sg13g2_nand3_1 _1793_ (.B(net795),
    .C(\logo_top[0] ),
    .A(\logo_top[2] ),
    .Y(_0827_));
 sg13g2_nor2_1 _1794_ (.A(_0761_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_nand3_1 _1795_ (.B(\logo_top[4] ),
    .C(_0828_),
    .A(\logo_top[5] ),
    .Y(_0829_));
 sg13g2_inv_1 _1796_ (.Y(_0830_),
    .A(_0829_));
 sg13g2_nor2_1 _1797_ (.A(_0013_),
    .B(_0829_),
    .Y(_0831_));
 sg13g2_xor2_1 _1798_ (.B(_0829_),
    .A(_0013_),
    .X(_0832_));
 sg13g2_inv_1 _1799_ (.Y(_0833_),
    .A(_0832_));
 sg13g2_xnor2_1 _1800_ (.Y(_0834_),
    .A(\logo_top[7] ),
    .B(_0831_));
 sg13g2_inv_1 _1801_ (.Y(_0835_),
    .A(_0834_));
 sg13g2_and3_1 _1802_ (.X(_0836_),
    .A(\logo_top[7] ),
    .B(\logo_top[6] ),
    .C(_0830_));
 sg13g2_and2_1 _1803_ (.A(_0793_),
    .B(_0836_),
    .X(_0837_));
 sg13g2_nor3_1 _1804_ (.A(\logo_top[9] ),
    .B(_0793_),
    .C(_0836_),
    .Y(_0838_));
 sg13g2_a21oi_1 _1805_ (.A1(net793),
    .A2(_0837_),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nor2_1 _1806_ (.A(net795),
    .B(\logo_top[0] ),
    .Y(_0840_));
 sg13g2_or2_1 _1807_ (.X(_0841_),
    .B(\logo_top[0] ),
    .A(net795));
 sg13g2_nand2_1 _1808_ (.Y(_0842_),
    .A(_0011_),
    .B(_0840_));
 sg13g2_xnor2_1 _1809_ (.Y(_0843_),
    .A(_0761_),
    .B(_0842_));
 sg13g2_nand4_1 _1810_ (.B(\logo_top[0] ),
    .C(_0011_),
    .A(_0760_),
    .Y(_0844_),
    .D(_0012_));
 sg13g2_nor3_1 _1811_ (.A(net789),
    .B(net795),
    .C(_0844_),
    .Y(_0845_));
 sg13g2_nand2_1 _1812_ (.Y(_0846_),
    .A(_0843_),
    .B(_0845_));
 sg13g2_nor4_2 _1813_ (.A(_0832_),
    .B(_0835_),
    .C(_0839_),
    .Y(_0847_),
    .D(_0846_));
 sg13g2_xnor2_1 _1814_ (.Y(_0848_),
    .A(_0014_),
    .B(_0836_));
 sg13g2_nor2b_1 _1815_ (.A(net793),
    .B_N(_0848_),
    .Y(_0849_));
 sg13g2_nor2_1 _1816_ (.A(net794),
    .B(_0833_),
    .Y(_0850_));
 sg13g2_a21oi_1 _1817_ (.A1(\logo_top[4] ),
    .A2(_0828_),
    .Y(_0851_),
    .B1(\logo_top[5] ));
 sg13g2_or2_1 _1818_ (.X(_0852_),
    .B(_0851_),
    .A(_0830_));
 sg13g2_xnor2_1 _1819_ (.Y(_0853_),
    .A(_0012_),
    .B(_0828_));
 sg13g2_nor2_1 _1820_ (.A(_0011_),
    .B(_0826_),
    .Y(_0854_));
 sg13g2_xnor2_1 _1821_ (.Y(_0855_),
    .A(_0761_),
    .B(_0854_));
 sg13g2_nor4_1 _1822_ (.A(_0827_),
    .B(_0852_),
    .C(_0853_),
    .D(_0855_),
    .Y(_0856_));
 sg13g2_and3_1 _1823_ (.X(_0857_),
    .A(_0849_),
    .B(_0850_),
    .C(_0856_));
 sg13g2_nand2_1 _1824_ (.Y(_0858_),
    .A(net790),
    .B(_0857_));
 sg13g2_a21oi_1 _1825_ (.A1(net790),
    .A2(_0857_),
    .Y(_0859_),
    .B1(_0847_));
 sg13g2_nand2_1 _1826_ (.Y(_0860_),
    .A(net803),
    .B(\logo_left[0] ));
 sg13g2_and4_1 _1827_ (.A(\logo_left[3] ),
    .B(\logo_left[2] ),
    .C(net802),
    .D(\logo_left[0] ),
    .X(_0861_));
 sg13g2_nand3_1 _1828_ (.B(net799),
    .C(_0861_),
    .A(\logo_left[5] ),
    .Y(_0862_));
 sg13g2_inv_1 _1829_ (.Y(_0863_),
    .A(_0862_));
 sg13g2_and3_1 _1830_ (.X(_0864_),
    .A(\logo_left[7] ),
    .B(\logo_left[6] ),
    .C(_0863_));
 sg13g2_and2_1 _1831_ (.A(_0792_),
    .B(_0864_),
    .X(_0865_));
 sg13g2_xnor2_1 _1832_ (.Y(_0866_),
    .A(\logo_left[9] ),
    .B(_0865_));
 sg13g2_xor2_1 _1833_ (.B(_0864_),
    .A(\logo_left[8] ),
    .X(_0867_));
 sg13g2_nor2_1 _1834_ (.A(_0009_),
    .B(_0862_),
    .Y(_0868_));
 sg13g2_xnor2_1 _1835_ (.Y(_0869_),
    .A(\logo_left[7] ),
    .B(_0868_));
 sg13g2_a21oi_1 _1836_ (.A1(net799),
    .A2(_0861_),
    .Y(_0870_),
    .B1(net798));
 sg13g2_or2_1 _1837_ (.X(_0871_),
    .B(_0870_),
    .A(_0863_));
 sg13g2_xor2_1 _1838_ (.B(_0861_),
    .A(_0008_),
    .X(_0872_));
 sg13g2_nand2_1 _1839_ (.Y(_0873_),
    .A(_0871_),
    .B(_0872_));
 sg13g2_xor2_1 _1840_ (.B(_0862_),
    .A(net797),
    .X(_0874_));
 sg13g2_nor2_1 _1841_ (.A(_0007_),
    .B(_0860_),
    .Y(_0875_));
 sg13g2_xnor2_1 _1842_ (.Y(_0876_),
    .A(\logo_left[3] ),
    .B(_0875_));
 sg13g2_nand4_1 _1843_ (.B(net801),
    .C(net802),
    .A(net792),
    .Y(_0877_),
    .D(\logo_left[0] ));
 sg13g2_nand2b_1 _1844_ (.Y(_0878_),
    .B(_0876_),
    .A_N(_0877_));
 sg13g2_nor2_1 _1845_ (.A(net802),
    .B(net804),
    .Y(_0879_));
 sg13g2_or2_1 _1846_ (.X(_0880_),
    .B(net801),
    .A(\logo_left[3] ));
 sg13g2_nor3_2 _1847_ (.A(net802),
    .B(net804),
    .C(_0880_),
    .Y(_0881_));
 sg13g2_nor2_2 _1848_ (.A(net798),
    .B(net799),
    .Y(_0882_));
 sg13g2_nand2_1 _1849_ (.Y(_0883_),
    .A(_0881_),
    .B(_0882_));
 sg13g2_or3_1 _1850_ (.A(net796),
    .B(net797),
    .C(_0883_),
    .X(_0884_));
 sg13g2_nor2_1 _1851_ (.A(_0792_),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_xnor2_1 _1852_ (.Y(_0886_),
    .A(_0792_),
    .B(_0884_));
 sg13g2_nand3_1 _1853_ (.B(_0881_),
    .C(_0882_),
    .A(_0009_),
    .Y(_0887_));
 sg13g2_xnor2_1 _1854_ (.Y(_0888_),
    .A(_0009_),
    .B(_0883_));
 sg13g2_nand3_1 _1855_ (.B(_0850_),
    .C(_0856_),
    .A(_0849_),
    .Y(_0889_));
 sg13g2_nand2_1 _1856_ (.Y(_0890_),
    .A(_0007_),
    .B(_0879_));
 sg13g2_xor2_1 _1857_ (.B(_0890_),
    .A(net800),
    .X(_0891_));
 sg13g2_nand2_1 _1858_ (.Y(_0892_),
    .A(net804),
    .B(_0007_));
 sg13g2_nor4_1 _1859_ (.A(net792),
    .B(net796),
    .C(net802),
    .D(_0892_),
    .Y(_0893_));
 sg13g2_nand3_1 _1860_ (.B(_0891_),
    .C(_0893_),
    .A(_0888_),
    .Y(_0894_));
 sg13g2_xor2_1 _1861_ (.B(_0885_),
    .A(\logo_left[9] ),
    .X(_0895_));
 sg13g2_nor2_1 _1862_ (.A(_0873_),
    .B(_0878_),
    .Y(_0896_));
 sg13g2_nand3_1 _1863_ (.B(\logo_left[8] ),
    .C(_0864_),
    .A(\logo_left[9] ),
    .Y(_0897_));
 sg13g2_nand4_1 _1864_ (.B(_0874_),
    .C(_0896_),
    .A(_0869_),
    .Y(_0898_),
    .D(_0897_));
 sg13g2_nor3_1 _1865_ (.A(_0866_),
    .B(_0867_),
    .C(_0898_),
    .Y(_0899_));
 sg13g2_nor4_1 _1866_ (.A(_0873_),
    .B(_0886_),
    .C(_0894_),
    .D(_0895_),
    .Y(_0900_));
 sg13g2_nor2_1 _1867_ (.A(_0899_),
    .B(_0900_),
    .Y(_0901_));
 sg13g2_a21o_2 _1868_ (.A2(_0901_),
    .A1(_0859_),
    .B1(_0825_),
    .X(_0902_));
 sg13g2_xor2_1 _1869_ (.B(_0902_),
    .A(net220),
    .X(_0903_));
 sg13g2_inv_1 _1870_ (.Y(_0904_),
    .A(_0903_));
 sg13g2_and2_1 _1871_ (.A(net809),
    .B(_0903_),
    .X(_0905_));
 sg13g2_nand2b_1 _1872_ (.Y(_0906_),
    .B(_0902_),
    .A_N(net250));
 sg13g2_nand2_1 _1873_ (.Y(_0907_),
    .A(net215),
    .B(\color_index[0] ));
 sg13g2_xor2_1 _1874_ (.B(_0907_),
    .A(_0015_),
    .X(_0908_));
 sg13g2_nand2b_1 _1875_ (.Y(_0909_),
    .B(_0908_),
    .A_N(_0902_));
 sg13g2_nand2_1 _1876_ (.Y(_0910_),
    .A(_0906_),
    .B(_0909_));
 sg13g2_nand2b_1 _1877_ (.Y(_0911_),
    .B(_0902_),
    .A_N(net252));
 sg13g2_nor2_1 _1878_ (.A(\color_index[1] ),
    .B(\color_index[0] ),
    .Y(_0912_));
 sg13g2_nand2b_1 _1879_ (.Y(_0913_),
    .B(_0907_),
    .A_N(_0902_));
 sg13g2_o21ai_1 _1880_ (.B1(_0911_),
    .Y(_0914_),
    .A1(_0912_),
    .A2(_0913_));
 sg13g2_nand2_1 _1881_ (.Y(_0915_),
    .A(_0910_),
    .B(_0914_));
 sg13g2_nand2_1 _1882_ (.Y(_0000_),
    .A(_0905_),
    .B(_0915_));
 sg13g2_nand2_1 _1883_ (.Y(_0916_),
    .A(_0905_),
    .B(_0910_));
 sg13g2_nand2_1 _1884_ (.Y(_0917_),
    .A(net809),
    .B(_0914_));
 sg13g2_mux2_1 _1885_ (.A0(_0914_),
    .A1(_0917_),
    .S(_0916_),
    .X(_0001_));
 sg13g2_nor2_1 _1886_ (.A(_0910_),
    .B(_0917_),
    .Y(_0918_));
 sg13g2_mux2_1 _1887_ (.A0(_0905_),
    .A1(_0904_),
    .S(_0918_),
    .X(_0002_));
 sg13g2_a21o_1 _1888_ (.A2(_0910_),
    .A1(net808),
    .B1(_0905_),
    .X(_0116_));
 sg13g2_nand2_1 _1889_ (.Y(_0919_),
    .A(_0916_),
    .B(_0116_));
 sg13g2_or2_1 _1890_ (.X(_0003_),
    .B(_0919_),
    .A(_0918_));
 sg13g2_nor2b_1 _1891_ (.A(\logo_top[3] ),
    .B_N(net782),
    .Y(_0920_));
 sg13g2_xnor2_1 _1892_ (.Y(_0921_),
    .A(\logo_top[3] ),
    .B(net782));
 sg13g2_nor2_1 _1893_ (.A(\logo_top[2] ),
    .B(_0770_),
    .Y(_0922_));
 sg13g2_nor2b_1 _1894_ (.A(net795),
    .B_N(\pix_y[1] ),
    .Y(_0923_));
 sg13g2_nand2b_2 _1895_ (.Y(_0924_),
    .B(\logo_top[0] ),
    .A_N(\pix_y[0] ));
 sg13g2_xnor2_1 _1896_ (.Y(_0925_),
    .A(net795),
    .B(\pix_y[1] ));
 sg13g2_a21o_1 _1897_ (.A2(_0925_),
    .A1(_0924_),
    .B1(_0923_),
    .X(_0926_));
 sg13g2_xnor2_1 _1898_ (.Y(_0927_),
    .A(\logo_top[2] ),
    .B(\pix_y[2] ));
 sg13g2_a21o_2 _1899_ (.A2(_0927_),
    .A1(_0926_),
    .B1(_0922_),
    .X(_0928_));
 sg13g2_xor2_1 _1900_ (.B(_0928_),
    .A(_0921_),
    .X(_0929_));
 sg13g2_xnor2_1 _1901_ (.Y(_0930_),
    .A(_0921_),
    .B(_0928_));
 sg13g2_xor2_1 _1902_ (.B(_0927_),
    .A(_0926_),
    .X(_0931_));
 sg13g2_xnor2_1 _1903_ (.Y(_0932_),
    .A(_0926_),
    .B(_0927_));
 sg13g2_nor2_1 _1904_ (.A(net718),
    .B(net741),
    .Y(_0933_));
 sg13g2_nand2_2 _1905_ (.Y(_0934_),
    .A(net726),
    .B(net746));
 sg13g2_nor2b_1 _1906_ (.A(net799),
    .B_N(\pix_x[4] ),
    .Y(_0935_));
 sg13g2_nor2b_1 _1907_ (.A(net803),
    .B_N(\pix_x[1] ),
    .Y(_0936_));
 sg13g2_nand2b_2 _1908_ (.Y(_0937_),
    .B(net804),
    .A_N(\pix_x[0] ));
 sg13g2_xnor2_1 _1909_ (.Y(_0938_),
    .A(net803),
    .B(\pix_x[1] ));
 sg13g2_a21oi_2 _1910_ (.B1(_0936_),
    .Y(_0939_),
    .A2(_0938_),
    .A1(_0937_));
 sg13g2_a21o_1 _1911_ (.A2(_0938_),
    .A1(_0937_),
    .B1(_0936_),
    .X(_0940_));
 sg13g2_nor2b_1 _1912_ (.A(net800),
    .B_N(\pix_x[3] ),
    .Y(_0941_));
 sg13g2_xnor2_1 _1913_ (.Y(_0942_),
    .A(net800),
    .B(\pix_x[3] ));
 sg13g2_nor2b_1 _1914_ (.A(net801),
    .B_N(\pix_x[2] ),
    .Y(_0943_));
 sg13g2_xnor2_1 _1915_ (.Y(_0944_),
    .A(net801),
    .B(\pix_x[2] ));
 sg13g2_nand2_1 _1916_ (.Y(_0945_),
    .A(_0942_),
    .B(_0944_));
 sg13g2_a21oi_1 _1917_ (.A1(_0942_),
    .A2(_0943_),
    .Y(_0946_),
    .B1(_0941_));
 sg13g2_o21ai_1 _1918_ (.B1(_0946_),
    .Y(_0947_),
    .A1(_0939_),
    .A2(_0945_));
 sg13g2_xnor2_1 _1919_ (.Y(_0948_),
    .A(net799),
    .B(\pix_x[4] ));
 sg13g2_a21o_1 _1920_ (.A2(_0948_),
    .A1(_0947_),
    .B1(_0935_),
    .X(_0949_));
 sg13g2_nor2b_1 _1921_ (.A(net798),
    .B_N(\pix_x[5] ),
    .Y(_0950_));
 sg13g2_nor2_2 _1922_ (.A(_0764_),
    .B(\pix_x[5] ),
    .Y(_0951_));
 sg13g2_inv_1 _1923_ (.Y(_0952_),
    .A(_0951_));
 sg13g2_nor2_1 _1924_ (.A(_0950_),
    .B(_0951_),
    .Y(_0953_));
 sg13g2_xor2_1 _1925_ (.B(_0953_),
    .A(_0949_),
    .X(_0954_));
 sg13g2_xnor2_1 _1926_ (.Y(_0955_),
    .A(_0949_),
    .B(_0953_));
 sg13g2_a21oi_2 _1927_ (.B1(_0943_),
    .Y(_0956_),
    .A2(_0944_),
    .A1(_0940_));
 sg13g2_xor2_1 _1928_ (.B(_0956_),
    .A(_0942_),
    .X(_0957_));
 sg13g2_xnor2_1 _1929_ (.Y(_0958_),
    .A(_0942_),
    .B(_0956_));
 sg13g2_nand2_2 _1930_ (.Y(_0959_),
    .A(net696),
    .B(net713));
 sg13g2_xor2_1 _1931_ (.B(_0948_),
    .A(_0947_),
    .X(_0960_));
 sg13g2_xnor2_1 _1932_ (.Y(_0961_),
    .A(_0947_),
    .B(_0948_));
 sg13g2_nor2_2 _1933_ (.A(net714),
    .B(net708),
    .Y(_0962_));
 sg13g2_nand2_1 _1934_ (.Y(_0963_),
    .A(net715),
    .B(net711));
 sg13g2_nor2_2 _1935_ (.A(net713),
    .B(net711),
    .Y(_0964_));
 sg13g2_nand2_2 _1936_ (.Y(_0965_),
    .A(net715),
    .B(net710));
 sg13g2_nor2_1 _1937_ (.A(net695),
    .B(net716),
    .Y(_0966_));
 sg13g2_nand2_2 _1938_ (.Y(_0967_),
    .A(net703),
    .B(net714));
 sg13g2_a21oi_2 _1939_ (.B1(_0962_),
    .Y(_0968_),
    .A2(net714),
    .A1(net695));
 sg13g2_nand2b_1 _1940_ (.Y(_0969_),
    .B(net797),
    .A_N(\pix_x[6] ));
 sg13g2_nand2b_1 _1941_ (.Y(_0970_),
    .B(\pix_x[6] ),
    .A_N(net797));
 sg13g2_and2_1 _1942_ (.A(_0969_),
    .B(_0970_),
    .X(_0971_));
 sg13g2_nand2_1 _1943_ (.Y(_0972_),
    .A(_0969_),
    .B(_0970_));
 sg13g2_a221oi_1 _1944_ (.B2(_0948_),
    .C1(_0935_),
    .B1(_0947_),
    .A1(_0764_),
    .Y(_0973_),
    .A2(\pix_x[5] ));
 sg13g2_nor3_2 _1945_ (.A(_0951_),
    .B(_0972_),
    .C(_0973_),
    .Y(_0974_));
 sg13g2_or3_1 _1946_ (.A(_0951_),
    .B(_0972_),
    .C(_0973_),
    .X(_0975_));
 sg13g2_a221oi_1 _1947_ (.B2(_0970_),
    .C1(_0950_),
    .B1(_0969_),
    .A1(_0949_),
    .Y(_0976_),
    .A2(_0952_));
 sg13g2_o21ai_1 _1948_ (.B1(_0972_),
    .Y(_0977_),
    .A1(_0951_),
    .A2(_0973_));
 sg13g2_o21ai_1 _1949_ (.B1(_0971_),
    .Y(_0978_),
    .A1(_0951_),
    .A2(_0973_));
 sg13g2_or3_1 _1950_ (.A(_0951_),
    .B(_0971_),
    .C(_0973_),
    .X(_0979_));
 sg13g2_nor2_1 _1951_ (.A(_0974_),
    .B(_0976_),
    .Y(_0980_));
 sg13g2_nand2_1 _1952_ (.Y(_0981_),
    .A(net687),
    .B(net683));
 sg13g2_nor2_2 _1953_ (.A(net716),
    .B(_0960_),
    .Y(_0982_));
 sg13g2_inv_1 _1954_ (.Y(_0983_),
    .A(_0982_));
 sg13g2_a22oi_1 _1955_ (.Y(_0984_),
    .B1(_0982_),
    .B2(net695),
    .A2(net683),
    .A1(net688));
 sg13g2_inv_1 _1956_ (.Y(_0985_),
    .A(net643));
 sg13g2_or2_1 _1957_ (.X(_0986_),
    .B(net643),
    .A(_0968_));
 sg13g2_xor2_1 _1958_ (.B(_0925_),
    .A(_0924_),
    .X(_0987_));
 sg13g2_xnor2_1 _1959_ (.Y(_0988_),
    .A(_0924_),
    .B(_0925_));
 sg13g2_nand2b_2 _1960_ (.Y(_0989_),
    .B(\pix_y[0] ),
    .A_N(\logo_top[0] ));
 sg13g2_and2_1 _1961_ (.A(_0924_),
    .B(_0989_),
    .X(_0990_));
 sg13g2_nand2_2 _1962_ (.Y(_0991_),
    .A(_0924_),
    .B(_0989_));
 sg13g2_nor2_1 _1963_ (.A(net766),
    .B(net760),
    .Y(_0992_));
 sg13g2_nand2_1 _1964_ (.Y(_0993_),
    .A(net773),
    .B(net755));
 sg13g2_nor3_1 _1965_ (.A(net711),
    .B(net690),
    .C(net685),
    .Y(_0994_));
 sg13g2_nand3_1 _1966_ (.B(net687),
    .C(net682),
    .A(net708),
    .Y(_0995_));
 sg13g2_nor4_2 _1967_ (.A(net692),
    .B(net715),
    .C(net690),
    .Y(_0996_),
    .D(net685));
 sg13g2_nor2_1 _1968_ (.A(net641),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_or3_1 _1969_ (.A(net643),
    .B(net640),
    .C(_0996_),
    .X(_0998_));
 sg13g2_nor2_1 _1970_ (.A(net773),
    .B(net756),
    .Y(_0999_));
 sg13g2_nand2_1 _1971_ (.Y(_1000_),
    .A(net763),
    .B(net757));
 sg13g2_nor2_1 _1972_ (.A(net715),
    .B(net710),
    .Y(_1001_));
 sg13g2_nand2_2 _1973_ (.Y(_1002_),
    .A(net713),
    .B(net711));
 sg13g2_nand2_2 _1974_ (.Y(_1003_),
    .A(net695),
    .B(net677));
 sg13g2_nand2_2 _1975_ (.Y(_1004_),
    .A(net703),
    .B(net716));
 sg13g2_inv_1 _1976_ (.Y(_1005_),
    .A(_1004_));
 sg13g2_a22oi_1 _1977_ (.Y(_1006_),
    .B1(net681),
    .B2(net679),
    .A2(net716),
    .A1(net703));
 sg13g2_nand2_1 _1978_ (.Y(_1007_),
    .A(_1003_),
    .B(_1006_));
 sg13g2_nand2_2 _1979_ (.Y(_1008_),
    .A(net701),
    .B(net712));
 sg13g2_nand2_1 _1980_ (.Y(_1009_),
    .A(net698),
    .B(_0962_));
 sg13g2_a22oi_1 _1981_ (.Y(_1010_),
    .B1(net681),
    .B2(net679),
    .A2(_0962_),
    .A1(net702));
 sg13g2_nand2_1 _1982_ (.Y(_1011_),
    .A(_1003_),
    .B(_1010_));
 sg13g2_and2_1 _1983_ (.A(_1003_),
    .B(_1010_),
    .X(_1012_));
 sg13g2_a22oi_1 _1984_ (.Y(_1013_),
    .B1(net733),
    .B2(_1012_),
    .A2(_0998_),
    .A1(net736));
 sg13g2_a221oi_1 _1985_ (.B2(_1012_),
    .C1(_0986_),
    .B1(net733),
    .A1(net736),
    .Y(_1014_),
    .A2(_0998_));
 sg13g2_nor2_1 _1986_ (.A(_0934_),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_nand2_1 _1987_ (.Y(_1016_),
    .A(net693),
    .B(net710));
 sg13g2_a22oi_1 _1988_ (.Y(_1017_),
    .B1(net688),
    .B2(net683),
    .A2(net709),
    .A1(net695));
 sg13g2_nand2_1 _1989_ (.Y(_1018_),
    .A(net645),
    .B(_1016_));
 sg13g2_a21oi_1 _1990_ (.A1(_1003_),
    .A2(_1010_),
    .Y(_1019_),
    .B1(_1017_));
 sg13g2_nor2_2 _1991_ (.A(net721),
    .B(net746),
    .Y(_1020_));
 sg13g2_nand2_2 _1992_ (.Y(_1021_),
    .A(net725),
    .B(net743));
 sg13g2_nor2_1 _1993_ (.A(net726),
    .B(net742),
    .Y(_1022_));
 sg13g2_nand2_1 _1994_ (.Y(_1023_),
    .A(net719),
    .B(net745));
 sg13g2_nor2_2 _1995_ (.A(net743),
    .B(net767),
    .Y(_1024_));
 sg13g2_nand2_2 _1996_ (.Y(_1025_),
    .A(net744),
    .B(net774));
 sg13g2_nor2_1 _1997_ (.A(net725),
    .B(_1025_),
    .Y(_1026_));
 sg13g2_nand2_1 _1998_ (.Y(_1027_),
    .A(net719),
    .B(_1024_));
 sg13g2_nand2_2 _1999_ (.Y(_1028_),
    .A(net744),
    .B(net754));
 sg13g2_nor2_1 _2000_ (.A(net741),
    .B(net734),
    .Y(_1029_));
 sg13g2_nand2_2 _2001_ (.Y(_1030_),
    .A(net745),
    .B(net739));
 sg13g2_nor2_2 _2002_ (.A(net723),
    .B(_1030_),
    .Y(_1031_));
 sg13g2_nand2_1 _2003_ (.Y(_1032_),
    .A(net693),
    .B(net675));
 sg13g2_a22oi_1 _2004_ (.Y(_1033_),
    .B1(net675),
    .B2(net692),
    .A2(net684),
    .A1(net686));
 sg13g2_inv_1 _2005_ (.Y(_1034_),
    .A(_1033_));
 sg13g2_nor2_2 _2006_ (.A(net640),
    .B(net637),
    .Y(_1035_));
 sg13g2_or2_1 _2007_ (.X(_1036_),
    .B(net637),
    .A(net640));
 sg13g2_nor2_1 _2008_ (.A(_0996_),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_a21oi_2 _2009_ (.B1(_0920_),
    .Y(_1038_),
    .A2(_0928_),
    .A1(_0921_));
 sg13g2_nand2b_1 _2010_ (.Y(_1039_),
    .B(\pix_y[4] ),
    .A_N(\logo_top[4] ));
 sg13g2_xor2_1 _2011_ (.B(\pix_y[4] ),
    .A(\logo_top[4] ),
    .X(_1040_));
 sg13g2_xor2_1 _2012_ (.B(_1040_),
    .A(_1038_),
    .X(_1041_));
 sg13g2_xnor2_1 _2013_ (.Y(_1042_),
    .A(_1038_),
    .B(_1040_));
 sg13g2_nor2_1 _2014_ (.A(net767),
    .B(net755),
    .Y(_1043_));
 sg13g2_nand2_2 _2015_ (.Y(_1044_),
    .A(net773),
    .B(net760));
 sg13g2_o21ai_1 _2016_ (.B1(net729),
    .Y(_1045_),
    .A1(net643),
    .A2(_1010_));
 sg13g2_o21ai_1 _2017_ (.B1(_1037_),
    .Y(_1046_),
    .A1(net735),
    .A2(_1019_));
 sg13g2_nand2_1 _2018_ (.Y(_1047_),
    .A(_1019_),
    .B(_1045_));
 sg13g2_a221oi_1 _2019_ (.B2(_1020_),
    .C1(net665),
    .B1(_1047_),
    .A1(net673),
    .Y(_1048_),
    .A2(_1046_));
 sg13g2_nor2_2 _2020_ (.A(net767),
    .B(_1021_),
    .Y(_1049_));
 sg13g2_a21oi_1 _2021_ (.A1(_0985_),
    .A2(_1011_),
    .Y(_1050_),
    .B1(net760));
 sg13g2_nor2_1 _2022_ (.A(net726),
    .B(net746),
    .Y(_1051_));
 sg13g2_nand2_1 _2023_ (.Y(_1052_),
    .A(net721),
    .B(net742));
 sg13g2_nand2_1 _2024_ (.Y(_1053_),
    .A(net773),
    .B(_0996_));
 sg13g2_o21ai_1 _2025_ (.B1(net675),
    .Y(_1054_),
    .A1(net696),
    .A2(net714));
 sg13g2_a21oi_2 _2026_ (.B1(net640),
    .Y(_1055_),
    .A2(_1054_),
    .A1(net647));
 sg13g2_a21o_1 _2027_ (.A2(_1054_),
    .A1(net647),
    .B1(net640),
    .X(_1056_));
 sg13g2_nand3_1 _2028_ (.B(_1053_),
    .C(_1055_),
    .A(net735),
    .Y(_1057_));
 sg13g2_a21oi_1 _2029_ (.A1(net739),
    .A2(_1037_),
    .Y(_1058_),
    .B1(net658));
 sg13g2_a221oi_1 _2030_ (.B2(_1058_),
    .C1(_1015_),
    .B1(_1057_),
    .A1(_1049_),
    .Y(_1059_),
    .A2(_1050_));
 sg13g2_o21ai_1 _2031_ (.B1(_1039_),
    .Y(_1060_),
    .A1(_1038_),
    .A2(_1040_));
 sg13g2_xnor2_1 _2032_ (.Y(_1061_),
    .A(\logo_top[5] ),
    .B(\pix_y[5] ));
 sg13g2_xnor2_1 _2033_ (.Y(_1062_),
    .A(_1060_),
    .B(_1061_));
 sg13g2_xor2_1 _2034_ (.B(_1061_),
    .A(_1060_),
    .X(_1063_));
 sg13g2_nor2_2 _2035_ (.A(net743),
    .B(net774),
    .Y(_1064_));
 sg13g2_nand2_2 _2036_ (.Y(_1065_),
    .A(net746),
    .B(net767));
 sg13g2_nor2_1 _2037_ (.A(net726),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_nand2_1 _2038_ (.Y(_1067_),
    .A(net702),
    .B(net708));
 sg13g2_and4_1 _2039_ (.A(net702),
    .B(net708),
    .C(net681),
    .D(net679),
    .X(_1068_));
 sg13g2_nand2b_1 _2040_ (.Y(_1069_),
    .B(net648),
    .A_N(_1067_));
 sg13g2_xnor2_1 _2041_ (.Y(_1070_),
    .A(net702),
    .B(net716));
 sg13g2_nand2_1 _2042_ (.Y(_1071_),
    .A(net641),
    .B(_1070_));
 sg13g2_nand2_1 _2043_ (.Y(_1072_),
    .A(_1069_),
    .B(_1071_));
 sg13g2_a22oi_1 _2044_ (.Y(_1073_),
    .B1(net686),
    .B2(net684),
    .A2(net710),
    .A1(net698));
 sg13g2_nand2_2 _2045_ (.Y(_1074_),
    .A(net693),
    .B(_0965_));
 sg13g2_xnor2_1 _2046_ (.Y(_1075_),
    .A(net715),
    .B(net712));
 sg13g2_xnor2_1 _2047_ (.Y(_1076_),
    .A(net713),
    .B(net712));
 sg13g2_nand2_1 _2048_ (.Y(_1077_),
    .A(net696),
    .B(net656));
 sg13g2_a22oi_1 _2049_ (.Y(_1078_),
    .B1(net681),
    .B2(net679),
    .A2(_0964_),
    .A1(net703));
 sg13g2_a21oi_2 _2050_ (.B1(net632),
    .Y(_1079_),
    .A2(_1078_),
    .A1(_1077_));
 sg13g2_a21oi_1 _2051_ (.A1(net762),
    .A2(_1079_),
    .Y(_1080_),
    .B1(_1072_));
 sg13g2_nand2b_1 _2052_ (.Y(_1081_),
    .B(_1066_),
    .A_N(_1080_));
 sg13g2_a21oi_1 _2053_ (.A1(net661),
    .A2(_1079_),
    .Y(_1082_),
    .B1(net668));
 sg13g2_nand2_2 _2054_ (.Y(_1083_),
    .A(net699),
    .B(_0965_));
 sg13g2_mux2_2 _2055_ (.A0(net691),
    .A1(net676),
    .S(net692),
    .X(_1084_));
 sg13g2_mux2_2 _2056_ (.A0(_0965_),
    .A1(net675),
    .S(net693),
    .X(_1085_));
 sg13g2_a21oi_1 _2057_ (.A1(net647),
    .A2(_1084_),
    .Y(_1086_),
    .B1(net640));
 sg13g2_o21ai_1 _2058_ (.B1(_0995_),
    .Y(_1087_),
    .A1(net652),
    .A2(_1085_));
 sg13g2_nor2_1 _2059_ (.A(net742),
    .B(_1086_),
    .Y(_1088_));
 sg13g2_nor2_1 _2060_ (.A(_1030_),
    .B(_1055_),
    .Y(_1089_));
 sg13g2_o21ai_1 _2061_ (.B1(net725),
    .Y(_1090_),
    .A1(_1088_),
    .A2(_1089_));
 sg13g2_a21oi_1 _2062_ (.A1(_0966_),
    .A2(net766),
    .Y(_1091_),
    .B1(_1086_));
 sg13g2_nor2_2 _2063_ (.A(net755),
    .B(_1068_),
    .Y(_1092_));
 sg13g2_a21oi_2 _2064_ (.B1(net761),
    .Y(_1093_),
    .A2(_1084_),
    .A1(net647));
 sg13g2_o21ai_1 _2065_ (.B1(_1071_),
    .Y(_1094_),
    .A1(_1092_),
    .A2(_1093_));
 sg13g2_a22oi_1 _2066_ (.Y(_1095_),
    .B1(_1094_),
    .B2(_1026_),
    .A2(_1091_),
    .A1(_1020_));
 sg13g2_and3_1 _2067_ (.X(_1096_),
    .A(_1082_),
    .B(_1090_),
    .C(_1095_));
 sg13g2_a221oi_1 _2068_ (.B2(_1096_),
    .C1(net633),
    .B1(_1081_),
    .A1(_1048_),
    .Y(_1097_),
    .A2(_1059_));
 sg13g2_xor2_1 _2069_ (.B(\pix_y[6] ),
    .A(\logo_top[6] ),
    .X(_1098_));
 sg13g2_a21oi_1 _2070_ (.A1(_0760_),
    .A2(\pix_y[5] ),
    .Y(_1099_),
    .B1(_1060_));
 sg13g2_a21oi_2 _2071_ (.B1(_1099_),
    .Y(_1100_),
    .A2(_0771_),
    .A1(\logo_top[5] ));
 sg13g2_nand2b_1 _2072_ (.Y(_1101_),
    .B(_1100_),
    .A_N(_1098_));
 sg13g2_xnor2_1 _2073_ (.Y(_1102_),
    .A(_1098_),
    .B(_1100_));
 sg13g2_xor2_1 _2074_ (.B(_1100_),
    .A(_1098_),
    .X(_1103_));
 sg13g2_o21ai_1 _2075_ (.B1(net732),
    .Y(_1104_),
    .A1(_0968_),
    .A2(net644));
 sg13g2_nor2_2 _2076_ (.A(net774),
    .B(net761),
    .Y(_1105_));
 sg13g2_nand2_2 _2077_ (.Y(_1106_),
    .A(net766),
    .B(net755));
 sg13g2_nor3_2 _2078_ (.A(net693),
    .B(net690),
    .C(net685),
    .Y(_1107_));
 sg13g2_nand3_1 _2079_ (.B(net686),
    .C(net684),
    .A(net698),
    .Y(_1108_));
 sg13g2_xnor2_1 _2080_ (.Y(_1109_),
    .A(net692),
    .B(net691));
 sg13g2_xnor2_1 _2081_ (.Y(_1110_),
    .A(net698),
    .B(net691));
 sg13g2_o21ai_1 _2082_ (.B1(_1108_),
    .Y(_1111_),
    .A1(net649),
    .A2(_1110_));
 sg13g2_a22oi_1 _2083_ (.Y(_1112_),
    .B1(_1109_),
    .B2(net646),
    .A2(net628),
    .A1(_0963_));
 sg13g2_o21ai_1 _2084_ (.B1(_1104_),
    .Y(_1113_),
    .A1(_1106_),
    .A2(_1112_));
 sg13g2_a21oi_1 _2085_ (.A1(net688),
    .A2(net682),
    .Y(_1114_),
    .B1(_1075_));
 sg13g2_a221oi_1 _2086_ (.B2(net682),
    .C1(net656),
    .B1(net687),
    .A1(net696),
    .Y(_1115_),
    .A2(net708));
 sg13g2_nand3b_1 _2087_ (.B(net737),
    .C(_1074_),
    .Y(_1116_),
    .A_N(_1115_));
 sg13g2_o21ai_1 _2088_ (.B1(_1116_),
    .Y(_1117_),
    .A1(_1044_),
    .A2(_1112_));
 sg13g2_o21ai_1 _2089_ (.B1(net660),
    .Y(_1118_),
    .A1(_1113_),
    .A2(_1117_));
 sg13g2_nand2_1 _2090_ (.Y(_1119_),
    .A(net702),
    .B(_1076_));
 sg13g2_nor2_1 _2091_ (.A(net712),
    .B(_1070_),
    .Y(_1120_));
 sg13g2_mux2_2 _2092_ (.A0(_0964_),
    .A1(net656),
    .S(net702),
    .X(_1121_));
 sg13g2_nand2_1 _2093_ (.Y(_1122_),
    .A(net733),
    .B(_1121_));
 sg13g2_nor4_2 _2094_ (.A(net692),
    .B(net691),
    .C(net690),
    .Y(_1123_),
    .D(net685));
 sg13g2_nand4_1 _2095_ (.B(_0965_),
    .C(net686),
    .A(net699),
    .Y(_1124_),
    .D(net684));
 sg13g2_nor3_1 _2096_ (.A(net712),
    .B(net653),
    .C(_1070_),
    .Y(_1125_));
 sg13g2_o21ai_1 _2097_ (.B1(net735),
    .Y(_1126_),
    .A1(_1123_),
    .A2(_1125_));
 sg13g2_a21o_1 _2098_ (.A2(_1126_),
    .A1(_1122_),
    .B1(net671),
    .X(_1127_));
 sg13g2_xnor2_1 _2099_ (.Y(_1128_),
    .A(net692),
    .B(net711));
 sg13g2_xnor2_1 _2100_ (.Y(_1129_),
    .A(net699),
    .B(net711));
 sg13g2_a21oi_2 _2101_ (.B1(net627),
    .Y(_1130_),
    .A2(_1129_),
    .A1(net645));
 sg13g2_o21ai_1 _2102_ (.B1(_1124_),
    .Y(_1131_),
    .A1(net649),
    .A2(_1128_));
 sg13g2_nor2_2 _2103_ (.A(net744),
    .B(net774),
    .Y(_1132_));
 sg13g2_nand2_2 _2104_ (.Y(_1133_),
    .A(net740),
    .B(net763));
 sg13g2_nand2_1 _2105_ (.Y(_1134_),
    .A(_1131_),
    .B(_1133_));
 sg13g2_nand2_1 _2106_ (.Y(_1135_),
    .A(net701),
    .B(net676));
 sg13g2_and4_2 _2107_ (.A(net700),
    .B(net713),
    .C(net681),
    .D(net679),
    .X(_1136_));
 sg13g2_and4_2 _2108_ (.A(net698),
    .B(net680),
    .C(net678),
    .D(net676),
    .X(_1137_));
 sg13g2_nand4_1 _2109_ (.B(net680),
    .C(net678),
    .A(net700),
    .Y(_1138_),
    .D(net677));
 sg13g2_and4_2 _2110_ (.A(net692),
    .B(net710),
    .C(net680),
    .D(net678),
    .X(_1139_));
 sg13g2_nand4_1 _2111_ (.B(net710),
    .C(net680),
    .A(net694),
    .Y(_1140_),
    .D(net678));
 sg13g2_nor2_2 _2112_ (.A(net627),
    .B(_1139_),
    .Y(_1141_));
 sg13g2_nand2_2 _2113_ (.Y(_1142_),
    .A(_1124_),
    .B(_1140_));
 sg13g2_nor3_2 _2114_ (.A(net627),
    .B(_1137_),
    .C(_1139_),
    .Y(_1143_));
 sg13g2_nand2_1 _2115_ (.Y(_1144_),
    .A(_1138_),
    .B(_1141_));
 sg13g2_o21ai_1 _2116_ (.B1(_1143_),
    .Y(_1145_),
    .A1(_1130_),
    .A2(_1132_));
 sg13g2_a21oi_1 _2117_ (.A1(net723),
    .A2(_1145_),
    .Y(_1146_),
    .B1(net667));
 sg13g2_nand2_1 _2118_ (.Y(_1147_),
    .A(_1031_),
    .B(_1144_));
 sg13g2_nand4_1 _2119_ (.B(_1127_),
    .C(_1146_),
    .A(_1118_),
    .Y(_1148_),
    .D(_1147_));
 sg13g2_nor3_2 _2120_ (.A(net698),
    .B(net690),
    .C(net685),
    .Y(_1149_));
 sg13g2_nand3_1 _2121_ (.B(net687),
    .C(net682),
    .A(net695),
    .Y(_1150_));
 sg13g2_nor2_2 _2122_ (.A(net631),
    .B(net628),
    .Y(_1151_));
 sg13g2_nor2_1 _2123_ (.A(net730),
    .B(_1151_),
    .Y(_1152_));
 sg13g2_nand2_1 _2124_ (.Y(_1153_),
    .A(net733),
    .B(_1003_));
 sg13g2_nor2_1 _2125_ (.A(_1151_),
    .B(_1153_),
    .Y(_1154_));
 sg13g2_a21oi_2 _2126_ (.B1(net628),
    .Y(_1155_),
    .A2(net630),
    .A1(net675));
 sg13g2_nor2_1 _2127_ (.A(_1106_),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_o21ai_1 _2128_ (.B1(net673),
    .Y(_1157_),
    .A1(_1154_),
    .A2(_1156_));
 sg13g2_nand4_1 _2129_ (.B(net687),
    .C(net682),
    .A(net695),
    .Y(_1158_),
    .D(_1002_));
 sg13g2_and3_1 _2130_ (.X(_1159_),
    .A(net772),
    .B(_1138_),
    .C(_1158_));
 sg13g2_a22oi_1 _2131_ (.Y(_1160_),
    .B1(_1076_),
    .B2(net702),
    .A2(net682),
    .A1(net687));
 sg13g2_nor3_2 _2132_ (.A(net690),
    .B(net685),
    .C(net757),
    .Y(_1161_));
 sg13g2_nor3_2 _2133_ (.A(net690),
    .B(net685),
    .C(net675),
    .Y(_1162_));
 sg13g2_nand3_1 _2134_ (.B(net684),
    .C(net676),
    .A(net686),
    .Y(_1163_));
 sg13g2_nor2_1 _2135_ (.A(net759),
    .B(_1163_),
    .Y(_1164_));
 sg13g2_or4_1 _2136_ (.A(net628),
    .B(_1159_),
    .C(_1160_),
    .D(_1164_),
    .X(_1165_));
 sg13g2_nand4_1 _2137_ (.B(net708),
    .C(net688),
    .A(net695),
    .Y(_1166_),
    .D(net683));
 sg13g2_a21oi_2 _2138_ (.B1(net699),
    .Y(_1167_),
    .A2(net684),
    .A1(net686));
 sg13g2_o21ai_1 _2139_ (.B1(net693),
    .Y(_1168_),
    .A1(net690),
    .A2(net685));
 sg13g2_nor2_2 _2140_ (.A(net628),
    .B(_1167_),
    .Y(_1169_));
 sg13g2_nand2_1 _2141_ (.Y(_1170_),
    .A(_1138_),
    .B(_1166_));
 sg13g2_a22oi_1 _2142_ (.Y(_1171_),
    .B1(net676),
    .B2(net698),
    .A2(net684),
    .A1(net686));
 sg13g2_a22oi_1 _2143_ (.Y(_1172_),
    .B1(net680),
    .B2(net678),
    .A2(net691),
    .A1(net692));
 sg13g2_o21ai_1 _2144_ (.B1(net737),
    .Y(_1173_),
    .A1(_1171_),
    .A2(_1172_));
 sg13g2_nand2_1 _2145_ (.Y(_1174_),
    .A(_1170_),
    .B(_1173_));
 sg13g2_a22oi_1 _2146_ (.Y(_1175_),
    .B1(_1174_),
    .B2(net705),
    .A2(_1165_),
    .A1(net674));
 sg13g2_o21ai_1 _2147_ (.B1(_1003_),
    .Y(_1176_),
    .A1(net631),
    .A2(_1123_));
 sg13g2_o21ai_1 _2148_ (.B1(net668),
    .Y(_1177_),
    .A1(net658),
    .A2(_1176_));
 sg13g2_inv_1 _2149_ (.Y(_1178_),
    .A(_1177_));
 sg13g2_nand3_1 _2150_ (.B(_1108_),
    .C(_1168_),
    .A(_1009_),
    .Y(_1179_));
 sg13g2_a21oi_1 _2151_ (.A1(_1026_),
    .A2(_1179_),
    .Y(_1180_),
    .B1(_1177_));
 sg13g2_nand3_1 _2152_ (.B(_1175_),
    .C(_1180_),
    .A(_1157_),
    .Y(_1181_));
 sg13g2_nand3_1 _2153_ (.B(_1148_),
    .C(_1181_),
    .A(_1063_),
    .Y(_1182_));
 sg13g2_nand3b_1 _2154_ (.B(net618),
    .C(_1182_),
    .Y(_1183_),
    .A_N(_1097_));
 sg13g2_xnor2_1 _2155_ (.Y(_1184_),
    .A(net804),
    .B(\pix_x[0] ));
 sg13g2_xor2_1 _2156_ (.B(\pix_x[0] ),
    .A(net804),
    .X(_1185_));
 sg13g2_nand2_2 _2157_ (.Y(_1186_),
    .A(net632),
    .B(net629));
 sg13g2_a21oi_2 _2158_ (.B1(_1162_),
    .Y(_1187_),
    .A2(_1074_),
    .A1(net632));
 sg13g2_a221oi_1 _2159_ (.B2(net629),
    .C1(net758),
    .B1(net632),
    .A1(net650),
    .Y(_1188_),
    .A2(net676));
 sg13g2_nor3_2 _2160_ (.A(_0974_),
    .B(_0976_),
    .C(net676),
    .Y(_1189_));
 sg13g2_and2_1 _2161_ (.A(net758),
    .B(_1189_),
    .X(_1190_));
 sg13g2_o21ai_1 _2162_ (.B1(net724),
    .Y(_1191_),
    .A1(_1188_),
    .A2(_1190_));
 sg13g2_nand2_2 _2163_ (.Y(_1192_),
    .A(net638),
    .B(_1189_));
 sg13g2_a21oi_1 _2164_ (.A1(_1025_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(_1191_));
 sg13g2_and2_1 _2165_ (.A(net638),
    .B(_1172_),
    .X(_1194_));
 sg13g2_nand2_1 _2166_ (.Y(_1195_),
    .A(net638),
    .B(_1172_));
 sg13g2_a21oi_1 _2167_ (.A1(net650),
    .A2(_1110_),
    .Y(_1196_),
    .B1(net758));
 sg13g2_o21ai_1 _2168_ (.B1(net753),
    .Y(_1197_),
    .A1(net646),
    .A2(_1109_));
 sg13g2_a21oi_2 _2169_ (.B1(net770),
    .Y(_1198_),
    .A2(_1197_),
    .A1(_1141_));
 sg13g2_nor2_1 _2170_ (.A(net734),
    .B(_1194_),
    .Y(_1199_));
 sg13g2_o21ai_1 _2171_ (.B1(net728),
    .Y(_1200_),
    .A1(net645),
    .A2(_1109_));
 sg13g2_nor3_1 _2172_ (.A(net659),
    .B(_1198_),
    .C(_1199_),
    .Y(_1201_));
 sg13g2_a22oi_1 _2173_ (.Y(_1202_),
    .B1(_1200_),
    .B2(_1201_),
    .A2(_1194_),
    .A1(net672));
 sg13g2_a21oi_2 _2174_ (.B1(net631),
    .Y(_1203_),
    .A2(_1109_),
    .A1(net652));
 sg13g2_nand2_1 _2175_ (.Y(_1204_),
    .A(net726),
    .B(_1203_));
 sg13g2_nand2_1 _2176_ (.Y(_1205_),
    .A(net702),
    .B(net656));
 sg13g2_and4_1 _2177_ (.A(net704),
    .B(net681),
    .C(net679),
    .D(net656),
    .X(_1206_));
 sg13g2_a22oi_1 _2178_ (.Y(_1207_),
    .B1(net680),
    .B2(net678),
    .A2(net710),
    .A1(net694));
 sg13g2_nand2_1 _2179_ (.Y(_1208_),
    .A(net650),
    .B(_1016_));
 sg13g2_nand2_1 _2180_ (.Y(_1209_),
    .A(_1083_),
    .B(net625));
 sg13g2_a21o_1 _2181_ (.A2(net625),
    .A1(_1083_),
    .B1(net626),
    .X(_1210_));
 sg13g2_nand2_1 _2182_ (.Y(_1211_),
    .A(net761),
    .B(net626));
 sg13g2_nand2_2 _2183_ (.Y(_1212_),
    .A(net703),
    .B(_0982_));
 sg13g2_nor2_1 _2184_ (.A(net652),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_nand2_1 _2185_ (.Y(_1214_),
    .A(net708),
    .B(_1136_));
 sg13g2_nand3_1 _2186_ (.B(_1211_),
    .C(_1214_),
    .A(_1209_),
    .Y(_1215_));
 sg13g2_and2_1 _2187_ (.A(net735),
    .B(_1203_),
    .X(_1216_));
 sg13g2_nor2_1 _2188_ (.A(net747),
    .B(_1187_),
    .Y(_1217_));
 sg13g2_a22oi_1 _2189_ (.Y(_1218_),
    .B1(net689),
    .B2(net684),
    .A2(net712),
    .A1(net701));
 sg13g2_and4_1 _2190_ (.A(net681),
    .B(net679),
    .C(net755),
    .D(_1076_),
    .X(_1219_));
 sg13g2_nor2_1 _2191_ (.A(_1218_),
    .B(_1219_),
    .Y(_1220_));
 sg13g2_o21ai_1 _2192_ (.B1(_1189_),
    .Y(_1221_),
    .A1(net694),
    .A2(_0965_));
 sg13g2_and3_1 _2193_ (.X(_1222_),
    .A(_1024_),
    .B(_1220_),
    .C(_1221_));
 sg13g2_o21ai_1 _2194_ (.B1(net720),
    .Y(_1223_),
    .A1(_1217_),
    .A2(_1222_));
 sg13g2_and2_1 _2195_ (.A(net772),
    .B(net623),
    .X(_1224_));
 sg13g2_a21o_2 _2196_ (.A2(_1207_),
    .A1(_1205_),
    .B1(net626),
    .X(_1225_));
 sg13g2_mux2_1 _2197_ (.A0(_1210_),
    .A1(_1225_),
    .S(net768),
    .X(_1226_));
 sg13g2_nand2_1 _2198_ (.Y(_1227_),
    .A(_1076_),
    .B(net625));
 sg13g2_o21ai_1 _2199_ (.B1(_1187_),
    .Y(_1228_),
    .A1(net761),
    .A2(_1227_));
 sg13g2_nand2_1 _2200_ (.Y(_1229_),
    .A(net645),
    .B(_1083_));
 sg13g2_nand2_1 _2201_ (.Y(_1230_),
    .A(_1208_),
    .B(_1229_));
 sg13g2_o21ai_1 _2202_ (.B1(net734),
    .Y(_1231_),
    .A1(net625),
    .A2(_1218_));
 sg13g2_o21ai_1 _2203_ (.B1(net758),
    .Y(_1232_),
    .A1(_1171_),
    .A2(_1172_));
 sg13g2_o21ai_1 _2204_ (.B1(_1231_),
    .Y(_1233_),
    .A1(net770),
    .A2(_1232_));
 sg13g2_o21ai_1 _2205_ (.B1(net660),
    .Y(_1234_),
    .A1(_1230_),
    .A2(_1233_));
 sg13g2_nor2_1 _2206_ (.A(net753),
    .B(_1163_),
    .Y(_1235_));
 sg13g2_nand4_1 _2207_ (.B(net682),
    .C(net762),
    .A(net687),
    .Y(_1236_),
    .D(net677));
 sg13g2_nand2_1 _2208_ (.Y(_1237_),
    .A(_1085_),
    .B(_1169_));
 sg13g2_o21ai_1 _2209_ (.B1(_1169_),
    .Y(_1238_),
    .A1(net770),
    .A2(_1085_));
 sg13g2_o21ai_1 _2210_ (.B1(net672),
    .Y(_1239_),
    .A1(_1235_),
    .A2(_1238_));
 sg13g2_nor2_1 _2211_ (.A(net637),
    .B(_1149_),
    .Y(_1240_));
 sg13g2_nand2b_1 _2212_ (.Y(_1241_),
    .B(_1150_),
    .A_N(net637));
 sg13g2_o21ai_1 _2213_ (.B1(_1241_),
    .Y(_1242_),
    .A1(net770),
    .A2(_1169_));
 sg13g2_o21ai_1 _2214_ (.B1(_1124_),
    .Y(_1243_),
    .A1(net649),
    .A2(_1032_));
 sg13g2_a21oi_2 _2215_ (.B1(net664),
    .Y(_1244_),
    .A2(_1210_),
    .A1(net720));
 sg13g2_a22oi_1 _2216_ (.Y(_1245_),
    .B1(_1204_),
    .B2(_1244_),
    .A2(net669),
    .A1(net744));
 sg13g2_o21ai_1 _2217_ (.B1(net706),
    .Y(_1246_),
    .A1(_1079_),
    .A2(_1216_));
 sg13g2_and2_1 _2218_ (.A(net768),
    .B(net623),
    .X(_1247_));
 sg13g2_o21ai_1 _2219_ (.B1(net673),
    .Y(_1248_),
    .A1(_1215_),
    .A2(_1247_));
 sg13g2_nand3b_1 _2220_ (.B(_1246_),
    .C(_1248_),
    .Y(_1249_),
    .A_N(_1245_));
 sg13g2_a22oi_1 _2221_ (.Y(_1250_),
    .B1(_1226_),
    .B2(net706),
    .A2(_1225_),
    .A1(net674));
 sg13g2_a21oi_1 _2222_ (.A1(_1066_),
    .A2(_1228_),
    .Y(_1251_),
    .B1(net669));
 sg13g2_nand3_1 _2223_ (.B(_1250_),
    .C(_1251_),
    .A(_1223_),
    .Y(_1252_));
 sg13g2_a21oi_1 _2224_ (.A1(_1249_),
    .A2(_1252_),
    .Y(_1253_),
    .B1(net636));
 sg13g2_a22oi_1 _2225_ (.Y(_1254_),
    .B1(net622),
    .B2(net705),
    .A2(_1242_),
    .A1(net674));
 sg13g2_nand3_1 _2226_ (.B(_1239_),
    .C(_1254_),
    .A(_1234_),
    .Y(_1255_));
 sg13g2_o21ai_1 _2227_ (.B1(_1189_),
    .Y(_1256_),
    .A1(net753),
    .A2(net638));
 sg13g2_a221oi_1 _2228_ (.B2(net764),
    .C1(_1191_),
    .B1(_1256_),
    .A1(net740),
    .Y(_1257_),
    .A2(_1192_));
 sg13g2_nor2_1 _2229_ (.A(net662),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_a221oi_1 _2230_ (.B2(_1202_),
    .C1(net633),
    .B1(_1258_),
    .A1(net662),
    .Y(_1259_),
    .A2(_1255_));
 sg13g2_o21ai_1 _2231_ (.B1(_1103_),
    .Y(_1260_),
    .A1(_1253_),
    .A2(_1259_));
 sg13g2_nand3_1 _2232_ (.B(_1185_),
    .C(_1260_),
    .A(_1183_),
    .Y(_1261_));
 sg13g2_xor2_1 _2233_ (.B(_0938_),
    .A(_0937_),
    .X(_1262_));
 sg13g2_xnor2_1 _2234_ (.Y(_1263_),
    .A(_0937_),
    .B(_0938_));
 sg13g2_o21ai_1 _2235_ (.B1(_1173_),
    .Y(_1264_),
    .A1(_1044_),
    .A2(_1170_));
 sg13g2_nand3_1 _2236_ (.B(_1138_),
    .C(_1166_),
    .A(net752),
    .Y(_1265_));
 sg13g2_a21oi_1 _2237_ (.A1(_1138_),
    .A2(_1158_),
    .Y(_1266_),
    .B1(net717));
 sg13g2_nand2_1 _2238_ (.Y(_1267_),
    .A(_1265_),
    .B(_1266_));
 sg13g2_o21ai_1 _2239_ (.B1(_1021_),
    .Y(_1268_),
    .A1(_1264_),
    .A2(_1267_));
 sg13g2_nor2_1 _2240_ (.A(net761),
    .B(_1003_),
    .Y(_1269_));
 sg13g2_nor3_1 _2241_ (.A(_1159_),
    .B(_1179_),
    .C(_1269_),
    .Y(_1270_));
 sg13g2_nand2_1 _2242_ (.Y(_1271_),
    .A(net755),
    .B(_1151_));
 sg13g2_a21oi_1 _2243_ (.A1(net761),
    .A2(_1176_),
    .Y(_1272_),
    .B1(_1065_));
 sg13g2_nand2_1 _2244_ (.Y(_1273_),
    .A(_1271_),
    .B(_1272_));
 sg13g2_a21o_1 _2245_ (.A2(_1150_),
    .A1(_1092_),
    .B1(_1179_),
    .X(_1274_));
 sg13g2_a221oi_1 _2246_ (.B2(net707),
    .C1(net725),
    .B1(_1274_),
    .A1(_1271_),
    .Y(_1275_),
    .A2(_1272_));
 sg13g2_a21o_1 _2247_ (.A2(_1270_),
    .A1(_1268_),
    .B1(_1275_),
    .X(_1276_));
 sg13g2_a21oi_1 _2248_ (.A1(net650),
    .A2(_1110_),
    .Y(_1277_),
    .B1(net764));
 sg13g2_a221oi_1 _2249_ (.B2(net652),
    .C1(net765),
    .B1(_1110_),
    .A1(_0983_),
    .Y(_1278_),
    .A2(_1017_));
 sg13g2_nand2_1 _2250_ (.Y(_1279_),
    .A(net646),
    .B(_1121_));
 sg13g2_mux2_1 _2251_ (.A0(net713),
    .A1(net691),
    .S(net694),
    .X(_1280_));
 sg13g2_mux2_1 _2252_ (.A0(_1121_),
    .A1(_1280_),
    .S(net651),
    .X(_1281_));
 sg13g2_a22oi_1 _2253_ (.Y(_1282_),
    .B1(_1281_),
    .B2(net732),
    .A2(_1278_),
    .A1(net759));
 sg13g2_nor2_2 _2254_ (.A(net648),
    .B(net638),
    .Y(_1283_));
 sg13g2_o21ai_1 _2255_ (.B1(_1105_),
    .Y(_1284_),
    .A1(_1120_),
    .A2(_1283_));
 sg13g2_a21o_1 _2256_ (.A2(_1284_),
    .A1(_1282_),
    .B1(net670),
    .X(_1285_));
 sg13g2_nor2_2 _2257_ (.A(net723),
    .B(_1133_),
    .Y(_1286_));
 sg13g2_nand2_2 _2258_ (.Y(_1287_),
    .A(net717),
    .B(_1132_));
 sg13g2_a21oi_1 _2259_ (.A1(net648),
    .A2(_1109_),
    .Y(_1288_),
    .B1(_0996_));
 sg13g2_or2_1 _2260_ (.X(_1289_),
    .B(_1288_),
    .A(net759));
 sg13g2_a21o_1 _2261_ (.A2(net629),
    .A1(net639),
    .B1(net643),
    .X(_1290_));
 sg13g2_nand2_2 _2262_ (.Y(_1291_),
    .A(net761),
    .B(_1290_));
 sg13g2_o21ai_1 _2263_ (.B1(_1031_),
    .Y(_1292_),
    .A1(_1136_),
    .A2(_1142_));
 sg13g2_nor2_1 _2264_ (.A(net728),
    .B(_1159_),
    .Y(_1293_));
 sg13g2_mux2_1 _2265_ (.A0(_1130_),
    .A1(_1176_),
    .S(net752),
    .X(_1294_));
 sg13g2_nor2_2 _2266_ (.A(net719),
    .B(_1025_),
    .Y(_1295_));
 sg13g2_nand2_1 _2267_ (.Y(_1296_),
    .A(net723),
    .B(net707));
 sg13g2_nand2b_1 _2268_ (.Y(_1297_),
    .B(net655),
    .A_N(_1294_));
 sg13g2_nor2_1 _2269_ (.A(_1288_),
    .B(_1293_),
    .Y(_1298_));
 sg13g2_a21oi_1 _2270_ (.A1(_1289_),
    .A2(_1291_),
    .Y(_1299_),
    .B1(net774));
 sg13g2_o21ai_1 _2271_ (.B1(net661),
    .Y(_1300_),
    .A1(_1298_),
    .A2(_1299_));
 sg13g2_and4_1 _2272_ (.A(_1146_),
    .B(_1285_),
    .C(_1292_),
    .D(_1297_),
    .X(_1301_));
 sg13g2_a221oi_1 _2273_ (.B2(_1301_),
    .C1(net635),
    .B1(_1300_),
    .A1(_1178_),
    .Y(_1302_),
    .A2(_1276_));
 sg13g2_nor2_1 _2274_ (.A(net742),
    .B(_1290_),
    .Y(_1303_));
 sg13g2_a22oi_1 _2275_ (.Y(_1304_),
    .B1(net656),
    .B2(net696),
    .A2(net682),
    .A1(net688));
 sg13g2_a21oi_2 _2276_ (.B1(net624),
    .Y(_1305_),
    .A2(net756),
    .A1(net643));
 sg13g2_and3_1 _2277_ (.X(_1306_),
    .A(_1011_),
    .B(_1045_),
    .C(_1305_));
 sg13g2_a221oi_1 _2278_ (.B2(net742),
    .C1(net719),
    .B1(_1306_),
    .A1(_1013_),
    .Y(_1307_),
    .A2(_1303_));
 sg13g2_nand3_1 _2279_ (.B(net756),
    .C(_1012_),
    .A(net773),
    .Y(_1308_));
 sg13g2_a221oi_1 _2280_ (.B2(_1308_),
    .C1(net671),
    .B1(_1037_),
    .A1(net733),
    .Y(_1309_),
    .A2(_1035_));
 sg13g2_nand2_2 _2281_ (.Y(_1310_),
    .A(net735),
    .B(_1206_));
 sg13g2_a22oi_1 _2282_ (.Y(_1311_),
    .B1(_1310_),
    .B2(_1036_),
    .A2(_1056_),
    .A1(net729));
 sg13g2_o21ai_1 _2283_ (.B1(net669),
    .Y(_1312_),
    .A1(net658),
    .A2(_1311_));
 sg13g2_nor3_1 _2284_ (.A(net760),
    .B(net658),
    .C(_1055_),
    .Y(_1313_));
 sg13g2_or4_1 _2285_ (.A(_1307_),
    .B(_1309_),
    .C(_1312_),
    .D(_1313_),
    .X(_1314_));
 sg13g2_mux2_1 _2286_ (.A0(_0960_),
    .A1(_1076_),
    .S(net697),
    .X(_1315_));
 sg13g2_mux2_1 _2287_ (.A0(net709),
    .A1(net656),
    .S(net697),
    .X(_1316_));
 sg13g2_nand2b_1 _2288_ (.Y(_1317_),
    .B(_1316_),
    .A_N(net631));
 sg13g2_nor3_1 _2289_ (.A(net631),
    .B(_1106_),
    .C(_1315_),
    .Y(_1318_));
 sg13g2_a221oi_1 _2290_ (.B2(_1078_),
    .C1(net730),
    .B1(_1077_),
    .A1(net647),
    .Y(_1319_),
    .A2(_1067_));
 sg13g2_a221oi_1 _2291_ (.B2(_0924_),
    .C1(_0982_),
    .B1(_0989_),
    .A1(net704),
    .Y(_1320_),
    .A2(net709));
 sg13g2_a221oi_1 _2292_ (.B2(net762),
    .C1(_1320_),
    .B1(_1315_),
    .A1(net647),
    .Y(_1321_),
    .A2(_1067_));
 sg13g2_a221oi_1 _2293_ (.B2(net775),
    .C1(_1318_),
    .B1(_1321_),
    .A1(net733),
    .Y(_1322_),
    .A2(_1079_));
 sg13g2_nand2b_1 _2294_ (.Y(_1323_),
    .B(net673),
    .A_N(_1322_));
 sg13g2_nor2_1 _2295_ (.A(_1035_),
    .B(net626),
    .Y(_1324_));
 sg13g2_nor3_1 _2296_ (.A(_1030_),
    .B(_1035_),
    .C(net626),
    .Y(_1325_));
 sg13g2_o21ai_1 _2297_ (.B1(net725),
    .Y(_1326_),
    .A1(_1088_),
    .A2(_1325_));
 sg13g2_nor2_2 _2298_ (.A(net717),
    .B(_1133_),
    .Y(_1327_));
 sg13g2_nand2_2 _2299_ (.Y(_1328_),
    .A(net725),
    .B(_1132_));
 sg13g2_a21o_1 _2300_ (.A2(_1067_),
    .A1(_0983_),
    .B1(net647),
    .X(_1329_));
 sg13g2_o21ai_1 _2301_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_1092_),
    .A2(_1093_));
 sg13g2_nand2_1 _2302_ (.Y(_1331_),
    .A(_1327_),
    .B(_1330_));
 sg13g2_a221oi_1 _2303_ (.B2(_1049_),
    .C1(net668),
    .B1(_1087_),
    .A1(_1051_),
    .Y(_1332_),
    .A2(_1079_));
 sg13g2_nand4_1 _2304_ (.B(_1326_),
    .C(_1331_),
    .A(_1323_),
    .Y(_1333_),
    .D(_1332_));
 sg13g2_nand3_1 _2305_ (.B(_1314_),
    .C(_1333_),
    .A(net636),
    .Y(_1334_));
 sg13g2_nand3b_1 _2306_ (.B(_1334_),
    .C(net618),
    .Y(_1335_),
    .A_N(_1302_));
 sg13g2_nand2_2 _2307_ (.Y(_1336_),
    .A(net740),
    .B(net734));
 sg13g2_o21ai_1 _2308_ (.B1(net661),
    .Y(_1337_),
    .A1(_1233_),
    .A2(_1237_));
 sg13g2_a21oi_1 _2309_ (.A1(_1084_),
    .A2(_1336_),
    .Y(_1338_),
    .B1(_1169_));
 sg13g2_nor2_1 _2310_ (.A(net666),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_nand3_1 _2311_ (.B(_1337_),
    .C(_1339_),
    .A(_1239_),
    .Y(_1340_));
 sg13g2_a21o_1 _2312_ (.A2(_1243_),
    .A1(net758),
    .B1(_1196_),
    .X(_1341_));
 sg13g2_nor3_1 _2313_ (.A(_0934_),
    .B(_1188_),
    .C(_1190_),
    .Y(_1342_));
 sg13g2_nor2_2 _2314_ (.A(net722),
    .B(_1065_),
    .Y(_1343_));
 sg13g2_nand2_1 _2315_ (.Y(_1344_),
    .A(net723),
    .B(_1064_));
 sg13g2_o21ai_1 _2316_ (.B1(net666),
    .Y(_1345_),
    .A1(_1189_),
    .A2(_1344_));
 sg13g2_nor3_1 _2317_ (.A(net723),
    .B(_1132_),
    .C(_1194_),
    .Y(_1346_));
 sg13g2_a21oi_1 _2318_ (.A1(_1195_),
    .A2(_1327_),
    .Y(_1347_),
    .B1(_1345_));
 sg13g2_a221oi_1 _2319_ (.B2(_1341_),
    .C1(_1346_),
    .B1(_1286_),
    .A1(_1049_),
    .Y(_1348_),
    .A2(_1256_));
 sg13g2_nand3b_1 _2320_ (.B(_1347_),
    .C(_1348_),
    .Y(_1349_),
    .A_N(_1342_));
 sg13g2_nand3_1 _2321_ (.B(_1340_),
    .C(_1349_),
    .A(net634),
    .Y(_1350_));
 sg13g2_nand2_2 _2322_ (.Y(_1351_),
    .A(_1186_),
    .B(_1227_));
 sg13g2_a221oi_1 _2323_ (.B2(net718),
    .C1(net667),
    .B1(_1351_),
    .A1(net706),
    .Y(_1352_),
    .A2(net623));
 sg13g2_nand3_1 _2324_ (.B(_1220_),
    .C(_1221_),
    .A(net768),
    .Y(_1353_));
 sg13g2_a22oi_1 _2325_ (.Y(_1354_),
    .B1(_1225_),
    .B2(net729),
    .A2(net623),
    .A1(net774));
 sg13g2_a21o_1 _2326_ (.A2(_1354_),
    .A1(_1353_),
    .B1(_1021_),
    .X(_1355_));
 sg13g2_nor2_2 _2327_ (.A(net717),
    .B(_1132_),
    .Y(_1356_));
 sg13g2_a22oi_1 _2328_ (.Y(_1357_),
    .B1(_1356_),
    .B2(_1079_),
    .A2(_1327_),
    .A1(_1215_));
 sg13g2_a221oi_1 _2329_ (.B2(_1244_),
    .C1(net634),
    .B1(_1357_),
    .A1(_1352_),
    .Y(_1358_),
    .A2(_1355_));
 sg13g2_nor2_1 _2330_ (.A(net619),
    .B(_1358_),
    .Y(_1359_));
 sg13g2_a21oi_1 _2331_ (.A1(_1350_),
    .A2(_1359_),
    .Y(_1360_),
    .B1(_1185_));
 sg13g2_a21oi_1 _2332_ (.A1(_1335_),
    .A2(_1360_),
    .Y(_1361_),
    .B1(_1262_));
 sg13g2_o21ai_1 _2333_ (.B1(net740),
    .Y(_1362_),
    .A1(_1198_),
    .A2(_1277_));
 sg13g2_a221oi_1 _2334_ (.B2(_1064_),
    .C1(net724),
    .B1(_1195_),
    .A1(net707),
    .Y(_1363_),
    .A2(_1192_));
 sg13g2_a21o_1 _2335_ (.A2(_1363_),
    .A1(_1362_),
    .B1(_1193_),
    .X(_1364_));
 sg13g2_nor2_1 _2336_ (.A(_1172_),
    .B(_1218_),
    .Y(_1365_));
 sg13g2_nand3_1 _2337_ (.B(_1232_),
    .C(_1365_),
    .A(net763),
    .Y(_1366_));
 sg13g2_nand3_1 _2338_ (.B(_1208_),
    .C(_1229_),
    .A(net770),
    .Y(_1367_));
 sg13g2_nand3_1 _2339_ (.B(_1366_),
    .C(_1367_),
    .A(net661),
    .Y(_1368_));
 sg13g2_nor2_1 _2340_ (.A(net731),
    .B(_1168_),
    .Y(_1369_));
 sg13g2_or2_1 _2341_ (.X(_1370_),
    .B(_1369_),
    .A(_1240_));
 sg13g2_nor2_1 _2342_ (.A(net753),
    .B(_1229_),
    .Y(_1371_));
 sg13g2_nand3_1 _2343_ (.B(net732),
    .C(_1083_),
    .A(net645),
    .Y(_1372_));
 sg13g2_a21oi_1 _2344_ (.A1(net650),
    .A2(_1032_),
    .Y(_1373_),
    .B1(_1167_));
 sg13g2_a21oi_1 _2345_ (.A1(_1372_),
    .A2(_1373_),
    .Y(_1374_),
    .B1(net670));
 sg13g2_a21oi_1 _2346_ (.A1(net770),
    .A2(_1142_),
    .Y(_1375_),
    .B1(net666));
 sg13g2_a21oi_1 _2347_ (.A1(net740),
    .A2(_1370_),
    .Y(_1376_),
    .B1(_1374_));
 sg13g2_and3_1 _2348_ (.X(_1377_),
    .A(_1368_),
    .B(_1375_),
    .C(_1376_));
 sg13g2_nand2_1 _2349_ (.Y(_1378_),
    .A(net764),
    .B(_1240_));
 sg13g2_a22oi_1 _2350_ (.Y(_1379_),
    .B1(net622),
    .B2(net734),
    .A2(_1240_),
    .A1(net732));
 sg13g2_a22oi_1 _2351_ (.Y(_1380_),
    .B1(_1377_),
    .B2(_1379_),
    .A2(_1364_),
    .A1(net666));
 sg13g2_or3_1 _2352_ (.A(_1189_),
    .B(_1218_),
    .C(_1219_),
    .X(_1381_));
 sg13g2_nor2_1 _2353_ (.A(_1065_),
    .B(_1381_),
    .Y(_1382_));
 sg13g2_o21ai_1 _2354_ (.B1(net720),
    .Y(_1383_),
    .A1(_1217_),
    .A2(_1382_));
 sg13g2_o21ai_1 _2355_ (.B1(_0995_),
    .Y(_1384_),
    .A1(net639),
    .A2(net626));
 sg13g2_nand2_1 _2356_ (.Y(_1385_),
    .A(net720),
    .B(_1025_));
 sg13g2_a21oi_1 _2357_ (.A1(_1027_),
    .A2(_1328_),
    .Y(_1386_),
    .B1(_1384_));
 sg13g2_a21oi_1 _2358_ (.A1(_1225_),
    .A2(_1356_),
    .Y(_1387_),
    .B1(_1386_));
 sg13g2_nand3_1 _2359_ (.B(_1383_),
    .C(_1387_),
    .A(net664),
    .Y(_1388_));
 sg13g2_nand2_1 _2360_ (.Y(_1389_),
    .A(net661),
    .B(_1226_));
 sg13g2_a221oi_1 _2361_ (.B2(_1203_),
    .C1(net664),
    .B1(_1385_),
    .A1(_1066_),
    .Y(_1390_),
    .A2(_1215_));
 sg13g2_a21oi_1 _2362_ (.A1(_1389_),
    .A2(_1390_),
    .Y(_1391_),
    .B1(net636));
 sg13g2_a221oi_1 _2363_ (.B2(_1391_),
    .C1(net619),
    .B1(_1388_),
    .A1(net636),
    .Y(_1392_),
    .A2(_1380_));
 sg13g2_nand2b_1 _2364_ (.Y(_1393_),
    .B(_1150_),
    .A_N(_1115_));
 sg13g2_nand3b_1 _2365_ (.B(_1150_),
    .C(net728),
    .Y(_1394_),
    .A_N(_1115_));
 sg13g2_o21ai_1 _2366_ (.B1(net737),
    .Y(_1395_),
    .A1(_1107_),
    .A2(_1160_));
 sg13g2_a221oi_1 _2367_ (.B2(net737),
    .C1(_1107_),
    .B1(_1160_),
    .A1(net675),
    .Y(_1396_),
    .A2(net631));
 sg13g2_a21oi_1 _2368_ (.A1(_1394_),
    .A2(_1396_),
    .Y(_1397_),
    .B1(net670));
 sg13g2_nor3_1 _2369_ (.A(net734),
    .B(net657),
    .C(_1155_),
    .Y(_1398_));
 sg13g2_nor3_1 _2370_ (.A(_1044_),
    .B(net657),
    .C(_1176_),
    .Y(_1399_));
 sg13g2_nor3_1 _2371_ (.A(_1397_),
    .B(_1398_),
    .C(_1399_),
    .Y(_1400_));
 sg13g2_a221oi_1 _2372_ (.B2(net738),
    .C1(net628),
    .B1(_1171_),
    .A1(net646),
    .Y(_1401_),
    .A2(_1119_));
 sg13g2_a21oi_1 _2373_ (.A1(_1163_),
    .A2(_1401_),
    .Y(_1402_),
    .B1(_1021_));
 sg13g2_o21ai_1 _2374_ (.B1(net655),
    .Y(_1403_),
    .A1(_1171_),
    .A2(_1172_));
 sg13g2_nand2_1 _2375_ (.Y(_1404_),
    .A(net667),
    .B(_1403_));
 sg13g2_nor2_1 _2376_ (.A(_0934_),
    .B(_1170_),
    .Y(_1405_));
 sg13g2_nor3_1 _2377_ (.A(_1402_),
    .B(_1404_),
    .C(_1405_),
    .Y(_1406_));
 sg13g2_nand2b_1 _2378_ (.Y(_1407_),
    .B(_1286_),
    .A_N(_1294_));
 sg13g2_nand3_1 _2379_ (.B(_1406_),
    .C(_1407_),
    .A(_1400_),
    .Y(_1408_));
 sg13g2_and2_1 _2380_ (.A(net660),
    .B(_1113_),
    .X(_1409_));
 sg13g2_a21o_1 _2381_ (.A2(_1121_),
    .A1(net645),
    .B1(net628),
    .X(_1410_));
 sg13g2_a22oi_1 _2382_ (.Y(_1411_),
    .B1(_1410_),
    .B2(net737),
    .A2(_1111_),
    .A1(net728));
 sg13g2_nor2_1 _2383_ (.A(net657),
    .B(_1411_),
    .Y(_1412_));
 sg13g2_a21oi_1 _2384_ (.A1(net763),
    .A2(_1410_),
    .Y(_1413_),
    .B1(net728));
 sg13g2_a221oi_1 _2385_ (.B2(net732),
    .C1(net649),
    .B1(_1121_),
    .A1(_1004_),
    .Y(_1414_),
    .A2(net629));
 sg13g2_nand3b_1 _2386_ (.B(net672),
    .C(_1150_),
    .Y(_1415_),
    .A_N(_1414_));
 sg13g2_a221oi_1 _2387_ (.B2(net683),
    .C1(_0962_),
    .B1(net687),
    .A1(net696),
    .Y(_1416_),
    .A2(net714));
 sg13g2_nand2_1 _2388_ (.Y(_1417_),
    .A(_0968_),
    .B(net630));
 sg13g2_a21o_1 _2389_ (.A2(net630),
    .A1(_0968_),
    .B1(net628),
    .X(_1418_));
 sg13g2_a21oi_1 _2390_ (.A1(_1031_),
    .A2(_1418_),
    .Y(_1419_),
    .B1(net667));
 sg13g2_o21ai_1 _2391_ (.B1(_1419_),
    .Y(_1420_),
    .A1(_1413_),
    .A2(_1415_));
 sg13g2_a21oi_1 _2392_ (.A1(net752),
    .A2(_1131_),
    .Y(_1421_),
    .B1(net627));
 sg13g2_a221oi_1 _2393_ (.B2(net752),
    .C1(net627),
    .B1(_1131_),
    .A1(_0968_),
    .Y(_1422_),
    .A2(net630));
 sg13g2_a21oi_1 _2394_ (.A1(_1134_),
    .A2(_1422_),
    .Y(_1423_),
    .B1(net717));
 sg13g2_or4_1 _2395_ (.A(_1409_),
    .B(_1412_),
    .C(_1420_),
    .D(_1423_),
    .X(_1424_));
 sg13g2_a21oi_1 _2396_ (.A1(_1408_),
    .A2(_1424_),
    .Y(_1425_),
    .B1(net635));
 sg13g2_nand2_1 _2397_ (.Y(_1426_),
    .A(net725),
    .B(_1019_));
 sg13g2_nand2_1 _2398_ (.Y(_1427_),
    .A(_0934_),
    .B(_1426_));
 sg13g2_o21ai_1 _2399_ (.B1(_1427_),
    .Y(_1428_),
    .A1(net742),
    .A2(_1014_));
 sg13g2_nand2_2 _2400_ (.Y(_1429_),
    .A(net745),
    .B(net730));
 sg13g2_nor3_1 _2401_ (.A(net641),
    .B(_0996_),
    .C(_1017_),
    .Y(_1430_));
 sg13g2_o21ai_1 _2402_ (.B1(net719),
    .Y(_1431_),
    .A1(_1429_),
    .A2(_1430_));
 sg13g2_a22oi_1 _2403_ (.Y(_1432_),
    .B1(net735),
    .B2(net743),
    .A2(net653),
    .A1(_0968_));
 sg13g2_a21oi_1 _2404_ (.A1(net648),
    .A2(_1054_),
    .Y(_1433_),
    .B1(_1336_));
 sg13g2_a22oi_1 _2405_ (.Y(_1434_),
    .B1(_1433_),
    .B2(_0997_),
    .A2(_1432_),
    .A1(_1034_));
 sg13g2_nor2_1 _2406_ (.A(_1431_),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_nor2_1 _2407_ (.A(net664),
    .B(_1435_),
    .Y(_1436_));
 sg13g2_nor2_2 _2408_ (.A(net718),
    .B(net707),
    .Y(_1437_));
 sg13g2_nand2_1 _2409_ (.Y(_1438_),
    .A(_0967_),
    .B(net637));
 sg13g2_o21ai_1 _2410_ (.B1(_1437_),
    .Y(_1439_),
    .A1(_1028_),
    .A2(_1438_));
 sg13g2_a22oi_1 _2411_ (.Y(_1440_),
    .B1(_1439_),
    .B2(_1027_),
    .A2(_1087_),
    .A1(_0967_));
 sg13g2_nor3_1 _2412_ (.A(net658),
    .B(_1072_),
    .C(_1216_),
    .Y(_1441_));
 sg13g2_o21ai_1 _2413_ (.B1(_1212_),
    .Y(_1442_),
    .A1(net641),
    .A2(_0996_));
 sg13g2_nand3_1 _2414_ (.B(_1438_),
    .C(_1442_),
    .A(net655),
    .Y(_1443_));
 sg13g2_a21o_1 _2415_ (.A2(_1161_),
    .A1(net708),
    .B1(_1443_),
    .X(_1444_));
 sg13g2_nor3_1 _2416_ (.A(net773),
    .B(net671),
    .C(_1094_),
    .Y(_1445_));
 sg13g2_nor4_1 _2417_ (.A(net668),
    .B(_1440_),
    .C(_1441_),
    .D(_1445_),
    .Y(_1446_));
 sg13g2_a221oi_1 _2418_ (.B2(_1446_),
    .C1(_1063_),
    .B1(_1444_),
    .A1(_1428_),
    .Y(_1447_),
    .A2(_1436_));
 sg13g2_o21ai_1 _2419_ (.B1(net618),
    .Y(_1448_),
    .A1(_1425_),
    .A2(_1447_));
 sg13g2_nand3b_1 _2420_ (.B(_1448_),
    .C(_1184_),
    .Y(_1449_),
    .A_N(_1392_));
 sg13g2_nor2_1 _2421_ (.A(_1065_),
    .B(_1430_),
    .Y(_1450_));
 sg13g2_a221oi_1 _2422_ (.B2(_0934_),
    .C1(_1450_),
    .B1(_1426_),
    .A1(_0986_),
    .Y(_1451_),
    .A2(net707));
 sg13g2_nor3_1 _2423_ (.A(net745),
    .B(net731),
    .C(_1166_),
    .Y(_1452_));
 sg13g2_nand3_1 _2424_ (.B(net652),
    .C(_1076_),
    .A(_0959_),
    .Y(_1453_));
 sg13g2_a22oi_1 _2425_ (.Y(_1454_),
    .B1(_1433_),
    .B2(_1453_),
    .A2(_1432_),
    .A1(_1018_));
 sg13g2_nor3_1 _2426_ (.A(_1431_),
    .B(_1452_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_o21ai_1 _2427_ (.B1(net668),
    .Y(_1456_),
    .A1(_1451_),
    .A2(_1455_));
 sg13g2_nand4_1 _2428_ (.B(net730),
    .C(_1438_),
    .A(net745),
    .Y(_1457_),
    .D(_1442_));
 sg13g2_a22oi_1 _2429_ (.Y(_1458_),
    .B1(_1084_),
    .B2(net647),
    .A2(net730),
    .A1(net745));
 sg13g2_a21oi_1 _2430_ (.A1(_1442_),
    .A2(_1458_),
    .Y(_1459_),
    .B1(net719));
 sg13g2_nor3_1 _2431_ (.A(_1092_),
    .B(_1093_),
    .C(_1105_),
    .Y(_1460_));
 sg13g2_nor2_1 _2432_ (.A(net774),
    .B(_1161_),
    .Y(_1461_));
 sg13g2_nand2_1 _2433_ (.Y(_1462_),
    .A(_0995_),
    .B(_1150_));
 sg13g2_a221oi_1 _2434_ (.B2(_1070_),
    .C1(_1460_),
    .B1(_1462_),
    .A1(_1203_),
    .Y(_1463_),
    .A2(_1461_));
 sg13g2_nor3_1 _2435_ (.A(_0962_),
    .B(_0966_),
    .C(_1139_),
    .Y(_1464_));
 sg13g2_a221oi_1 _2436_ (.B2(net673),
    .C1(net668),
    .B1(_1464_),
    .A1(_1457_),
    .Y(_1465_),
    .A2(_1459_));
 sg13g2_o21ai_1 _2437_ (.B1(_1465_),
    .Y(_1466_),
    .A1(net658),
    .A2(_1463_));
 sg13g2_nand3_1 _2438_ (.B(_1456_),
    .C(_1466_),
    .A(net636),
    .Y(_1467_));
 sg13g2_o21ai_1 _2439_ (.B1(_1108_),
    .Y(_1468_),
    .A1(net649),
    .A2(_1128_));
 sg13g2_nand3_1 _2440_ (.B(_1429_),
    .C(_1468_),
    .A(_1356_),
    .Y(_1469_));
 sg13g2_nand3_1 _2441_ (.B(net731),
    .C(_1131_),
    .A(net705),
    .Y(_1470_));
 sg13g2_nand2_1 _2442_ (.Y(_1471_),
    .A(_1469_),
    .B(_1470_));
 sg13g2_nor2_1 _2443_ (.A(net757),
    .B(_1009_),
    .Y(_1472_));
 sg13g2_o21ai_1 _2444_ (.B1(_1327_),
    .Y(_1473_),
    .A1(_1418_),
    .A2(_1472_));
 sg13g2_a21o_1 _2445_ (.A2(_1109_),
    .A1(net649),
    .B1(net644),
    .X(_1474_));
 sg13g2_nand2_1 _2446_ (.Y(_1475_),
    .A(net757),
    .B(_1474_));
 sg13g2_a21oi_1 _2447_ (.A1(net757),
    .A2(_1474_),
    .Y(_1476_),
    .B1(_1111_));
 sg13g2_o21ai_1 _2448_ (.B1(_1473_),
    .Y(_1477_),
    .A1(_1287_),
    .A2(_1476_));
 sg13g2_nor4_1 _2449_ (.A(_1412_),
    .B(_1420_),
    .C(_1471_),
    .D(_1477_),
    .Y(_1478_));
 sg13g2_nand4_1 _2450_ (.B(_0962_),
    .C(net680),
    .A(net700),
    .Y(_1479_),
    .D(net678));
 sg13g2_nand3_1 _2451_ (.B(_1140_),
    .C(_1479_),
    .A(_1124_),
    .Y(_1480_));
 sg13g2_nand2_2 _2452_ (.Y(_1481_),
    .A(net772),
    .B(net661));
 sg13g2_a21oi_1 _2453_ (.A1(net772),
    .A2(_1155_),
    .Y(_1482_),
    .B1(net657));
 sg13g2_o21ai_1 _2454_ (.B1(net769),
    .Y(_1483_),
    .A1(net752),
    .A2(_1130_));
 sg13g2_o21ai_1 _2455_ (.B1(_1482_),
    .Y(_1484_),
    .A1(_1480_),
    .A2(_1483_));
 sg13g2_a21oi_1 _2456_ (.A1(_1393_),
    .A2(_1395_),
    .Y(_1485_),
    .B1(net670));
 sg13g2_nor4_1 _2457_ (.A(_1402_),
    .B(_1404_),
    .C(_1405_),
    .D(_1485_),
    .Y(_1486_));
 sg13g2_a21oi_1 _2458_ (.A1(_1484_),
    .A2(_1486_),
    .Y(_1487_),
    .B1(net635));
 sg13g2_nand2b_1 _2459_ (.Y(_1488_),
    .B(_1487_),
    .A_N(_1478_));
 sg13g2_nand3_1 _2460_ (.B(_1467_),
    .C(_1488_),
    .A(net618),
    .Y(_1489_));
 sg13g2_o21ai_1 _2461_ (.B1(net660),
    .Y(_1490_),
    .A1(_1198_),
    .A2(_1277_));
 sg13g2_a21oi_1 _2462_ (.A1(_1030_),
    .A2(_1192_),
    .Y(_1491_),
    .B1(_1283_));
 sg13g2_a21o_1 _2463_ (.A2(_1491_),
    .A1(_1187_),
    .B1(net720),
    .X(_1492_));
 sg13g2_nor2_1 _2464_ (.A(net730),
    .B(_1212_),
    .Y(_1493_));
 sg13g2_o21ai_1 _2465_ (.B1(net673),
    .Y(_1494_),
    .A1(_1192_),
    .A2(_1493_));
 sg13g2_nand4_1 _2466_ (.B(_1490_),
    .C(_1492_),
    .A(net666),
    .Y(_1495_),
    .D(_1494_));
 sg13g2_nand4_1 _2467_ (.B(_1375_),
    .C(_1376_),
    .A(_1368_),
    .Y(_1496_),
    .D(_1378_));
 sg13g2_nand3_1 _2468_ (.B(_1495_),
    .C(_1496_),
    .A(net635),
    .Y(_1497_));
 sg13g2_nand2b_1 _2469_ (.Y(_1498_),
    .B(_1381_),
    .A_N(_1481_));
 sg13g2_a221oi_1 _2470_ (.B2(net659),
    .C1(_1295_),
    .B1(_1384_),
    .A1(_1187_),
    .Y(_1499_),
    .A2(_1286_));
 sg13g2_a22oi_1 _2471_ (.Y(_1500_),
    .B1(_1498_),
    .B2(_1499_),
    .A2(_1295_),
    .A1(_1225_));
 sg13g2_a21oi_1 _2472_ (.A1(_1205_),
    .A2(net625),
    .Y(_1501_),
    .B1(_1213_));
 sg13g2_a21o_1 _2473_ (.A2(_1501_),
    .A1(_1310_),
    .B1(net658),
    .X(_1502_));
 sg13g2_a21o_1 _2474_ (.A2(_1205_),
    .A1(_1172_),
    .B1(_1068_),
    .X(_1503_));
 sg13g2_a221oi_1 _2475_ (.B2(net673),
    .C1(net664),
    .B1(_1503_),
    .A1(net726),
    .Y(_1504_),
    .A2(_1203_));
 sg13g2_a221oi_1 _2476_ (.B2(_1504_),
    .C1(net636),
    .B1(_1502_),
    .A1(net664),
    .Y(_1505_),
    .A2(_1500_));
 sg13g2_nor2_1 _2477_ (.A(net618),
    .B(_1505_),
    .Y(_1506_));
 sg13g2_a21oi_1 _2478_ (.A1(_1497_),
    .A2(_1506_),
    .Y(_1507_),
    .B1(_1184_));
 sg13g2_a21oi_1 _2479_ (.A1(_1489_),
    .A2(_1507_),
    .Y(_1508_),
    .B1(_1263_));
 sg13g2_xnor2_1 _2480_ (.Y(_1509_),
    .A(_0939_),
    .B(_0944_));
 sg13g2_inv_1 _2481_ (.Y(_1510_),
    .A(_1509_));
 sg13g2_a221oi_1 _2482_ (.B2(_1508_),
    .C1(_1510_),
    .B1(_1449_),
    .A1(_1261_),
    .Y(_1511_),
    .A2(_1361_));
 sg13g2_nand2_1 _2483_ (.Y(_1512_),
    .A(net650),
    .B(_1084_));
 sg13g2_a22oi_1 _2484_ (.Y(_1513_),
    .B1(_1084_),
    .B2(net650),
    .A2(net629),
    .A1(net632));
 sg13g2_nand2_1 _2485_ (.Y(_1514_),
    .A(_1186_),
    .B(_1512_));
 sg13g2_o21ai_1 _2486_ (.B1(net724),
    .Y(_1515_),
    .A1(net747),
    .A2(_1513_));
 sg13g2_nand3_1 _2487_ (.B(net630),
    .C(net629),
    .A(net759),
    .Y(_1516_));
 sg13g2_nand3_1 _2488_ (.B(net645),
    .C(_1129_),
    .A(net715),
    .Y(_1517_));
 sg13g2_nand2_1 _2489_ (.Y(_0117_),
    .A(_1512_),
    .B(_1517_));
 sg13g2_nand3_1 _2490_ (.B(_1516_),
    .C(_1517_),
    .A(_1512_),
    .Y(_0118_));
 sg13g2_a21o_1 _2491_ (.A2(_0118_),
    .A1(net765),
    .B1(_1224_),
    .X(_0119_));
 sg13g2_a21oi_1 _2492_ (.A1(net747),
    .A2(_0119_),
    .Y(_0120_),
    .B1(_1515_));
 sg13g2_a221oi_1 _2493_ (.B2(net772),
    .C1(net724),
    .B1(_1514_),
    .A1(_1025_),
    .Y(_0121_),
    .A2(_1351_));
 sg13g2_o21ai_1 _2494_ (.B1(net663),
    .Y(_0122_),
    .A1(_0120_),
    .A2(_0121_));
 sg13g2_nand2_1 _2495_ (.Y(_0123_),
    .A(net638),
    .B(net625));
 sg13g2_nand2b_2 _2496_ (.Y(_0124_),
    .B(_0123_),
    .A_N(net626));
 sg13g2_nand2_1 _2497_ (.Y(_0125_),
    .A(net714),
    .B(_1069_));
 sg13g2_a221oi_1 _2498_ (.B2(_0125_),
    .C1(net744),
    .B1(_0124_),
    .A1(net735),
    .Y(_0126_),
    .A2(net623));
 sg13g2_nand3_1 _2499_ (.B(net638),
    .C(net625),
    .A(_0959_),
    .Y(_0127_));
 sg13g2_nand2_1 _2500_ (.Y(_0128_),
    .A(net755),
    .B(_1068_));
 sg13g2_nand3_1 _2501_ (.B(_0127_),
    .C(_0128_),
    .A(_1211_),
    .Y(_0129_));
 sg13g2_a21oi_1 _2502_ (.A1(net707),
    .A2(_1317_),
    .Y(_0130_),
    .B1(net720));
 sg13g2_o21ai_1 _2503_ (.B1(_0130_),
    .Y(_0131_),
    .A1(_1065_),
    .A2(_0129_));
 sg13g2_o21ai_1 _2504_ (.B1(_1244_),
    .Y(_0132_),
    .A1(_0126_),
    .A2(_0131_));
 sg13g2_and2_1 _2505_ (.A(net633),
    .B(_0132_),
    .X(_0133_));
 sg13g2_a221oi_1 _2506_ (.B2(net700),
    .C1(net691),
    .B1(net676),
    .A1(net680),
    .Y(_0134_),
    .A2(net678));
 sg13g2_a21oi_1 _2507_ (.A1(_0995_),
    .A2(_1150_),
    .Y(_0135_),
    .B1(net691));
 sg13g2_o21ai_1 _2508_ (.B1(_0134_),
    .Y(_0136_),
    .A1(net771),
    .A2(_0135_));
 sg13g2_a22oi_1 _2509_ (.Y(_0137_),
    .B1(_1351_),
    .B2(net738),
    .A2(_1221_),
    .A1(net728));
 sg13g2_o21ai_1 _2510_ (.B1(net757),
    .Y(_0138_),
    .A1(net642),
    .A2(_1241_));
 sg13g2_nor2_1 _2511_ (.A(net657),
    .B(_1194_),
    .Y(_0139_));
 sg13g2_a21oi_1 _2512_ (.A1(_0138_),
    .A2(_0139_),
    .Y(_0140_),
    .B1(net662));
 sg13g2_a21oi_1 _2513_ (.A1(net753),
    .A2(_0134_),
    .Y(_0141_),
    .B1(_1021_));
 sg13g2_o21ai_1 _2514_ (.B1(_0140_),
    .Y(_0142_),
    .A1(_1344_),
    .A2(_0134_));
 sg13g2_a221oi_1 _2515_ (.B2(_0141_),
    .C1(_1346_),
    .B1(_0136_),
    .A1(_1005_),
    .Y(_0143_),
    .A2(_1031_));
 sg13g2_o21ai_1 _2516_ (.B1(_0143_),
    .Y(_0144_),
    .A1(_0934_),
    .A2(_0137_));
 sg13g2_or2_1 _2517_ (.X(_0145_),
    .B(_0144_),
    .A(_0142_));
 sg13g2_a21o_1 _2518_ (.A2(_1032_),
    .A1(net650),
    .B1(_1218_),
    .X(_0146_));
 sg13g2_o21ai_1 _2519_ (.B1(net660),
    .Y(_0147_),
    .A1(_1233_),
    .A2(_0146_));
 sg13g2_o21ai_1 _2520_ (.B1(net672),
    .Y(_0148_),
    .A1(_1238_),
    .A2(_1371_));
 sg13g2_nor2_2 _2521_ (.A(net627),
    .B(_1167_),
    .Y(_0149_));
 sg13g2_o21ai_1 _2522_ (.B1(_0149_),
    .Y(_0150_),
    .A1(net770),
    .A2(_1169_));
 sg13g2_a22oi_1 _2523_ (.Y(_0151_),
    .B1(_0150_),
    .B2(net674),
    .A2(net622),
    .A1(net705));
 sg13g2_nand4_1 _2524_ (.B(_0147_),
    .C(_0148_),
    .A(net662),
    .Y(_0152_),
    .D(_0151_));
 sg13g2_and2_1 _2525_ (.A(net634),
    .B(_0152_),
    .X(_0153_));
 sg13g2_a221oi_1 _2526_ (.B2(_0153_),
    .C1(net618),
    .B1(_0145_),
    .A1(_0122_),
    .Y(_0154_),
    .A2(_0133_));
 sg13g2_or2_1 _2527_ (.X(_0155_),
    .B(net624),
    .A(_1006_));
 sg13g2_o21ai_1 _2528_ (.B1(net775),
    .Y(_0156_),
    .A1(net639),
    .A2(net624));
 sg13g2_nor2_1 _2529_ (.A(net767),
    .B(_1162_),
    .Y(_0157_));
 sg13g2_or2_1 _2530_ (.X(_0158_),
    .B(net624),
    .A(net641));
 sg13g2_a221oi_1 _2531_ (.B2(net766),
    .C1(net671),
    .B1(_0158_),
    .A1(_0155_),
    .Y(_0159_),
    .A2(_0157_));
 sg13g2_nand3_1 _2532_ (.B(_1305_),
    .C(_1343_),
    .A(_1007_),
    .Y(_0160_));
 sg13g2_nand2_1 _2533_ (.Y(_0161_),
    .A(_0967_),
    .B(_1166_));
 sg13g2_nand4_1 _2534_ (.B(_0985_),
    .C(_1166_),
    .A(_0967_),
    .Y(_0162_),
    .D(net655));
 sg13g2_nand3_1 _2535_ (.B(_0160_),
    .C(_0162_),
    .A(net636),
    .Y(_0163_));
 sg13g2_o21ai_1 _2536_ (.B1(net760),
    .Y(_0164_),
    .A1(net641),
    .A2(_1114_));
 sg13g2_o21ai_1 _2537_ (.B1(net756),
    .Y(_0165_),
    .A1(net641),
    .A2(net624));
 sg13g2_a21oi_1 _2538_ (.A1(_0164_),
    .A2(_0165_),
    .Y(_0166_),
    .B1(net766));
 sg13g2_nor3_1 _2539_ (.A(net659),
    .B(_1324_),
    .C(_0166_),
    .Y(_0167_));
 sg13g2_nor2b_1 _2540_ (.A(_1008_),
    .B_N(_1161_),
    .Y(_0168_));
 sg13g2_o21ai_1 _2541_ (.B1(_1236_),
    .Y(_0169_),
    .A1(net639),
    .A2(_1304_));
 sg13g2_o21ai_1 _2542_ (.B1(_0156_),
    .Y(_0170_),
    .A1(_0168_),
    .A2(_0169_));
 sg13g2_nor2_1 _2543_ (.A(_1021_),
    .B(_0170_),
    .Y(_0171_));
 sg13g2_nor4_2 _2544_ (.A(_0159_),
    .B(_0163_),
    .C(_0167_),
    .Y(_0172_),
    .D(_0171_));
 sg13g2_o21ai_1 _2545_ (.B1(net728),
    .Y(_0173_),
    .A1(net652),
    .A2(_1212_));
 sg13g2_o21ai_1 _2546_ (.B1(_0173_),
    .Y(_0174_),
    .A1(net735),
    .A2(_1136_));
 sg13g2_nor2_1 _2547_ (.A(_1149_),
    .B(_1213_),
    .Y(_0175_));
 sg13g2_a221oi_1 _2548_ (.B2(_1105_),
    .C1(_1152_),
    .B1(_0175_),
    .A1(_1158_),
    .Y(_0176_),
    .A2(_0174_));
 sg13g2_o21ai_1 _2549_ (.B1(_1268_),
    .Y(_0177_),
    .A1(net744),
    .A2(_0176_));
 sg13g2_o21ai_1 _2550_ (.B1(net744),
    .Y(_0178_),
    .A1(net631),
    .A2(_1123_));
 sg13g2_nor2_1 _2551_ (.A(net744),
    .B(_1176_),
    .Y(_0179_));
 sg13g2_o21ai_1 _2552_ (.B1(net717),
    .Y(_0180_),
    .A1(_1025_),
    .A2(_1151_));
 sg13g2_nor2_1 _2553_ (.A(_0179_),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_a21oi_1 _2554_ (.A1(_0178_),
    .A2(_0181_),
    .Y(_0182_),
    .B1(net635));
 sg13g2_a21o_1 _2555_ (.A2(_0182_),
    .A1(_0177_),
    .B1(_0172_),
    .X(_0183_));
 sg13g2_a21oi_2 _2556_ (.B1(_1017_),
    .Y(_0184_),
    .A2(_1110_),
    .A1(net652));
 sg13g2_a221oi_1 _2557_ (.B2(net711),
    .C1(_1139_),
    .B1(_1136_),
    .A1(net651),
    .Y(_0185_),
    .A2(_1109_));
 sg13g2_nand2b_1 _2558_ (.Y(_0186_),
    .B(net674),
    .A_N(_0185_));
 sg13g2_a21oi_1 _2559_ (.A1(_1186_),
    .A2(_1421_),
    .Y(_0187_),
    .B1(_1481_));
 sg13g2_a22oi_1 _2560_ (.Y(_0188_),
    .B1(_1109_),
    .B2(net649),
    .A2(net629),
    .A1(net630));
 sg13g2_or2_1 _2561_ (.X(_0189_),
    .B(_0188_),
    .A(net757));
 sg13g2_a21oi_1 _2562_ (.A1(_1291_),
    .A2(_0189_),
    .Y(_0190_),
    .B1(_1287_));
 sg13g2_mux2_1 _2563_ (.A0(_1143_),
    .A1(_0185_),
    .S(net757),
    .X(_0191_));
 sg13g2_nor2b_1 _2564_ (.A(_0191_),
    .B_N(_1049_),
    .Y(_0192_));
 sg13g2_o21ai_1 _2565_ (.B1(net633),
    .Y(_0193_),
    .A1(_1328_),
    .A2(_0185_));
 sg13g2_nor4_1 _2566_ (.A(_0187_),
    .B(_0190_),
    .C(_0192_),
    .D(_0193_),
    .Y(_0194_));
 sg13g2_o21ai_1 _2567_ (.B1(_1105_),
    .Y(_0195_),
    .A1(net626),
    .A2(_0184_));
 sg13g2_a21oi_1 _2568_ (.A1(net765),
    .A2(_1480_),
    .Y(_0196_),
    .B1(_1278_));
 sg13g2_nand2_1 _2569_ (.Y(_0197_),
    .A(_0195_),
    .B(_0196_));
 sg13g2_o21ai_1 _2570_ (.B1(net752),
    .Y(_0198_),
    .A1(_1137_),
    .A2(net622));
 sg13g2_o21ai_1 _2571_ (.B1(net771),
    .Y(_0199_),
    .A1(net630),
    .A2(net627));
 sg13g2_o21ai_1 _2572_ (.B1(_1143_),
    .Y(_0200_),
    .A1(net763),
    .A2(_1176_));
 sg13g2_nand2b_1 _2573_ (.Y(_0201_),
    .B(_0198_),
    .A_N(_0200_));
 sg13g2_a22oi_1 _2574_ (.Y(_0202_),
    .B1(_0201_),
    .B2(net705),
    .A2(_0197_),
    .A1(net672));
 sg13g2_nand2_1 _2575_ (.Y(_0203_),
    .A(_0194_),
    .B(_0202_));
 sg13g2_nand2_1 _2576_ (.Y(_0204_),
    .A(_1330_),
    .B(_1343_));
 sg13g2_o21ai_1 _2577_ (.B1(net636),
    .Y(_0205_),
    .A1(_1317_),
    .A2(_1356_));
 sg13g2_a221oi_1 _2578_ (.B2(_1295_),
    .C1(_0205_),
    .B1(_1324_),
    .A1(_1049_),
    .Y(_0206_),
    .A2(_1321_));
 sg13g2_a21oi_1 _2579_ (.A1(_0204_),
    .A2(_0206_),
    .Y(_0207_),
    .B1(net668));
 sg13g2_a221oi_1 _2580_ (.B2(_0207_),
    .C1(_1103_),
    .B1(_0203_),
    .A1(net667),
    .Y(_0208_),
    .A2(_0183_));
 sg13g2_or3_1 _2581_ (.A(_1185_),
    .B(_0154_),
    .C(_0208_),
    .X(_0209_));
 sg13g2_or3_1 _2582_ (.A(net732),
    .B(_1136_),
    .C(_1149_),
    .X(_0210_));
 sg13g2_o21ai_1 _2583_ (.B1(_0210_),
    .Y(_0211_),
    .A1(net769),
    .A2(_1163_));
 sg13g2_o21ai_1 _2584_ (.B1(net740),
    .Y(_0212_),
    .A1(_1152_),
    .A2(_0211_));
 sg13g2_a22oi_1 _2585_ (.Y(_0213_),
    .B1(_0212_),
    .B2(_1268_),
    .A2(_0181_),
    .A1(_1273_));
 sg13g2_o21ai_1 _2586_ (.B1(net737),
    .Y(_0214_),
    .A1(_1136_),
    .A2(_0184_));
 sg13g2_nand3_1 _2587_ (.B(_0195_),
    .C(_0214_),
    .A(_1282_),
    .Y(_0215_));
 sg13g2_nor2b_1 _2588_ (.A(_0996_),
    .B_N(_1289_),
    .Y(_0216_));
 sg13g2_o21ai_1 _2589_ (.B1(_1186_),
    .Y(_0217_),
    .A1(net765),
    .A2(_0216_));
 sg13g2_o21ai_1 _2590_ (.B1(_1130_),
    .Y(_0218_),
    .A1(net763),
    .A2(_1176_));
 sg13g2_a22oi_1 _2591_ (.Y(_0219_),
    .B1(net639),
    .B2(net629),
    .A2(net761),
    .A1(net643));
 sg13g2_nor2_1 _2592_ (.A(_1287_),
    .B(_0219_),
    .Y(_0220_));
 sg13g2_a21oi_1 _2593_ (.A1(net705),
    .A2(_0218_),
    .Y(_0221_),
    .B1(_0220_));
 sg13g2_nand2b_1 _2594_ (.Y(_0222_),
    .B(_1327_),
    .A_N(_0191_));
 sg13g2_a21oi_1 _2595_ (.A1(_1049_),
    .A2(_1144_),
    .Y(_0223_),
    .B1(net667));
 sg13g2_nand3_1 _2596_ (.B(_0222_),
    .C(_0223_),
    .A(_0221_),
    .Y(_0224_));
 sg13g2_a221oi_1 _2597_ (.B2(net660),
    .C1(_0224_),
    .B1(_0217_),
    .A1(net672),
    .Y(_0225_),
    .A2(_0215_));
 sg13g2_o21ai_1 _2598_ (.B1(_1063_),
    .Y(_0226_),
    .A1(net663),
    .A2(_0213_));
 sg13g2_nor2_2 _2599_ (.A(net739),
    .B(net733),
    .Y(_0227_));
 sg13g2_o21ai_1 _2600_ (.B1(_0227_),
    .Y(_0228_),
    .A1(net644),
    .A2(_0161_));
 sg13g2_a21o_1 _2601_ (.A2(net639),
    .A1(_1003_),
    .B1(net643),
    .X(_0229_));
 sg13g2_a221oi_1 _2602_ (.B2(net733),
    .C1(net742),
    .B1(_0229_),
    .A1(net773),
    .Y(_0230_),
    .A2(_1290_));
 sg13g2_o21ai_1 _2603_ (.B1(net766),
    .Y(_0231_),
    .A1(_1012_),
    .A2(net624));
 sg13g2_a221oi_1 _2604_ (.B2(net739),
    .C1(net745),
    .B1(_0229_),
    .A1(net729),
    .Y(_0232_),
    .A2(_0155_));
 sg13g2_a221oi_1 _2605_ (.B2(_0232_),
    .C1(net719),
    .B1(_0231_),
    .A1(_0228_),
    .Y(_0233_),
    .A2(_0230_));
 sg13g2_and3_1 _2606_ (.X(_0234_),
    .A(net766),
    .B(_1035_),
    .C(_0165_));
 sg13g2_nor2_1 _2607_ (.A(net760),
    .B(_1158_),
    .Y(_0235_));
 sg13g2_nor3_1 _2608_ (.A(net766),
    .B(_0158_),
    .C(_0235_),
    .Y(_0236_));
 sg13g2_nor3_1 _2609_ (.A(net671),
    .B(_0234_),
    .C(_0236_),
    .Y(_0237_));
 sg13g2_or3_1 _2610_ (.A(_1312_),
    .B(_0233_),
    .C(_0237_),
    .X(_0238_));
 sg13g2_nor3_1 _2611_ (.A(net631),
    .B(_1132_),
    .C(_1315_),
    .Y(_0239_));
 sg13g2_or3_1 _2612_ (.A(_1318_),
    .B(_1319_),
    .C(_0239_),
    .X(_0240_));
 sg13g2_a21o_1 _2613_ (.A2(_1327_),
    .A1(_1321_),
    .B1(net668),
    .X(_0241_));
 sg13g2_a221oi_1 _2614_ (.B2(net721),
    .C1(_0241_),
    .B1(_0240_),
    .A1(_1049_),
    .Y(_0242_),
    .A2(_1330_));
 sg13g2_a21oi_1 _2615_ (.A1(_1326_),
    .A2(_0242_),
    .Y(_0243_),
    .B1(net633));
 sg13g2_a21oi_1 _2616_ (.A1(_0238_),
    .A2(_0243_),
    .Y(_0244_),
    .B1(_1103_));
 sg13g2_o21ai_1 _2617_ (.B1(_0244_),
    .Y(_0245_),
    .A1(_0225_),
    .A2(_0226_));
 sg13g2_nand3_1 _2618_ (.B(_1339_),
    .C(_0148_),
    .A(_1337_),
    .Y(_0246_));
 sg13g2_mux2_1 _2619_ (.A0(_1221_),
    .A1(_1351_),
    .S(net738),
    .X(_0247_));
 sg13g2_nor2_2 _2620_ (.A(net731),
    .B(net659),
    .Y(_0248_));
 sg13g2_a21oi_1 _2621_ (.A1(_1135_),
    .A2(_1172_),
    .Y(_0249_),
    .B1(_1021_));
 sg13g2_nor2_1 _2622_ (.A(net662),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_or2_1 _2623_ (.X(_0251_),
    .B(_0248_),
    .A(_1194_));
 sg13g2_o21ai_1 _2624_ (.B1(_0250_),
    .Y(_0252_),
    .A1(_1356_),
    .A2(_0251_));
 sg13g2_a221oi_1 _2625_ (.B2(net622),
    .C1(_0252_),
    .B1(_0248_),
    .A1(net705),
    .Y(_0253_),
    .A2(_0247_));
 sg13g2_nand3b_1 _2626_ (.B(net634),
    .C(_0246_),
    .Y(_0254_),
    .A_N(_0253_));
 sg13g2_a22oi_1 _2627_ (.Y(_0255_),
    .B1(_0124_),
    .B2(_0125_),
    .A2(net623),
    .A1(net732));
 sg13g2_o21ai_1 _2628_ (.B1(net674),
    .Y(_0256_),
    .A1(net734),
    .A2(_1128_));
 sg13g2_a221oi_1 _2629_ (.B2(net718),
    .C1(net663),
    .B1(net623),
    .A1(net706),
    .Y(_0257_),
    .A2(_1079_));
 sg13g2_o21ai_1 _2630_ (.B1(_0257_),
    .Y(_0258_),
    .A1(_0255_),
    .A2(_0256_));
 sg13g2_nor2_1 _2631_ (.A(net738),
    .B(_1513_),
    .Y(_0259_));
 sg13g2_nand2_1 _2632_ (.Y(_0260_),
    .A(_1479_),
    .B(_1512_));
 sg13g2_o21ai_1 _2633_ (.B1(net674),
    .Y(_0261_),
    .A1(_0259_),
    .A2(_0260_));
 sg13g2_a21oi_1 _2634_ (.A1(_1352_),
    .A2(_0261_),
    .Y(_0262_),
    .B1(net634));
 sg13g2_a21oi_1 _2635_ (.A1(_0258_),
    .A2(_0262_),
    .Y(_0263_),
    .B1(net618));
 sg13g2_a21oi_1 _2636_ (.A1(_0254_),
    .A2(_0263_),
    .Y(_0264_),
    .B1(_1184_));
 sg13g2_a21oi_1 _2637_ (.A1(_0245_),
    .A2(_0264_),
    .Y(_0265_),
    .B1(_1263_));
 sg13g2_a22oi_1 _2638_ (.Y(_0266_),
    .B1(_0184_),
    .B2(net731),
    .A2(_1480_),
    .A1(net765));
 sg13g2_nand2_1 _2639_ (.Y(_0267_),
    .A(net754),
    .B(_1278_));
 sg13g2_a21oi_1 _2640_ (.A1(_0266_),
    .A2(_0267_),
    .Y(_0268_),
    .B1(net670));
 sg13g2_a21oi_1 _2641_ (.A1(_1475_),
    .A2(_0189_),
    .Y(_0269_),
    .B1(_1287_));
 sg13g2_o21ai_1 _2642_ (.B1(net655),
    .Y(_0270_),
    .A1(_1137_),
    .A2(net622));
 sg13g2_nand2b_1 _2643_ (.Y(_0271_),
    .B(_1131_),
    .A_N(_1481_));
 sg13g2_nand4_1 _2644_ (.B(_0186_),
    .C(_0270_),
    .A(net662),
    .Y(_0272_),
    .D(_0271_));
 sg13g2_a21o_1 _2645_ (.A2(_1110_),
    .A1(net651),
    .B1(net637),
    .X(_0273_));
 sg13g2_a21o_1 _2646_ (.A2(_0273_),
    .A1(_1138_),
    .B1(net752),
    .X(_0274_));
 sg13g2_a21oi_1 _2647_ (.A1(_0198_),
    .A2(_0274_),
    .Y(_0275_),
    .B1(_1344_));
 sg13g2_or4_1 _2648_ (.A(_0268_),
    .B(_0269_),
    .C(_0272_),
    .D(_0275_),
    .X(_0276_));
 sg13g2_a221oi_1 _2649_ (.B2(net675),
    .C1(net771),
    .B1(_1149_),
    .A1(net752),
    .Y(_0277_),
    .A2(_1137_));
 sg13g2_o21ai_1 _2650_ (.B1(net705),
    .Y(_0278_),
    .A1(_1264_),
    .A2(_0277_));
 sg13g2_a221oi_1 _2651_ (.B2(net674),
    .C1(net663),
    .B1(_0175_),
    .A1(_1049_),
    .Y(_0279_),
    .A2(_1164_));
 sg13g2_o21ai_1 _2652_ (.B1(_0178_),
    .Y(_0280_),
    .A1(_1030_),
    .A2(_1151_));
 sg13g2_o21ai_1 _2653_ (.B1(net737),
    .Y(_0281_),
    .A1(net630),
    .A2(net627));
 sg13g2_nand2_1 _2654_ (.Y(_0282_),
    .A(_1176_),
    .B(_0281_));
 sg13g2_o21ai_1 _2655_ (.B1(net717),
    .Y(_0283_),
    .A1(_0280_),
    .A2(_0282_));
 sg13g2_nand3_1 _2656_ (.B(_0279_),
    .C(_0283_),
    .A(_0278_),
    .Y(_0284_));
 sg13g2_nand3_1 _2657_ (.B(_0276_),
    .C(_0284_),
    .A(net618),
    .Y(_0285_));
 sg13g2_nand2_1 _2658_ (.Y(_0286_),
    .A(_1209_),
    .B(_1279_));
 sg13g2_a21oi_1 _2659_ (.A1(_1209_),
    .A2(_1279_),
    .Y(_0287_),
    .B1(net772));
 sg13g2_o21ai_1 _2660_ (.B1(net661),
    .Y(_0288_),
    .A1(_1224_),
    .A2(_0287_));
 sg13g2_nand2_1 _2661_ (.Y(_0289_),
    .A(net655),
    .B(_0129_));
 sg13g2_o21ai_1 _2662_ (.B1(_1437_),
    .Y(_0290_),
    .A1(_0959_),
    .A2(_1028_));
 sg13g2_nand2b_1 _2663_ (.Y(_0291_),
    .B(_0290_),
    .A_N(_1031_));
 sg13g2_a21oi_1 _2664_ (.A1(_0124_),
    .A2(_0291_),
    .Y(_0292_),
    .B1(net663));
 sg13g2_nand3_1 _2665_ (.B(net672),
    .C(net623),
    .A(net736),
    .Y(_0293_));
 sg13g2_nand4_1 _2666_ (.B(_0289_),
    .C(_0292_),
    .A(_0288_),
    .Y(_0294_),
    .D(_0293_));
 sg13g2_nor3_1 _2667_ (.A(_1515_),
    .B(_0117_),
    .C(_0259_),
    .Y(_0295_));
 sg13g2_nand2_1 _2668_ (.Y(_0296_),
    .A(net672),
    .B(_1513_));
 sg13g2_o21ai_1 _2669_ (.B1(_0296_),
    .Y(_0297_),
    .A1(net657),
    .A2(_1351_));
 sg13g2_o21ai_1 _2670_ (.B1(net663),
    .Y(_0298_),
    .A1(_0295_),
    .A2(_0297_));
 sg13g2_nand3_1 _2671_ (.B(_0294_),
    .C(_0298_),
    .A(_1103_),
    .Y(_0299_));
 sg13g2_nand3_1 _2672_ (.B(_0285_),
    .C(_0299_),
    .A(net633),
    .Y(_0300_));
 sg13g2_a21o_1 _2673_ (.A2(_1029_),
    .A1(net646),
    .B1(_0134_),
    .X(_0301_));
 sg13g2_nand3_1 _2674_ (.B(_1186_),
    .C(_0301_),
    .A(net723),
    .Y(_0302_));
 sg13g2_o21ai_1 _2675_ (.B1(net718),
    .Y(_0303_),
    .A1(_1028_),
    .A2(_0134_));
 sg13g2_nor3_1 _2676_ (.A(_1029_),
    .B(_1132_),
    .C(_0135_),
    .Y(_0304_));
 sg13g2_o21ai_1 _2677_ (.B1(_0302_),
    .Y(_0305_),
    .A1(_0303_),
    .A2(_0304_));
 sg13g2_nand2_1 _2678_ (.Y(_0306_),
    .A(_0140_),
    .B(_0305_));
 sg13g2_nand3_1 _2679_ (.B(_1232_),
    .C(_1265_),
    .A(net764),
    .Y(_0307_));
 sg13g2_a21o_1 _2680_ (.A2(_0146_),
    .A1(net660),
    .B1(_1286_),
    .X(_0308_));
 sg13g2_a22oi_1 _2681_ (.Y(_0309_),
    .B1(_1162_),
    .B2(net732),
    .A2(_1083_),
    .A1(net645));
 sg13g2_a21oi_1 _2682_ (.A1(_1108_),
    .A2(_0309_),
    .Y(_0310_),
    .B1(net670));
 sg13g2_o21ai_1 _2683_ (.B1(_0149_),
    .Y(_0311_),
    .A1(net731),
    .A2(_1108_));
 sg13g2_a221oi_1 _2684_ (.B2(net740),
    .C1(_0310_),
    .B1(_0311_),
    .A1(_0307_),
    .Y(_0312_),
    .A2(_0308_));
 sg13g2_or4_1 _2685_ (.A(net764),
    .B(net642),
    .C(net637),
    .D(_1149_),
    .X(_0313_));
 sg13g2_a21oi_1 _2686_ (.A1(net734),
    .A2(net622),
    .Y(_0314_),
    .B1(_1369_));
 sg13g2_nand4_1 _2687_ (.B(_0312_),
    .C(_0313_),
    .A(net662),
    .Y(_0315_),
    .D(_0314_));
 sg13g2_a21oi_1 _2688_ (.A1(_0306_),
    .A2(_0315_),
    .Y(_0316_),
    .B1(net619));
 sg13g2_nand2_1 _2689_ (.Y(_0317_),
    .A(net742),
    .B(_0170_));
 sg13g2_a21oi_1 _2690_ (.A1(_1085_),
    .A2(_1161_),
    .Y(_0318_),
    .B1(_1304_));
 sg13g2_nand2_1 _2691_ (.Y(_0319_),
    .A(_1007_),
    .B(_0318_));
 sg13g2_nand3_1 _2692_ (.B(_1166_),
    .C(_1305_),
    .A(_1124_),
    .Y(_0320_));
 sg13g2_a221oi_1 _2693_ (.B2(net707),
    .C1(net719),
    .B1(_0320_),
    .A1(_1064_),
    .Y(_0321_),
    .A2(_0319_));
 sg13g2_o21ai_1 _2694_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_1283_),
    .A2(_0317_));
 sg13g2_a221oi_1 _2695_ (.B2(net679),
    .C1(net712),
    .B1(net681),
    .A1(net703),
    .Y(_0323_),
    .A2(net715));
 sg13g2_nand2_1 _2696_ (.Y(_0324_),
    .A(net640),
    .B(_1004_));
 sg13g2_nor2_1 _2697_ (.A(_1114_),
    .B(_0323_),
    .Y(_0325_));
 sg13g2_o21ai_1 _2698_ (.B1(_0164_),
    .Y(_0326_),
    .A1(net760),
    .A2(_0325_));
 sg13g2_nand2_1 _2699_ (.Y(_0327_),
    .A(net767),
    .B(_0326_));
 sg13g2_o21ai_1 _2700_ (.B1(net739),
    .Y(_0328_),
    .A1(net624),
    .A2(_0323_));
 sg13g2_o21ai_1 _2701_ (.B1(_0328_),
    .Y(_0329_),
    .A1(_1044_),
    .A2(_0325_));
 sg13g2_nor2_1 _2702_ (.A(net658),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_a221oi_1 _2703_ (.B2(_0157_),
    .C1(_1304_),
    .B1(net639),
    .A1(net640),
    .Y(_0331_),
    .A2(_1004_));
 sg13g2_nand2b_1 _2704_ (.Y(_0332_),
    .B(net746),
    .A_N(_0331_));
 sg13g2_a221oi_1 _2705_ (.B2(net673),
    .C1(net664),
    .B1(_0331_),
    .A1(_0327_),
    .Y(_0333_),
    .A2(_0330_));
 sg13g2_nand2b_1 _2706_ (.Y(_0334_),
    .B(_1343_),
    .A_N(_1321_));
 sg13g2_a21oi_1 _2707_ (.A1(net760),
    .A2(_1416_),
    .Y(_0335_),
    .B1(_1219_));
 sg13g2_and2_1 _2708_ (.A(net655),
    .B(_1329_),
    .X(_0336_));
 sg13g2_a221oi_1 _2709_ (.B2(_0336_),
    .C1(net669),
    .B1(_0335_),
    .A1(_0934_),
    .Y(_0337_),
    .A2(_1317_));
 sg13g2_a221oi_1 _2710_ (.B2(_0337_),
    .C1(_1103_),
    .B1(_0334_),
    .A1(_0322_),
    .Y(_0338_),
    .A2(_0333_));
 sg13g2_o21ai_1 _2711_ (.B1(net634),
    .Y(_0339_),
    .A1(_0316_),
    .A2(_0338_));
 sg13g2_nand3_1 _2712_ (.B(_0300_),
    .C(_0339_),
    .A(_1185_),
    .Y(_0340_));
 sg13g2_a21oi_1 _2713_ (.A1(_0324_),
    .A2(_0335_),
    .Y(_0341_),
    .B1(net773));
 sg13g2_nor3_1 _2714_ (.A(net725),
    .B(_0329_),
    .C(_0341_),
    .Y(_0342_));
 sg13g2_nand3_1 _2715_ (.B(_1124_),
    .C(_1166_),
    .A(net707),
    .Y(_0343_));
 sg13g2_nand2_1 _2716_ (.Y(_0344_),
    .A(net730),
    .B(_1065_));
 sg13g2_a21oi_1 _2717_ (.A1(net652),
    .A2(_1119_),
    .Y(_0345_),
    .B1(net745));
 sg13g2_a22oi_1 _2718_ (.Y(_0346_),
    .B1(_0345_),
    .B2(net730),
    .A2(_0344_),
    .A1(_1221_));
 sg13g2_nand2_1 _2719_ (.Y(_0347_),
    .A(_0343_),
    .B(_0346_));
 sg13g2_nor2_1 _2720_ (.A(net720),
    .B(net624),
    .Y(_0348_));
 sg13g2_a221oi_1 _2721_ (.B2(_0348_),
    .C1(net664),
    .B1(_0347_),
    .A1(_0332_),
    .Y(_0349_),
    .A2(_0342_));
 sg13g2_nand2_1 _2722_ (.Y(_0350_),
    .A(_1286_),
    .B(_0129_));
 sg13g2_a22oi_1 _2723_ (.Y(_0351_),
    .B1(_1316_),
    .B2(net653),
    .A2(_1218_),
    .A1(_1074_));
 sg13g2_nor3_1 _2724_ (.A(net648),
    .B(_1028_),
    .C(_1085_),
    .Y(_0352_));
 sg13g2_nor4_1 _2725_ (.A(net720),
    .B(_1024_),
    .C(_0351_),
    .D(_0352_),
    .Y(_0353_));
 sg13g2_a21oi_1 _2726_ (.A1(net639),
    .A2(net656),
    .Y(_0354_),
    .B1(_1416_));
 sg13g2_inv_1 _2727_ (.Y(_0355_),
    .A(_0354_));
 sg13g2_a21oi_1 _2728_ (.A1(_0962_),
    .A2(net755),
    .Y(_0356_),
    .B1(_1296_));
 sg13g2_a221oi_1 _2729_ (.B2(_0356_),
    .C1(_0353_),
    .B1(_0355_),
    .A1(net721),
    .Y(_0357_),
    .A2(_0239_));
 sg13g2_a21oi_1 _2730_ (.A1(_0350_),
    .A2(_0357_),
    .Y(_0358_),
    .B1(net669));
 sg13g2_o21ai_1 _2731_ (.B1(_1062_),
    .Y(_0359_),
    .A1(_0349_),
    .A2(_0358_));
 sg13g2_a21o_1 _2732_ (.A2(_0274_),
    .A1(_0198_),
    .B1(_1296_),
    .X(_0360_));
 sg13g2_nor2b_1 _2733_ (.A(_0186_),
    .B_N(_0227_),
    .Y(_0361_));
 sg13g2_nand2_1 _2734_ (.Y(_0362_),
    .A(_1336_),
    .B(_1437_));
 sg13g2_a21oi_1 _2735_ (.A1(_1138_),
    .A2(_0273_),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_nor3_1 _2736_ (.A(net698),
    .B(_0965_),
    .C(_1287_),
    .Y(_0364_));
 sg13g2_a22oi_1 _2737_ (.Y(_0365_),
    .B1(_0248_),
    .B2(net637),
    .A2(_1131_),
    .A1(net660));
 sg13g2_a22oi_1 _2738_ (.Y(_0366_),
    .B1(_0364_),
    .B2(net649),
    .A2(_0184_),
    .A1(_1327_));
 sg13g2_nand3_1 _2739_ (.B(_0365_),
    .C(_0366_),
    .A(net662),
    .Y(_0367_));
 sg13g2_or2_1 _2740_ (.X(_0368_),
    .B(_1479_),
    .A(_1044_));
 sg13g2_a21oi_1 _2741_ (.A1(_0266_),
    .A2(_0368_),
    .Y(_0369_),
    .B1(net670));
 sg13g2_nor4_1 _2742_ (.A(_0361_),
    .B(_0363_),
    .C(_0367_),
    .D(_0369_),
    .Y(_0370_));
 sg13g2_o21ai_1 _2743_ (.B1(net763),
    .Y(_0371_),
    .A1(_1137_),
    .A2(net622));
 sg13g2_nand3b_1 _2744_ (.B(_0371_),
    .C(_0199_),
    .Y(_0372_),
    .A_N(_0280_));
 sg13g2_a22oi_1 _2745_ (.Y(_0373_),
    .B1(_1158_),
    .B2(net763),
    .A2(net737),
    .A1(net713));
 sg13g2_nor2_1 _2746_ (.A(_0934_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_a221oi_1 _2747_ (.B2(net717),
    .C1(_0374_),
    .B1(_0372_),
    .A1(_1166_),
    .Y(_0375_),
    .A2(net655));
 sg13g2_a221oi_1 _2748_ (.B2(_0279_),
    .C1(net635),
    .B1(_0375_),
    .A1(_0360_),
    .Y(_0376_),
    .A2(_0370_));
 sg13g2_nand3b_1 _2749_ (.B(net619),
    .C(_0359_),
    .Y(_0377_),
    .A_N(_0376_));
 sg13g2_nor2_1 _2750_ (.A(net764),
    .B(_0135_),
    .Y(_0378_));
 sg13g2_a21oi_1 _2751_ (.A1(net638),
    .A2(net625),
    .Y(_0379_),
    .B1(_1106_));
 sg13g2_nor3_1 _2752_ (.A(net771),
    .B(net642),
    .C(_1241_),
    .Y(_0380_));
 sg13g2_nor4_1 _2753_ (.A(net657),
    .B(_0378_),
    .C(_0379_),
    .D(_0380_),
    .Y(_0381_));
 sg13g2_nand4_1 _2754_ (.B(_1138_),
    .C(_1140_),
    .A(net723),
    .Y(_0382_),
    .D(_0301_));
 sg13g2_o21ai_1 _2755_ (.B1(_0382_),
    .Y(_0383_),
    .A1(net670),
    .A2(_0136_));
 sg13g2_o21ai_1 _2756_ (.B1(net666),
    .Y(_0384_),
    .A1(_0381_),
    .A2(_0383_));
 sg13g2_o21ai_1 _2757_ (.B1(_0313_),
    .Y(_0385_),
    .A1(net770),
    .A2(_0149_));
 sg13g2_nor2_1 _2758_ (.A(net666),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_a21oi_1 _2759_ (.A1(_0312_),
    .A2(_0386_),
    .Y(_0387_),
    .B1(net633));
 sg13g2_a22oi_1 _2760_ (.Y(_0388_),
    .B1(_0286_),
    .B2(net728),
    .A2(_0118_),
    .A1(net765));
 sg13g2_a22oi_1 _2761_ (.Y(_0389_),
    .B1(_1279_),
    .B2(_0123_),
    .A2(net736),
    .A1(net740));
 sg13g2_nor2_1 _2762_ (.A(_0959_),
    .B(_1030_),
    .Y(_0390_));
 sg13g2_nor2_1 _2763_ (.A(net718),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_a221oi_1 _2764_ (.B2(_0124_),
    .C1(net663),
    .B1(_0391_),
    .A1(net718),
    .Y(_0392_),
    .A2(_0389_));
 sg13g2_o21ai_1 _2765_ (.B1(_0392_),
    .Y(_0393_),
    .A1(net657),
    .A2(_0388_));
 sg13g2_nand2_1 _2766_ (.Y(_0394_),
    .A(_1287_),
    .B(_1514_));
 sg13g2_a21o_1 _2767_ (.A2(_1453_),
    .A1(_1417_),
    .B1(_1287_),
    .X(_0395_));
 sg13g2_nand3_1 _2768_ (.B(_0394_),
    .C(_0395_),
    .A(net663),
    .Y(_0396_));
 sg13g2_nand3_1 _2769_ (.B(_0393_),
    .C(_0396_),
    .A(net633),
    .Y(_0397_));
 sg13g2_a21oi_1 _2770_ (.A1(_0384_),
    .A2(_0387_),
    .Y(_0398_),
    .B1(net619));
 sg13g2_a21oi_1 _2771_ (.A1(_0397_),
    .A2(_0398_),
    .Y(_0399_),
    .B1(_1185_));
 sg13g2_a21oi_1 _2772_ (.A1(_0377_),
    .A2(_0399_),
    .Y(_0400_),
    .B1(_1262_));
 sg13g2_a221oi_1 _2773_ (.B2(_0400_),
    .C1(_1509_),
    .B1(_0340_),
    .A1(_0209_),
    .Y(_0401_),
    .A2(_0265_));
 sg13g2_xor2_1 _2774_ (.B(\pix_y[9] ),
    .A(net793),
    .X(_0402_));
 sg13g2_a21oi_1 _2775_ (.A1(_0759_),
    .A2(\pix_y[8] ),
    .Y(_0403_),
    .B1(_0402_));
 sg13g2_nand2_1 _2776_ (.Y(_0404_),
    .A(net794),
    .B(_0775_));
 sg13g2_o21ai_1 _2777_ (.B1(_1101_),
    .Y(_0405_),
    .A1(\logo_top[6] ),
    .A2(_0772_));
 sg13g2_nor2_1 _2778_ (.A(net794),
    .B(_0775_),
    .Y(_0406_));
 sg13g2_a21oi_1 _2779_ (.A1(_0404_),
    .A2(_0405_),
    .Y(_0407_),
    .B1(_0406_));
 sg13g2_nor2b_1 _2780_ (.A(\pix_x[8] ),
    .B_N(\logo_left[8] ),
    .Y(_0408_));
 sg13g2_xor2_1 _2781_ (.B(\pix_x[8] ),
    .A(\logo_left[8] ),
    .X(_0409_));
 sg13g2_nor2b_1 _2782_ (.A(net796),
    .B_N(\pix_x[7] ),
    .Y(_0410_));
 sg13g2_and2_1 _2783_ (.A(_0970_),
    .B(net686),
    .X(_0411_));
 sg13g2_nor2b_1 _2784_ (.A(\pix_x[7] ),
    .B_N(net796),
    .Y(_0412_));
 sg13g2_nor3_1 _2785_ (.A(_0410_),
    .B(_0411_),
    .C(_0412_),
    .Y(_0413_));
 sg13g2_o21ai_1 _2786_ (.B1(_0409_),
    .Y(_0414_),
    .A1(_0410_),
    .A2(_0413_));
 sg13g2_a21o_1 _2787_ (.A2(_0412_),
    .A1(_0409_),
    .B1(_0410_),
    .X(_0415_));
 sg13g2_a21o_1 _2788_ (.A2(_0415_),
    .A1(_0411_),
    .B1(_0413_),
    .X(_0416_));
 sg13g2_nor2_1 _2789_ (.A(_0759_),
    .B(\pix_y[8] ),
    .Y(_0417_));
 sg13g2_xnor2_1 _2790_ (.Y(_0418_),
    .A(_0402_),
    .B(_0417_));
 sg13g2_xor2_1 _2791_ (.B(\pix_x[9] ),
    .A(\logo_left[9] ),
    .X(_0419_));
 sg13g2_xnor2_1 _2792_ (.Y(_0420_),
    .A(_0408_),
    .B(_0419_));
 sg13g2_nand4_1 _2793_ (.B(_0416_),
    .C(_0418_),
    .A(_0414_),
    .Y(_0421_),
    .D(_0420_));
 sg13g2_a21oi_1 _2794_ (.A1(_0405_),
    .A2(_0406_),
    .Y(_0422_),
    .B1(_0421_));
 sg13g2_nor2_1 _2795_ (.A(_0404_),
    .B(_0405_),
    .Y(_0423_));
 sg13g2_o21ai_1 _2796_ (.B1(_0422_),
    .Y(_0424_),
    .A1(_0403_),
    .A2(_0423_));
 sg13g2_a21oi_1 _2797_ (.A1(_0403_),
    .A2(_0407_),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_or2_1 _2798_ (.X(_0426_),
    .B(_0425_),
    .A(net2));
 sg13g2_nor2_1 _2799_ (.A(net805),
    .B(\pix_y[9] ),
    .Y(_0427_));
 sg13g2_o21ai_1 _2800_ (.B1(\pix_x[9] ),
    .Y(_0428_),
    .A1(\pix_x[7] ),
    .A2(\pix_x[8] ));
 sg13g2_nand4_1 _2801_ (.B(_0426_),
    .C(_0427_),
    .A(_0797_),
    .Y(_0429_),
    .D(_0428_));
 sg13g2_xnor2_1 _2802_ (.Y(_0430_),
    .A(net799),
    .B(net666));
 sg13g2_nand2b_1 _2803_ (.Y(_0431_),
    .B(net669),
    .A_N(_0008_));
 sg13g2_o21ai_1 _2804_ (.B1(_0431_),
    .Y(_0432_),
    .A1(net711),
    .A2(_0430_));
 sg13g2_nor2_1 _2805_ (.A(_0764_),
    .B(net634),
    .Y(_0433_));
 sg13g2_xnor2_1 _2806_ (.Y(_0434_),
    .A(net798),
    .B(net634));
 sg13g2_xnor2_1 _2807_ (.Y(_0435_),
    .A(net701),
    .B(_0434_));
 sg13g2_xnor2_1 _2808_ (.Y(_0436_),
    .A(net710),
    .B(_0430_));
 sg13g2_nand2_1 _2809_ (.Y(_0437_),
    .A(net800),
    .B(net724));
 sg13g2_xnor2_1 _2810_ (.Y(_0438_),
    .A(net800),
    .B(net724));
 sg13g2_o21ai_1 _2811_ (.B1(_0437_),
    .Y(_0439_),
    .A1(net713),
    .A2(_0438_));
 sg13g2_nand2_1 _2812_ (.Y(_0440_),
    .A(_0436_),
    .B(_0439_));
 sg13g2_nand2_1 _2813_ (.Y(_0441_),
    .A(_0007_),
    .B(_1509_));
 sg13g2_xnor2_1 _2814_ (.Y(_0442_),
    .A(net715),
    .B(_0438_));
 sg13g2_and2_1 _2815_ (.A(_0441_),
    .B(_0442_),
    .X(_0443_));
 sg13g2_xnor2_1 _2816_ (.Y(_0444_),
    .A(\pix_x[2] ),
    .B(_0939_));
 sg13g2_nor2_1 _2817_ (.A(net741),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_xnor2_1 _2818_ (.Y(_0446_),
    .A(_0441_),
    .B(_0442_));
 sg13g2_nor3_1 _2819_ (.A(net741),
    .B(_0444_),
    .C(_0446_),
    .Y(_0447_));
 sg13g2_xor2_1 _2820_ (.B(_0439_),
    .A(_0436_),
    .X(_0448_));
 sg13g2_o21ai_1 _2821_ (.B1(_0448_),
    .Y(_0449_),
    .A1(_0443_),
    .A2(_0447_));
 sg13g2_xnor2_1 _2822_ (.Y(_0450_),
    .A(_0432_),
    .B(_0435_));
 sg13g2_a21oi_1 _2823_ (.A1(_0440_),
    .A2(_0449_),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_a21oi_1 _2824_ (.A1(_0432_),
    .A2(_0435_),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_a21oi_1 _2825_ (.A1(net694),
    .A2(_0434_),
    .Y(_0453_),
    .B1(_0433_));
 sg13g2_xnor2_1 _2826_ (.Y(_0454_),
    .A(net797),
    .B(net651));
 sg13g2_xnor2_1 _2827_ (.Y(_0455_),
    .A(_1103_),
    .B(_0454_));
 sg13g2_xnor2_1 _2828_ (.Y(_0456_),
    .A(_0453_),
    .B(_0455_));
 sg13g2_xor2_1 _2829_ (.B(_0456_),
    .A(_0452_),
    .X(_0457_));
 sg13g2_nor2_1 _2830_ (.A(net806),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_a21oi_1 _2831_ (.A1(net806),
    .A2(net171),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_nor4_1 _2832_ (.A(_1511_),
    .B(_0401_),
    .C(_0429_),
    .D(_0459_),
    .Y(_0022_));
 sg13g2_nor2b_1 _2833_ (.A(net168),
    .B_N(net807),
    .Y(_0460_));
 sg13g2_nor4_1 _2834_ (.A(_1511_),
    .B(_0401_),
    .C(_0429_),
    .D(_0460_),
    .Y(_0023_));
 sg13g2_nor2b_1 _2835_ (.A(\gamepad.driver.pmod_latch_prev ),
    .B_N(\gamepad.driver.pmod_latch_sync[1] ),
    .Y(_0461_));
 sg13g2_nor2_1 _2836_ (.A(_0773_),
    .B(net779),
    .Y(_0462_));
 sg13g2_a22oi_1 _2837_ (.Y(_0024_),
    .B1(net750),
    .B2(_0781_),
    .A2(net778),
    .A1(_0754_));
 sg13g2_a22oi_1 _2838_ (.Y(_0025_),
    .B1(net750),
    .B2(_0780_),
    .A2(net778),
    .A1(_0753_));
 sg13g2_a22oi_1 _2839_ (.Y(_0026_),
    .B1(net750),
    .B2(_0783_),
    .A2(net778),
    .A1(_0752_));
 sg13g2_a22oi_1 _2840_ (.Y(_0027_),
    .B1(net750),
    .B2(_0782_),
    .A2(net778),
    .A1(_0751_));
 sg13g2_a22oi_1 _2841_ (.Y(_0028_),
    .B1(net751),
    .B2(_0785_),
    .A2(net779),
    .A1(_0750_));
 sg13g2_a22oi_1 _2842_ (.Y(_0029_),
    .B1(net751),
    .B2(_0784_),
    .A2(net779),
    .A1(_0749_));
 sg13g2_a22oi_1 _2843_ (.Y(_0030_),
    .B1(net751),
    .B2(_0787_),
    .A2(net779),
    .A1(_0748_));
 sg13g2_a22oi_1 _2844_ (.Y(_0031_),
    .B1(net751),
    .B2(_0786_),
    .A2(net779),
    .A1(_0747_));
 sg13g2_a22oi_1 _2845_ (.Y(_0032_),
    .B1(net750),
    .B2(_0789_),
    .A2(net778),
    .A1(_0746_));
 sg13g2_a22oi_1 _2846_ (.Y(_0033_),
    .B1(net750),
    .B2(_0788_),
    .A2(net778),
    .A1(_0745_));
 sg13g2_a22oi_1 _2847_ (.Y(_0034_),
    .B1(net750),
    .B2(_0791_),
    .A2(net778),
    .A1(_0744_));
 sg13g2_a22oi_1 _2848_ (.Y(_0035_),
    .B1(net750),
    .B2(_0790_),
    .A2(net778),
    .A1(_0767_));
 sg13g2_nand2_1 _2849_ (.Y(_0463_),
    .A(net152),
    .B(_0824_));
 sg13g2_nand4_1 _2850_ (.B(\gamepad.decoder.data_reg[8] ),
    .C(\gamepad.decoder.data_reg[11] ),
    .A(\gamepad.decoder.data_reg[9] ),
    .Y(_0464_),
    .D(\gamepad.decoder.data_reg[10] ));
 sg13g2_nand4_1 _2851_ (.B(\gamepad.decoder.data_reg[4] ),
    .C(\gamepad.decoder.data_reg[7] ),
    .A(\gamepad.decoder.data_reg[5] ),
    .Y(_0465_),
    .D(\gamepad.decoder.data_reg[6] ));
 sg13g2_nand4_1 _2852_ (.B(\gamepad.decoder.data_reg[0] ),
    .C(\gamepad.decoder.data_reg[3] ),
    .A(\gamepad.decoder.data_reg[1] ),
    .Y(_0466_),
    .D(\gamepad.decoder.data_reg[2] ));
 sg13g2_or3_2 _2853_ (.A(_0464_),
    .B(_0465_),
    .C(_0466_),
    .X(_0467_));
 sg13g2_nand3_1 _2854_ (.B(_0823_),
    .C(_0467_),
    .A(\gamepad.decoder.data_reg[8] ),
    .Y(_0468_));
 sg13g2_a21oi_1 _2855_ (.A1(_0463_),
    .A2(_0468_),
    .Y(_0036_),
    .B1(_0773_));
 sg13g2_and3_1 _2856_ (.X(_0469_),
    .A(\pix_x[0] ),
    .B(net211),
    .C(\pix_x[1] ));
 sg13g2_and2_1 _2857_ (.A(net227),
    .B(_0469_),
    .X(_0470_));
 sg13g2_nand2_1 _2858_ (.Y(_0471_),
    .A(net235),
    .B(_0470_));
 sg13g2_nand3b_1 _2859_ (.B(\pix_x[8] ),
    .C(\pix_x[9] ),
    .Y(_0472_),
    .A_N(\pix_x[7] ));
 sg13g2_nor4_2 _2860_ (.A(\pix_x[5] ),
    .B(net217),
    .C(_0471_),
    .Y(_0473_),
    .D(_0472_));
 sg13g2_nand2b_1 _2861_ (.Y(_0474_),
    .B(net810),
    .A_N(_0473_));
 sg13g2_nor2_1 _2862_ (.A(_0794_),
    .B(net654),
    .Y(_0037_));
 sg13g2_xnor2_1 _2863_ (.Y(_0475_),
    .A(\pix_x[0] ),
    .B(net222));
 sg13g2_nor2_1 _2864_ (.A(_0474_),
    .B(net223),
    .Y(_0038_));
 sg13g2_a21oi_1 _2865_ (.A1(\pix_x[0] ),
    .A2(\pix_x[1] ),
    .Y(_0476_),
    .B1(net211));
 sg13g2_nor3_1 _2866_ (.A(net805),
    .B(_0469_),
    .C(net212),
    .Y(_0039_));
 sg13g2_o21ai_1 _2867_ (.B1(net810),
    .Y(_0477_),
    .A1(net227),
    .A2(_0469_));
 sg13g2_nor2_1 _2868_ (.A(_0470_),
    .B(net228),
    .Y(_0040_));
 sg13g2_o21ai_1 _2869_ (.B1(net810),
    .Y(_0478_),
    .A1(net235),
    .A2(_0470_));
 sg13g2_nor2b_1 _2870_ (.A(_0478_),
    .B_N(_0471_),
    .Y(_0041_));
 sg13g2_xor2_1 _2871_ (.B(_0471_),
    .A(net249),
    .X(_0479_));
 sg13g2_nor2_1 _2872_ (.A(net654),
    .B(_0479_),
    .Y(_0042_));
 sg13g2_a21oi_1 _2873_ (.A1(_0801_),
    .A2(_0470_),
    .Y(_0480_),
    .B1(net217));
 sg13g2_and2_1 _2874_ (.A(_0802_),
    .B(_0470_),
    .X(_0481_));
 sg13g2_nor3_1 _2875_ (.A(net654),
    .B(net218),
    .C(_0481_),
    .Y(_0043_));
 sg13g2_xnor2_1 _2876_ (.Y(_0482_),
    .A(net243),
    .B(_0481_));
 sg13g2_nor2_1 _2877_ (.A(net654),
    .B(_0482_),
    .Y(_0044_));
 sg13g2_a21oi_1 _2878_ (.A1(\pix_x[7] ),
    .A2(_0481_),
    .Y(_0483_),
    .B1(net233));
 sg13g2_and3_1 _2879_ (.X(_0484_),
    .A(net246),
    .B(\pix_x[8] ),
    .C(_0481_));
 sg13g2_nor3_1 _2880_ (.A(net654),
    .B(net234),
    .C(_0484_),
    .Y(_0045_));
 sg13g2_a21oi_1 _2881_ (.A1(net224),
    .A2(_0484_),
    .Y(_0485_),
    .B1(net654));
 sg13g2_o21ai_1 _2882_ (.B1(_0485_),
    .Y(_0486_),
    .A1(net224),
    .A2(_0484_));
 sg13g2_inv_1 _2883_ (.Y(_0046_),
    .A(_0486_));
 sg13g2_and2_1 _2884_ (.A(\gamepad.decoder.data_reg[5] ),
    .B(_0467_),
    .X(_0487_));
 sg13g2_or2_1 _2885_ (.X(_0488_),
    .B(\logo_left[8] ),
    .A(\logo_left[9] ));
 sg13g2_o21ai_1 _2886_ (.B1(_0487_),
    .Y(_0489_),
    .A1(_0884_),
    .A2(_0488_));
 sg13g2_and4_1 _2887_ (.A(\gamepad.decoder.data_reg[4] ),
    .B(_0866_),
    .C(_0897_),
    .D(_0467_),
    .X(_0490_));
 sg13g2_nor2_1 _2888_ (.A(net780),
    .B(net620),
    .Y(_0491_));
 sg13g2_a21oi_1 _2889_ (.A1(_0489_),
    .A2(_0491_),
    .Y(_0492_),
    .B1(_0824_));
 sg13g2_o21ai_1 _2890_ (.B1(net811),
    .Y(_0493_),
    .A1(net804),
    .A2(net616));
 sg13g2_a21oi_1 _2891_ (.A1(_0766_),
    .A2(net616),
    .Y(_0047_),
    .B1(_0493_));
 sg13g2_xor2_1 _2892_ (.B(net804),
    .A(net802),
    .X(_0494_));
 sg13g2_xnor2_1 _2893_ (.Y(_0495_),
    .A(net620),
    .B(_0494_));
 sg13g2_xor2_1 _2894_ (.B(net802),
    .A(net792),
    .X(_0496_));
 sg13g2_xnor2_1 _2895_ (.Y(_0497_),
    .A(net133),
    .B(_0496_));
 sg13g2_o21ai_1 _2896_ (.B1(net616),
    .Y(_0498_),
    .A1(net784),
    .A2(_0497_));
 sg13g2_a21oi_1 _2897_ (.A1(net784),
    .A2(_0495_),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_o21ai_1 _2898_ (.B1(net811),
    .Y(_0500_),
    .A1(net802),
    .A2(net616));
 sg13g2_nor2_1 _2899_ (.A(_0499_),
    .B(_0500_),
    .Y(_0048_));
 sg13g2_xnor2_1 _2900_ (.Y(_0501_),
    .A(_0007_),
    .B(_0879_));
 sg13g2_nor2_1 _2901_ (.A(net620),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_xor2_1 _2902_ (.B(_0860_),
    .A(net801),
    .X(_0503_));
 sg13g2_a21oi_1 _2903_ (.A1(net620),
    .A2(_0503_),
    .Y(_0504_),
    .B1(_0502_));
 sg13g2_xnor2_1 _2904_ (.Y(_0505_),
    .A(net792),
    .B(net801));
 sg13g2_a21oi_1 _2905_ (.A1(net792),
    .A2(_0860_),
    .Y(_0506_),
    .B1(_0879_));
 sg13g2_and2_1 _2906_ (.A(_0505_),
    .B(_0506_),
    .X(_0507_));
 sg13g2_o21ai_1 _2907_ (.B1(net780),
    .Y(_0508_),
    .A1(_0505_),
    .A2(_0506_));
 sg13g2_o21ai_1 _2908_ (.B1(net616),
    .Y(_0509_),
    .A1(_0507_),
    .A2(_0508_));
 sg13g2_a21oi_1 _2909_ (.A1(net784),
    .A2(_0504_),
    .Y(_0510_),
    .B1(_0509_));
 sg13g2_o21ai_1 _2910_ (.B1(net811),
    .Y(_0511_),
    .A1(net801),
    .A2(net616));
 sg13g2_nor2_1 _2911_ (.A(_0510_),
    .B(_0511_),
    .Y(_0049_));
 sg13g2_mux2_1 _2912_ (.A0(_0891_),
    .A1(_0876_),
    .S(net620),
    .X(_0512_));
 sg13g2_nand2b_1 _2913_ (.Y(_0513_),
    .B(net792),
    .A_N(net800));
 sg13g2_xnor2_1 _2914_ (.Y(_0514_),
    .A(net792),
    .B(net800));
 sg13g2_a21oi_1 _2915_ (.A1(_0758_),
    .A2(net801),
    .Y(_0515_),
    .B1(_0507_));
 sg13g2_xnor2_1 _2916_ (.Y(_0516_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_o21ai_1 _2917_ (.B1(net616),
    .Y(_0517_),
    .A1(net784),
    .A2(_0516_));
 sg13g2_a21o_1 _2918_ (.A2(_0512_),
    .A1(net784),
    .B1(_0517_),
    .X(_0518_));
 sg13g2_nand2b_1 _2919_ (.Y(_0519_),
    .B(net800),
    .A_N(net616));
 sg13g2_nand3_1 _2920_ (.B(_0518_),
    .C(_0519_),
    .A(net815),
    .Y(_0050_));
 sg13g2_nand2_1 _2921_ (.Y(_0520_),
    .A(_0008_),
    .B(_0881_));
 sg13g2_xnor2_1 _2922_ (.Y(_0521_),
    .A(net258),
    .B(_0881_));
 sg13g2_a21oi_1 _2923_ (.A1(_0872_),
    .A2(net621),
    .Y(_0522_),
    .B1(net780));
 sg13g2_o21ai_1 _2924_ (.B1(_0522_),
    .Y(_0523_),
    .A1(net620),
    .A2(_0521_));
 sg13g2_xnor2_1 _2925_ (.Y(_0524_),
    .A(net791),
    .B(net799));
 sg13g2_a22oi_1 _2926_ (.Y(_0525_),
    .B1(_0507_),
    .B2(_0513_),
    .A2(_0880_),
    .A1(_0758_));
 sg13g2_nand2b_1 _2927_ (.Y(_0526_),
    .B(_0524_),
    .A_N(_0525_));
 sg13g2_xnor2_1 _2928_ (.Y(_0527_),
    .A(_0524_),
    .B(_0525_));
 sg13g2_a221oi_1 _2929_ (.B2(net780),
    .C1(_0824_),
    .B1(_0527_),
    .A1(_0489_),
    .Y(_0528_),
    .A2(_0491_));
 sg13g2_o21ai_1 _2930_ (.B1(net815),
    .Y(_0529_),
    .A1(net799),
    .A2(net615));
 sg13g2_a21oi_1 _2931_ (.A1(_0523_),
    .A2(_0528_),
    .Y(_0051_),
    .B1(_0529_));
 sg13g2_xnor2_1 _2932_ (.Y(_0530_),
    .A(net798),
    .B(_0520_));
 sg13g2_xor2_1 _2933_ (.B(net798),
    .A(net791),
    .X(_0531_));
 sg13g2_o21ai_1 _2934_ (.B1(_0526_),
    .Y(_0532_),
    .A1(net791),
    .A2(_0765_));
 sg13g2_nor2_1 _2935_ (.A(net621),
    .B(_0530_),
    .Y(_0533_));
 sg13g2_a21oi_1 _2936_ (.A1(_0871_),
    .A2(net621),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_xor2_1 _2937_ (.B(_0532_),
    .A(_0531_),
    .X(_0535_));
 sg13g2_o21ai_1 _2938_ (.B1(net615),
    .Y(_0536_),
    .A1(net784),
    .A2(_0535_));
 sg13g2_a21oi_1 _2939_ (.A1(net784),
    .A2(_0534_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_o21ai_1 _2940_ (.B1(net815),
    .Y(_0538_),
    .A1(net798),
    .A2(net615));
 sg13g2_nor2_1 _2941_ (.A(_0537_),
    .B(_0538_),
    .Y(_0052_));
 sg13g2_mux2_1 _2942_ (.A0(_0888_),
    .A1(_0874_),
    .S(net621),
    .X(_0539_));
 sg13g2_nor2_1 _2943_ (.A(net780),
    .B(_0539_),
    .Y(_0540_));
 sg13g2_nand2_1 _2944_ (.Y(_0541_),
    .A(_0758_),
    .B(net797));
 sg13g2_xor2_1 _2945_ (.B(net797),
    .A(net791),
    .X(_0542_));
 sg13g2_nor2_1 _2946_ (.A(_0526_),
    .B(_0531_),
    .Y(_0543_));
 sg13g2_nor2_1 _2947_ (.A(dir_x),
    .B(_0882_),
    .Y(_0544_));
 sg13g2_nor2_1 _2948_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_or2_1 _2949_ (.X(_0546_),
    .B(_0545_),
    .A(_0542_));
 sg13g2_a21oi_1 _2950_ (.A1(_0542_),
    .A2(_0545_),
    .Y(_0547_),
    .B1(net786));
 sg13g2_and2_1 _2951_ (.A(_0546_),
    .B(_0547_),
    .X(_0548_));
 sg13g2_nand2b_1 _2952_ (.Y(_0549_),
    .B(net797),
    .A_N(net615));
 sg13g2_o21ai_1 _2953_ (.B1(net617),
    .Y(_0550_),
    .A1(_0540_),
    .A2(_0548_));
 sg13g2_nand3_1 _2954_ (.B(_0549_),
    .C(_0550_),
    .A(net814),
    .Y(_0053_));
 sg13g2_xnor2_1 _2955_ (.Y(_0551_),
    .A(net796),
    .B(_0887_));
 sg13g2_o21ai_1 _2956_ (.B1(net786),
    .Y(_0552_),
    .A1(net621),
    .A2(_0551_));
 sg13g2_a21oi_1 _2957_ (.A1(_0869_),
    .A2(net620),
    .Y(_0553_),
    .B1(_0552_));
 sg13g2_xor2_1 _2958_ (.B(net796),
    .A(net791),
    .X(_0554_));
 sg13g2_a21oi_1 _2959_ (.A1(_0541_),
    .A2(_0546_),
    .Y(_0555_),
    .B1(_0554_));
 sg13g2_and3_1 _2960_ (.X(_0556_),
    .A(_0541_),
    .B(_0546_),
    .C(_0554_));
 sg13g2_nor3_1 _2961_ (.A(net786),
    .B(_0555_),
    .C(_0556_),
    .Y(_0557_));
 sg13g2_o21ai_1 _2962_ (.B1(net615),
    .Y(_0558_),
    .A1(_0553_),
    .A2(_0557_));
 sg13g2_nand2b_1 _2963_ (.Y(_0559_),
    .B(net796),
    .A_N(net615));
 sg13g2_nand3_1 _2964_ (.B(_0558_),
    .C(_0559_),
    .A(net814),
    .Y(_0054_));
 sg13g2_mux2_1 _2965_ (.A0(_0886_),
    .A1(_0867_),
    .S(net620),
    .X(_0560_));
 sg13g2_xor2_1 _2966_ (.B(\logo_left[8] ),
    .A(net791),
    .X(_0561_));
 sg13g2_nor2_1 _2967_ (.A(_0542_),
    .B(_0554_),
    .Y(_0562_));
 sg13g2_o21ai_1 _2968_ (.B1(_0541_),
    .Y(_0563_),
    .A1(net791),
    .A2(_0882_));
 sg13g2_a221oi_1 _2969_ (.B2(_0562_),
    .C1(_0563_),
    .B1(_0543_),
    .A1(_0758_),
    .Y(_0564_),
    .A2(net796));
 sg13g2_nor2_1 _2970_ (.A(_0561_),
    .B(_0564_),
    .Y(_0565_));
 sg13g2_a21o_1 _2971_ (.A2(_0564_),
    .A1(_0561_),
    .B1(net786),
    .X(_0566_));
 sg13g2_o21ai_1 _2972_ (.B1(net617),
    .Y(_0567_),
    .A1(_0565_),
    .A2(_0566_));
 sg13g2_a21oi_1 _2973_ (.A1(net786),
    .A2(_0560_),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_o21ai_1 _2974_ (.B1(net814),
    .Y(_0569_),
    .A1(net256),
    .A2(net617));
 sg13g2_nor2_1 _2975_ (.A(_0568_),
    .B(_0569_),
    .Y(_0055_));
 sg13g2_a21oi_1 _2976_ (.A1(_0758_),
    .A2(\logo_left[8] ),
    .Y(_0570_),
    .B1(_0565_));
 sg13g2_xor2_1 _2977_ (.B(\logo_left[9] ),
    .A(net791),
    .X(_0571_));
 sg13g2_a21oi_1 _2978_ (.A1(_0570_),
    .A2(_0571_),
    .Y(_0572_),
    .B1(net786));
 sg13g2_o21ai_1 _2979_ (.B1(_0572_),
    .Y(_0573_),
    .A1(_0570_),
    .A2(_0571_));
 sg13g2_nand2_1 _2980_ (.Y(_0574_),
    .A(_0895_),
    .B(_0491_));
 sg13g2_and2_1 _2981_ (.A(net615),
    .B(_0574_),
    .X(_0575_));
 sg13g2_o21ai_1 _2982_ (.B1(net815),
    .Y(_0576_),
    .A1(net263),
    .A2(net615));
 sg13g2_a21oi_1 _2983_ (.A1(_0573_),
    .A2(_0575_),
    .Y(_0056_),
    .B1(_0576_));
 sg13g2_a22oi_1 _2984_ (.Y(_0577_),
    .B1(_0850_),
    .B2(_0852_),
    .A2(_0834_),
    .A1(_0833_));
 sg13g2_nand2b_1 _2985_ (.Y(_0578_),
    .B(_0849_),
    .A_N(_0577_));
 sg13g2_a22oi_1 _2986_ (.Y(_0579_),
    .B1(_0839_),
    .B2(_0578_),
    .A2(\logo_top[8] ),
    .A1(net793));
 sg13g2_nand4_1 _2987_ (.B(_0889_),
    .C(_0467_),
    .A(\gamepad.decoder.data_reg[6] ),
    .Y(_0580_),
    .D(_0579_));
 sg13g2_inv_1 _2988_ (.Y(_0581_),
    .A(net614));
 sg13g2_nand2_1 _2989_ (.Y(_0582_),
    .A(net194),
    .B(_0467_));
 sg13g2_nor2_1 _2990_ (.A(\logo_top[3] ),
    .B(\logo_top[2] ),
    .Y(_0583_));
 sg13g2_and2_1 _2991_ (.A(_0840_),
    .B(_0583_),
    .X(_0584_));
 sg13g2_nor2_1 _2992_ (.A(\logo_top[5] ),
    .B(\logo_top[4] ),
    .Y(_0585_));
 sg13g2_nand2_1 _2993_ (.Y(_0586_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_nor3_2 _2994_ (.A(net794),
    .B(\logo_top[6] ),
    .C(_0586_),
    .Y(_0587_));
 sg13g2_nor2_1 _2995_ (.A(net793),
    .B(\logo_top[8] ),
    .Y(_0588_));
 sg13g2_a21o_1 _2996_ (.A2(_0588_),
    .A1(_0587_),
    .B1(_0582_),
    .X(_0589_));
 sg13g2_nand3_1 _2997_ (.B(net614),
    .C(_0589_),
    .A(net786),
    .Y(_0590_));
 sg13g2_and2_1 _2998_ (.A(_0823_),
    .B(_0590_),
    .X(_0591_));
 sg13g2_nand2_2 _2999_ (.Y(_0592_),
    .A(_0823_),
    .B(_0590_));
 sg13g2_o21ai_1 _3000_ (.B1(net812),
    .Y(_0593_),
    .A1(\logo_top[0] ),
    .A2(net611));
 sg13g2_a21oi_1 _3001_ (.A1(_0763_),
    .A2(net611),
    .Y(_0057_),
    .B1(_0593_));
 sg13g2_a21oi_1 _3002_ (.A1(_0826_),
    .A2(_0841_),
    .Y(_0594_),
    .B1(_0580_));
 sg13g2_nand3_1 _3003_ (.B(_0841_),
    .C(_0580_),
    .A(_0826_),
    .Y(_0595_));
 sg13g2_nor2_1 _3004_ (.A(net781),
    .B(_0594_),
    .Y(_0596_));
 sg13g2_xor2_1 _3005_ (.B(net795),
    .A(net790),
    .X(_0597_));
 sg13g2_xnor2_1 _3006_ (.Y(_0598_),
    .A(_0763_),
    .B(_0597_));
 sg13g2_a221oi_1 _3007_ (.B2(net781),
    .C1(_0592_),
    .B1(_0598_),
    .A1(_0595_),
    .Y(_0599_),
    .A2(_0596_));
 sg13g2_o21ai_1 _3008_ (.B1(net812),
    .Y(_0600_),
    .A1(net795),
    .A2(net612));
 sg13g2_nor2_1 _3009_ (.A(_0599_),
    .B(_0600_),
    .Y(_0058_));
 sg13g2_xnor2_1 _3010_ (.Y(_0601_),
    .A(\logo_top[2] ),
    .B(_0826_));
 sg13g2_xnor2_1 _3011_ (.Y(_0602_),
    .A(_0011_),
    .B(_0841_));
 sg13g2_o21ai_1 _3012_ (.B1(net785),
    .Y(_0603_),
    .A1(net613),
    .A2(_0601_));
 sg13g2_a21oi_1 _3013_ (.A1(net613),
    .A2(_0602_),
    .Y(_0604_),
    .B1(_0603_));
 sg13g2_xnor2_1 _3014_ (.Y(_0605_),
    .A(net788),
    .B(\logo_top[2] ));
 sg13g2_a21oi_1 _3015_ (.A1(net789),
    .A2(_0826_),
    .Y(_0606_),
    .B1(_0840_));
 sg13g2_and2_1 _3016_ (.A(_0605_),
    .B(_0606_),
    .X(_0607_));
 sg13g2_o21ai_1 _3017_ (.B1(net781),
    .Y(_0608_),
    .A1(_0605_),
    .A2(_0606_));
 sg13g2_o21ai_1 _3018_ (.B1(net611),
    .Y(_0609_),
    .A1(_0607_),
    .A2(_0608_));
 sg13g2_o21ai_1 _3019_ (.B1(net815),
    .Y(_0610_),
    .A1(_0604_),
    .A2(_0609_));
 sg13g2_a21oi_1 _3020_ (.A1(_0762_),
    .A2(_0592_),
    .Y(_0059_),
    .B1(_0610_));
 sg13g2_o21ai_1 _3021_ (.B1(net785),
    .Y(_0611_),
    .A1(_0855_),
    .A2(net613));
 sg13g2_a21oi_1 _3022_ (.A1(_0843_),
    .A2(net613),
    .Y(_0612_),
    .B1(_0611_));
 sg13g2_xor2_1 _3023_ (.B(\logo_top[3] ),
    .A(net788),
    .X(_0613_));
 sg13g2_a21oi_1 _3024_ (.A1(_0757_),
    .A2(\logo_top[2] ),
    .Y(_0614_),
    .B1(_0607_));
 sg13g2_xnor2_1 _3025_ (.Y(_0615_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_nor2_1 _3026_ (.A(net787),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_o21ai_1 _3027_ (.B1(net611),
    .Y(_0617_),
    .A1(_0612_),
    .A2(_0616_));
 sg13g2_a21oi_1 _3028_ (.A1(net247),
    .A2(_0592_),
    .Y(_0618_),
    .B1(_0773_));
 sg13g2_nand2_1 _3029_ (.Y(_0060_),
    .A(_0617_),
    .B(_0618_));
 sg13g2_nand2_1 _3030_ (.Y(_0619_),
    .A(_0012_),
    .B(_0584_));
 sg13g2_xor2_1 _3031_ (.B(_0584_),
    .A(_0012_),
    .X(_0620_));
 sg13g2_or2_1 _3032_ (.X(_0621_),
    .B(net614),
    .A(_0853_));
 sg13g2_a21oi_1 _3033_ (.A1(net613),
    .A2(_0620_),
    .Y(_0622_),
    .B1(net781));
 sg13g2_nor2b_1 _3034_ (.A(net788),
    .B_N(\logo_top[4] ),
    .Y(_0623_));
 sg13g2_xnor2_1 _3035_ (.Y(_0624_),
    .A(net788),
    .B(\logo_top[4] ));
 sg13g2_o21ai_1 _3036_ (.B1(_0607_),
    .Y(_0625_),
    .A1(_0757_),
    .A2(\logo_top[3] ));
 sg13g2_o21ai_1 _3037_ (.B1(_0625_),
    .Y(_0626_),
    .A1(net788),
    .A2(_0583_));
 sg13g2_xor2_1 _3038_ (.B(_0626_),
    .A(_0624_),
    .X(_0627_));
 sg13g2_a221oi_1 _3039_ (.B2(net781),
    .C1(_0592_),
    .B1(_0627_),
    .A1(_0621_),
    .Y(_0628_),
    .A2(_0622_));
 sg13g2_o21ai_1 _3040_ (.B1(net815),
    .Y(_0629_),
    .A1(net251),
    .A2(net611));
 sg13g2_nor2_1 _3041_ (.A(_0628_),
    .B(_0629_),
    .Y(_0061_));
 sg13g2_xnor2_1 _3042_ (.Y(_0630_),
    .A(\logo_top[5] ),
    .B(_0619_));
 sg13g2_a21o_1 _3043_ (.A2(_0626_),
    .A1(_0624_),
    .B1(_0623_),
    .X(_0631_));
 sg13g2_xnor2_1 _3044_ (.Y(_0632_),
    .A(net788),
    .B(\logo_top[5] ));
 sg13g2_xnor2_1 _3045_ (.Y(_0633_),
    .A(_0631_),
    .B(_0632_));
 sg13g2_o21ai_1 _3046_ (.B1(net611),
    .Y(_0634_),
    .A1(net787),
    .A2(_0633_));
 sg13g2_o21ai_1 _3047_ (.B1(net785),
    .Y(_0635_),
    .A1(_0581_),
    .A2(_0630_));
 sg13g2_a21oi_1 _3048_ (.A1(_0852_),
    .A2(_0581_),
    .Y(_0636_),
    .B1(_0635_));
 sg13g2_o21ai_1 _3049_ (.B1(net815),
    .Y(_0637_),
    .A1(_0634_),
    .A2(_0636_));
 sg13g2_a21oi_1 _3050_ (.A1(_0760_),
    .A2(_0592_),
    .Y(_0062_),
    .B1(_0637_));
 sg13g2_nand3_1 _3051_ (.B(_0584_),
    .C(_0585_),
    .A(_0013_),
    .Y(_0638_));
 sg13g2_xnor2_1 _3052_ (.Y(_0639_),
    .A(_0013_),
    .B(_0586_));
 sg13g2_nor2_1 _3053_ (.A(_0832_),
    .B(net613),
    .Y(_0640_));
 sg13g2_a21oi_1 _3054_ (.A1(net613),
    .A2(_0639_),
    .Y(_0641_),
    .B1(_0640_));
 sg13g2_xor2_1 _3055_ (.B(\logo_top[6] ),
    .A(net788),
    .X(_0642_));
 sg13g2_or2_1 _3056_ (.X(_0643_),
    .B(_0585_),
    .A(net789));
 sg13g2_nand3_1 _3057_ (.B(_0626_),
    .C(_0632_),
    .A(_0624_),
    .Y(_0644_));
 sg13g2_nand3_1 _3058_ (.B(_0643_),
    .C(_0644_),
    .A(_0642_),
    .Y(_0645_));
 sg13g2_a21oi_1 _3059_ (.A1(_0643_),
    .A2(_0644_),
    .Y(_0646_),
    .B1(_0642_));
 sg13g2_nor2_1 _3060_ (.A(net785),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_a22oi_1 _3061_ (.Y(_0648_),
    .B1(_0645_),
    .B2(_0647_),
    .A2(_0641_),
    .A1(net785));
 sg13g2_a21oi_1 _3062_ (.A1(net255),
    .A2(_0592_),
    .Y(_0649_),
    .B1(net805));
 sg13g2_o21ai_1 _3063_ (.B1(_0649_),
    .Y(_0063_),
    .A1(_0592_),
    .A2(_0648_));
 sg13g2_xor2_1 _3064_ (.B(_0638_),
    .A(net794),
    .X(_0650_));
 sg13g2_o21ai_1 _3065_ (.B1(net787),
    .Y(_0651_),
    .A1(_0835_),
    .A2(net614));
 sg13g2_a21oi_1 _3066_ (.A1(net613),
    .A2(_0650_),
    .Y(_0652_),
    .B1(_0651_));
 sg13g2_xor2_1 _3067_ (.B(net794),
    .A(net788),
    .X(_0653_));
 sg13g2_a21oi_1 _3068_ (.A1(_0757_),
    .A2(\logo_top[6] ),
    .Y(_0654_),
    .B1(_0646_));
 sg13g2_xnor2_1 _3069_ (.Y(_0655_),
    .A(_0653_),
    .B(_0654_));
 sg13g2_nor2_1 _3070_ (.A(net785),
    .B(_0655_),
    .Y(_0656_));
 sg13g2_nand2_1 _3071_ (.Y(_0657_),
    .A(net794),
    .B(_0592_));
 sg13g2_o21ai_1 _3072_ (.B1(net611),
    .Y(_0658_),
    .A1(_0652_),
    .A2(_0656_));
 sg13g2_nand3_1 _3073_ (.B(_0657_),
    .C(_0658_),
    .A(net813),
    .Y(_0064_));
 sg13g2_nand2_1 _3074_ (.Y(_0659_),
    .A(_0014_),
    .B(_0587_));
 sg13g2_xnor2_1 _3075_ (.Y(_0660_),
    .A(_0793_),
    .B(_0587_));
 sg13g2_o21ai_1 _3076_ (.B1(net785),
    .Y(_0661_),
    .A1(_0848_),
    .A2(net614));
 sg13g2_a21o_1 _3077_ (.A2(_0660_),
    .A1(net614),
    .B1(_0661_),
    .X(_0662_));
 sg13g2_nand2_1 _3078_ (.Y(_0663_),
    .A(_0757_),
    .B(\logo_top[8] ));
 sg13g2_xnor2_1 _3079_ (.Y(_0664_),
    .A(net790),
    .B(\logo_top[8] ));
 sg13g2_nor3_1 _3080_ (.A(_0642_),
    .B(_0644_),
    .C(_0653_),
    .Y(_0665_));
 sg13g2_o21ai_1 _3081_ (.B1(_0757_),
    .Y(_0666_),
    .A1(net794),
    .A2(\logo_top[6] ));
 sg13g2_nand2_1 _3082_ (.Y(_0667_),
    .A(_0643_),
    .B(_0666_));
 sg13g2_o21ai_1 _3083_ (.B1(_0664_),
    .Y(_0668_),
    .A1(_0665_),
    .A2(_0667_));
 sg13g2_or3_1 _3084_ (.A(_0664_),
    .B(_0665_),
    .C(_0667_),
    .X(_0669_));
 sg13g2_nand3_1 _3085_ (.B(_0668_),
    .C(_0669_),
    .A(net780),
    .Y(_0670_));
 sg13g2_nand3_1 _3086_ (.B(_0662_),
    .C(_0670_),
    .A(net612),
    .Y(_0671_));
 sg13g2_o21ai_1 _3087_ (.B1(_0671_),
    .Y(_0672_),
    .A1(net248),
    .A2(net612));
 sg13g2_nor2_1 _3088_ (.A(net805),
    .B(_0672_),
    .Y(_0065_));
 sg13g2_and2_1 _3089_ (.A(_0663_),
    .B(_0668_),
    .X(_0673_));
 sg13g2_xor2_1 _3090_ (.B(net793),
    .A(net790),
    .X(_0674_));
 sg13g2_a21oi_1 _3091_ (.A1(_0673_),
    .A2(_0674_),
    .Y(_0675_),
    .B1(net787));
 sg13g2_o21ai_1 _3092_ (.B1(_0675_),
    .Y(_0676_),
    .A1(_0673_),
    .A2(_0674_));
 sg13g2_xnor2_1 _3093_ (.Y(_0677_),
    .A(net793),
    .B(_0659_));
 sg13g2_nand3_1 _3094_ (.B(net614),
    .C(_0677_),
    .A(net785),
    .Y(_0678_));
 sg13g2_nand3_1 _3095_ (.B(_0676_),
    .C(_0678_),
    .A(net612),
    .Y(_0679_));
 sg13g2_o21ai_1 _3096_ (.B1(net812),
    .Y(_0680_),
    .A1(net793),
    .A2(net611));
 sg13g2_nor2b_1 _3097_ (.A(_0680_),
    .B_N(_0679_),
    .Y(_0066_));
 sg13g2_o21ai_1 _3098_ (.B1(_0467_),
    .Y(_0681_),
    .A1(\gamepad.decoder.data_reg[5] ),
    .A2(\gamepad.decoder.data_reg[4] ));
 sg13g2_a21oi_1 _3099_ (.A1(_0901_),
    .A2(_0681_),
    .Y(_0682_),
    .B1(_0825_));
 sg13g2_nand2b_1 _3100_ (.Y(_0683_),
    .B(_0487_),
    .A_N(_0900_));
 sg13g2_nand3b_1 _3101_ (.B(_0682_),
    .C(_0683_),
    .Y(_0684_),
    .A_N(_0899_));
 sg13g2_o21ai_1 _3102_ (.B1(net814),
    .Y(_0685_),
    .A1(_0758_),
    .A2(_0682_));
 sg13g2_nand2b_1 _3103_ (.Y(_0067_),
    .B(_0684_),
    .A_N(_0685_));
 sg13g2_o21ai_1 _3104_ (.B1(_0467_),
    .Y(_0686_),
    .A1(net194),
    .A2(net209));
 sg13g2_a21oi_1 _3105_ (.A1(_0859_),
    .A2(_0686_),
    .Y(_0687_),
    .B1(_0825_));
 sg13g2_o21ai_1 _3106_ (.B1(_0858_),
    .Y(_0688_),
    .A1(_0847_),
    .A2(_0582_));
 sg13g2_o21ai_1 _3107_ (.B1(net812),
    .Y(_0689_),
    .A1(net790),
    .A2(_0687_));
 sg13g2_a21oi_1 _3108_ (.A1(_0687_),
    .A2(_0688_),
    .Y(_0068_),
    .B1(_0689_));
 sg13g2_or2_1 _3109_ (.X(_0690_),
    .B(_0468_),
    .A(gamepad_start_prev));
 sg13g2_o21ai_1 _3110_ (.B1(net814),
    .Y(_0691_),
    .A1(net135),
    .A2(_0690_));
 sg13g2_a21oi_1 _3111_ (.A1(net780),
    .A2(_0690_),
    .Y(_0069_),
    .B1(net136));
 sg13g2_mux2_1 _3112_ (.A0(net220),
    .A1(\color_index[0] ),
    .S(_0902_),
    .X(_0692_));
 sg13g2_and2_1 _3113_ (.A(net808),
    .B(net221),
    .X(_0070_));
 sg13g2_nand2_1 _3114_ (.Y(_0693_),
    .A(net215),
    .B(_0902_));
 sg13g2_o21ai_1 _3115_ (.B1(net808),
    .Y(_0694_),
    .A1(net215),
    .A2(\color_index[0] ));
 sg13g2_a21oi_1 _3116_ (.A1(_0913_),
    .A2(_0693_),
    .Y(_0071_),
    .B1(_0694_));
 sg13g2_nand2_1 _3117_ (.Y(_0695_),
    .A(net146),
    .B(_0902_));
 sg13g2_a21oi_1 _3118_ (.A1(_0909_),
    .A2(_0695_),
    .Y(_0072_),
    .B1(net805));
 sg13g2_nor2_1 _3119_ (.A(net810),
    .B(net190),
    .Y(_0696_));
 sg13g2_a21oi_1 _3120_ (.A1(_0768_),
    .A2(net809),
    .Y(_0073_),
    .B1(_0696_));
 sg13g2_mux2_1 _3121_ (.A0(net184),
    .A1(\pix_y[1] ),
    .S(net810),
    .X(_0074_));
 sg13g2_nor2_1 _3122_ (.A(net809),
    .B(net169),
    .Y(_0697_));
 sg13g2_a21oi_1 _3123_ (.A1(_0770_),
    .A2(net809),
    .Y(_0075_),
    .B1(_0697_));
 sg13g2_mux2_1 _3124_ (.A0(net176),
    .A1(net783),
    .S(net808),
    .X(_0076_));
 sg13g2_mux2_1 _3125_ (.A0(net174),
    .A1(\pix_y[4] ),
    .S(net808),
    .X(_0077_));
 sg13g2_nor2_1 _3126_ (.A(net808),
    .B(net165),
    .Y(_0698_));
 sg13g2_nand3_1 _3127_ (.B(net782),
    .C(\pix_y[9] ),
    .A(\pix_y[2] ),
    .Y(_0699_));
 sg13g2_o21ai_1 _3128_ (.B1(net1),
    .Y(_0700_),
    .A1(_0821_),
    .A2(_0699_));
 sg13g2_nand2_2 _3129_ (.Y(_0701_),
    .A(_0474_),
    .B(_0700_));
 sg13g2_a21oi_1 _3130_ (.A1(_0771_),
    .A2(net808),
    .Y(_0078_),
    .B1(_0698_));
 sg13g2_nor2_1 _3131_ (.A(net811),
    .B(net172),
    .Y(_0702_));
 sg13g2_a21oi_1 _3132_ (.A1(_0772_),
    .A2(net811),
    .Y(_0079_),
    .B1(_0702_));
 sg13g2_nor2_1 _3133_ (.A(net811),
    .B(net157),
    .Y(_0703_));
 sg13g2_a21oi_1 _3134_ (.A1(net811),
    .A2(_0775_),
    .Y(_0080_),
    .B1(_0703_));
 sg13g2_nor2_1 _3135_ (.A(net809),
    .B(net163),
    .Y(_0704_));
 sg13g2_a21oi_1 _3136_ (.A1(net809),
    .A2(_0774_),
    .Y(_0081_),
    .B1(_0704_));
 sg13g2_a21oi_1 _3137_ (.A1(net805),
    .A2(_0779_),
    .Y(_0082_),
    .B1(_0427_));
 sg13g2_nand2_1 _3138_ (.Y(_0705_),
    .A(net741),
    .B(_0444_));
 sg13g2_nor2_1 _3139_ (.A(net806),
    .B(_0445_),
    .Y(_0706_));
 sg13g2_a22oi_1 _3140_ (.Y(_0707_),
    .B1(_0705_),
    .B2(_0706_),
    .A2(net806),
    .A1(net156));
 sg13g2_nor4_1 _3141_ (.A(_1511_),
    .B(_0401_),
    .C(_0429_),
    .D(_0707_),
    .Y(_0083_));
 sg13g2_nand2b_1 _3142_ (.Y(_0708_),
    .B(net806),
    .A_N(net229));
 sg13g2_xnor2_1 _3143_ (.Y(_0709_),
    .A(_0445_),
    .B(_0446_));
 sg13g2_o21ai_1 _3144_ (.B1(_0708_),
    .Y(_0710_),
    .A1(net806),
    .A2(_0709_));
 sg13g2_nor4_1 _3145_ (.A(_1511_),
    .B(_0401_),
    .C(_0429_),
    .D(_0710_),
    .Y(_0084_));
 sg13g2_or3_1 _3146_ (.A(_0443_),
    .B(_0447_),
    .C(_0448_),
    .X(_0711_));
 sg13g2_nor2b_1 _3147_ (.A(net806),
    .B_N(_0449_),
    .Y(_0712_));
 sg13g2_a22oi_1 _3148_ (.Y(_0713_),
    .B1(_0711_),
    .B2(_0712_),
    .A2(net167),
    .A1(net806));
 sg13g2_nor4_1 _3149_ (.A(_1511_),
    .B(_0401_),
    .C(_0429_),
    .D(_0713_),
    .Y(_0085_));
 sg13g2_nand2b_1 _3150_ (.Y(_0714_),
    .B(net807),
    .A_N(net219));
 sg13g2_nand3_1 _3151_ (.B(_0449_),
    .C(_0450_),
    .A(_0440_),
    .Y(_0715_));
 sg13g2_nor2b_2 _3152_ (.A(_0451_),
    .B_N(_0715_),
    .Y(_0716_));
 sg13g2_o21ai_1 _3153_ (.B1(_0714_),
    .Y(_0717_),
    .A1(net807),
    .A2(_0716_));
 sg13g2_nor4_1 _3154_ (.A(_1511_),
    .B(_0401_),
    .C(_0429_),
    .D(_0717_),
    .Y(_0086_));
 sg13g2_nor2b_1 _3155_ (.A(\gamepad.driver.pmod_clk_prev ),
    .B_N(\gamepad.driver.pmod_clk_sync[1] ),
    .Y(_0718_));
 sg13g2_nor2_1 _3156_ (.A(net805),
    .B(net777),
    .Y(_0719_));
 sg13g2_a22oi_1 _3157_ (.Y(_0087_),
    .B1(net748),
    .B2(_0754_),
    .A2(net776),
    .A1(_0755_));
 sg13g2_a22oi_1 _3158_ (.Y(_0088_),
    .B1(net748),
    .B2(_0753_),
    .A2(net776),
    .A1(_0754_));
 sg13g2_a22oi_1 _3159_ (.Y(_0089_),
    .B1(net748),
    .B2(_0752_),
    .A2(net776),
    .A1(_0753_));
 sg13g2_a22oi_1 _3160_ (.Y(_0090_),
    .B1(net748),
    .B2(_0751_),
    .A2(net776),
    .A1(_0752_));
 sg13g2_a22oi_1 _3161_ (.Y(_0091_),
    .B1(net748),
    .B2(_0750_),
    .A2(net776),
    .A1(_0751_));
 sg13g2_a22oi_1 _3162_ (.Y(_0092_),
    .B1(net749),
    .B2(_0749_),
    .A2(net777),
    .A1(_0750_));
 sg13g2_a22oi_1 _3163_ (.Y(_0093_),
    .B1(net749),
    .B2(_0748_),
    .A2(net777),
    .A1(_0749_));
 sg13g2_a22oi_1 _3164_ (.Y(_0094_),
    .B1(net749),
    .B2(_0747_),
    .A2(net777),
    .A1(_0748_));
 sg13g2_a22oi_1 _3165_ (.Y(_0095_),
    .B1(net749),
    .B2(_0746_),
    .A2(net777),
    .A1(_0747_));
 sg13g2_a22oi_1 _3166_ (.Y(_0096_),
    .B1(net748),
    .B2(_0745_),
    .A2(net776),
    .A1(_0746_));
 sg13g2_a22oi_1 _3167_ (.Y(_0097_),
    .B1(net748),
    .B2(_0744_),
    .A2(net776),
    .A1(_0745_));
 sg13g2_a22oi_1 _3168_ (.Y(_0098_),
    .B1(net748),
    .B2(_0767_),
    .A2(net776),
    .A1(_0744_));
 sg13g2_and2_1 _3169_ (.A(net813),
    .B(net5),
    .X(_0099_));
 sg13g2_and2_1 _3170_ (.A(net812),
    .B(net131),
    .X(_0100_));
 sg13g2_and2_1 _3171_ (.A(net812),
    .B(net4),
    .X(_0101_));
 sg13g2_and2_1 _3172_ (.A(net812),
    .B(net132),
    .X(_0102_));
 sg13g2_and2_1 _3173_ (.A(net812),
    .B(net3),
    .X(_0103_));
 sg13g2_and2_1 _3174_ (.A(net813),
    .B(net130),
    .X(_0104_));
 sg13g2_or2_1 _3175_ (.X(_0720_),
    .B(net654),
    .A(_0768_));
 sg13g2_nand2_1 _3176_ (.Y(_0721_),
    .A(net128),
    .B(_0473_));
 sg13g2_o21ai_1 _3177_ (.B1(_0720_),
    .Y(_0105_),
    .A1(_0700_),
    .A2(net129));
 sg13g2_a21oi_1 _3178_ (.A1(\pix_y[0] ),
    .A2(_0473_),
    .Y(_0722_),
    .B1(net239));
 sg13g2_nand3_1 _3179_ (.B(\pix_y[1] ),
    .C(_0473_),
    .A(\pix_y[0] ),
    .Y(_0723_));
 sg13g2_nand2_1 _3180_ (.Y(_0724_),
    .A(net810),
    .B(_0723_));
 sg13g2_nor2_1 _3181_ (.A(net240),
    .B(_0724_),
    .Y(_0106_));
 sg13g2_nand3_1 _3182_ (.B(net239),
    .C(net654),
    .A(net244),
    .Y(_0725_));
 sg13g2_or2_1 _3183_ (.X(_0726_),
    .B(_0725_),
    .A(_0770_));
 sg13g2_inv_1 _3184_ (.Y(_0727_),
    .A(_0726_));
 sg13g2_nand2_1 _3185_ (.Y(_0728_),
    .A(_0701_),
    .B(_0726_));
 sg13g2_a21oi_1 _3186_ (.A1(_0770_),
    .A2(_0725_),
    .Y(_0107_),
    .B1(_0728_));
 sg13g2_nand3_1 _3187_ (.B(_0701_),
    .C(_0726_),
    .A(net782),
    .Y(_0729_));
 sg13g2_or3_1 _3188_ (.A(_0770_),
    .B(net805),
    .C(_0723_),
    .X(_0730_));
 sg13g2_o21ai_1 _3189_ (.B1(_0729_),
    .Y(_0108_),
    .A1(net782),
    .A2(_0730_));
 sg13g2_nand2_1 _3190_ (.Y(_0731_),
    .A(net782),
    .B(\pix_y[4] ));
 sg13g2_or2_2 _3191_ (.X(_0732_),
    .B(_0731_),
    .A(_0726_));
 sg13g2_nand2_1 _3192_ (.Y(_0733_),
    .A(_0701_),
    .B(_0732_));
 sg13g2_a21oi_1 _3193_ (.A1(net782),
    .A2(_0727_),
    .Y(_0734_),
    .B1(net241));
 sg13g2_nor2_1 _3194_ (.A(_0733_),
    .B(_0734_),
    .Y(_0109_));
 sg13g2_nor2_1 _3195_ (.A(_0700_),
    .B(_0732_),
    .Y(_0735_));
 sg13g2_nor2_1 _3196_ (.A(net236),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_a21oi_1 _3197_ (.A1(net236),
    .A2(_0733_),
    .Y(_0110_),
    .B1(_0736_));
 sg13g2_o21ai_1 _3198_ (.B1(_0772_),
    .Y(_0737_),
    .A1(_0771_),
    .A2(_0732_));
 sg13g2_o21ai_1 _3199_ (.B1(_0701_),
    .Y(_0738_),
    .A1(_0795_),
    .A2(_0732_));
 sg13g2_nor2b_1 _3200_ (.A(_0738_),
    .B_N(_0737_),
    .Y(_0111_));
 sg13g2_or4_1 _3201_ (.A(net231),
    .B(_0795_),
    .C(_0730_),
    .D(_0731_),
    .X(_0739_));
 sg13g2_o21ai_1 _3202_ (.B1(_0739_),
    .Y(_0112_),
    .A1(_0775_),
    .A2(_0738_));
 sg13g2_o21ai_1 _3203_ (.B1(_0733_),
    .Y(_0740_),
    .A1(_0798_),
    .A2(_0700_));
 sg13g2_o21ai_1 _3204_ (.B1(_0774_),
    .Y(_0741_),
    .A1(_0796_),
    .A2(_0732_));
 sg13g2_nand2_1 _3205_ (.Y(_0742_),
    .A(_0740_),
    .B(net262));
 sg13g2_inv_1 _3206_ (.Y(_0113_),
    .A(_0742_));
 sg13g2_a22oi_1 _3207_ (.Y(_0743_),
    .B1(_0740_),
    .B2(net230),
    .A2(_0735_),
    .A1(_0799_));
 sg13g2_inv_1 _3208_ (.Y(_0114_),
    .A(_0743_));
 sg13g2_a21o_1 _3209_ (.A2(_0914_),
    .A1(net808),
    .B1(_0116_),
    .X(_0115_));
 sg13g2_dfrbp_1 _3210_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net87),
    .D(_0022_),
    .Q_N(_1596_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _3211_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net97),
    .D(_0023_),
    .Q_N(_1595_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _3212_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net96),
    .D(net143),
    .Q_N(_1594_),
    .Q(\gamepad.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _3213_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net94),
    .D(net151),
    .Q_N(_1593_),
    .Q(\gamepad.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net92),
    .D(net149),
    .Q_N(_1592_),
    .Q(\gamepad.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net90),
    .D(net141),
    .Q_N(_1591_),
    .Q(\gamepad.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net86),
    .D(net199),
    .Q_N(_1590_),
    .Q(\gamepad.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net84),
    .D(_0029_),
    .Q_N(_1589_),
    .Q(\gamepad.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net82),
    .D(_0030_),
    .Q_N(_1588_),
    .Q(\gamepad.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net80),
    .D(net195),
    .Q_N(_1587_),
    .Q(\gamepad.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net78),
    .D(net183),
    .Q_N(_1586_),
    .Q(\gamepad.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net76),
    .D(net162),
    .Q_N(_1585_),
    .Q(\gamepad.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(net155),
    .Q_N(_1584_),
    .Q(\gamepad.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net72),
    .D(net145),
    .Q_N(_1583_),
    .Q(\gamepad.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _3224_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net70),
    .D(net153),
    .Q_N(_1582_),
    .Q(gamepad_start_prev));
 sg13g2_dfrbp_1 _3225_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net68),
    .D(_0037_),
    .Q_N(_0021_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _3226_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net67),
    .D(_0038_),
    .Q_N(_1581_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _3227_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net66),
    .D(net213),
    .Q_N(_1580_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _3228_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net65),
    .D(_0040_),
    .Q_N(_1579_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _3229_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net64),
    .D(_0041_),
    .Q_N(_1578_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _3230_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net63),
    .D(_0042_),
    .Q_N(_1577_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _3231_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net62),
    .D(_0043_),
    .Q_N(_1576_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _3232_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net61),
    .D(_0044_),
    .Q_N(_1575_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net60),
    .D(_0045_),
    .Q_N(_1574_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net59),
    .D(_0046_),
    .Q_N(_1573_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net58),
    .D(net134),
    .Q_N(_0020_),
    .Q(\logo_left[0] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net56),
    .D(_0048_),
    .Q_N(_1572_),
    .Q(\logo_left[1] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net54),
    .D(_0049_),
    .Q_N(_0007_),
    .Q(\logo_left[2] ));
 sg13g2_dfrbp_1 _3238_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(_0050_),
    .Q_N(_1571_),
    .Q(\logo_left[3] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net50),
    .D(net259),
    .Q_N(_0008_),
    .Q(\logo_left[4] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net48),
    .D(_0052_),
    .Q_N(_1570_),
    .Q(\logo_left[5] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net46),
    .D(_0053_),
    .Q_N(_0009_),
    .Q(\logo_left[6] ));
 sg13g2_dfrbp_1 _3242_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net44),
    .D(_0054_),
    .Q_N(_1569_),
    .Q(\logo_left[7] ));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net42),
    .D(_0055_),
    .Q_N(_0010_),
    .Q(\logo_left[8] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net40),
    .D(_0056_),
    .Q_N(_1568_),
    .Q(\logo_left[9] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net38),
    .D(net139),
    .Q_N(_0019_),
    .Q(\logo_top[0] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net36),
    .D(_0058_),
    .Q_N(_1567_),
    .Q(\logo_top[1] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net34),
    .D(_0059_),
    .Q_N(_0011_),
    .Q(\logo_top[2] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net32),
    .D(_0060_),
    .Q_N(_1566_),
    .Q(\logo_top[3] ));
 sg13g2_dfrbp_1 _3249_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net30),
    .D(_0061_),
    .Q_N(_0012_),
    .Q(\logo_top[4] ));
 sg13g2_dfrbp_1 _3250_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net28),
    .D(_0062_),
    .Q_N(_1565_),
    .Q(\logo_top[5] ));
 sg13g2_dfrbp_1 _3251_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net26),
    .D(_0063_),
    .Q_N(_0013_),
    .Q(\logo_top[6] ));
 sg13g2_dfrbp_1 _3252_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net24),
    .D(_0064_),
    .Q_N(_1564_),
    .Q(\logo_top[7] ));
 sg13g2_dfrbp_1 _3253_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net22),
    .D(_0065_),
    .Q_N(_0014_),
    .Q(\logo_top[8] ));
 sg13g2_dfrbp_1 _3254_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net119),
    .D(_0066_),
    .Q_N(_1563_),
    .Q(\logo_top[9] ));
 sg13g2_dfrbp_1 _3255_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net116),
    .D(_0067_),
    .Q_N(_1562_),
    .Q(dir_x));
 sg13g2_dfrbp_1 _3256_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net114),
    .D(_0068_),
    .Q_N(_1561_),
    .Q(dir_y));
 sg13g2_dfrbp_1 _3257_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net112),
    .D(net137),
    .Q_N(_0004_),
    .Q(manual_mode));
 sg13g2_dfrbp_1 _3258_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net110),
    .D(_0070_),
    .Q_N(_0018_),
    .Q(\color_index[0] ));
 sg13g2_dfrbp_1 _3259_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net108),
    .D(net216),
    .Q_N(_0016_),
    .Q(\color_index[1] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net105),
    .D(net147),
    .Q_N(_0015_),
    .Q(\color_index[2] ));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net103),
    .D(net191),
    .Q_N(_1560_),
    .Q(\prev_y[0] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net102),
    .D(net185),
    .Q_N(_1559_),
    .Q(\prev_y[1] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net101),
    .D(net170),
    .Q_N(_1558_),
    .Q(\prev_y[2] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net100),
    .D(net177),
    .Q_N(_1557_),
    .Q(\prev_y[3] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net99),
    .D(net175),
    .Q_N(_1556_),
    .Q(\prev_y[4] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net98),
    .D(net166),
    .Q_N(_1555_),
    .Q(\prev_y[5] ));
 sg13g2_dfrbp_1 _3267_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net95),
    .D(net173),
    .Q_N(_1554_),
    .Q(\prev_y[6] ));
 sg13g2_dfrbp_1 _3268_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net93),
    .D(net158),
    .Q_N(_1553_),
    .Q(\prev_y[7] ));
 sg13g2_dfrbp_1 _3269_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net91),
    .D(net164),
    .Q_N(_1552_),
    .Q(\prev_y[8] ));
 sg13g2_dfrbp_1 _3270_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net89),
    .D(net160),
    .Q_N(_1551_),
    .Q(\prev_y[9] ));
 sg13g2_dfrbp_1 _3271_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net85),
    .D(_0083_),
    .Q_N(_1550_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _3272_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net83),
    .D(_0084_),
    .Q_N(_1549_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _3273_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(_0085_),
    .Q_N(_1548_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _3274_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net88),
    .D(_0086_),
    .Q_N(_1597_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _3275_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net107),
    .D(net126),
    .Q_N(_1598_),
    .Q(\gamepad.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _3276_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net79),
    .D(net125),
    .Q_N(_1547_),
    .Q(\gamepad.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _3277_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net77),
    .D(net203),
    .Q_N(_1546_),
    .Q(\gamepad.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _3278_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net73),
    .D(_0088_),
    .Q_N(_1545_),
    .Q(\gamepad.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _3279_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net69),
    .D(net201),
    .Q_N(_1544_),
    .Q(\gamepad.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _3280_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net55),
    .D(net181),
    .Q_N(_1543_),
    .Q(\gamepad.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _3281_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net51),
    .D(_0091_),
    .Q_N(_1542_),
    .Q(\gamepad.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _3282_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net47),
    .D(net189),
    .Q_N(_1541_),
    .Q(\gamepad.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _3283_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net43),
    .D(net193),
    .Q_N(_1540_),
    .Q(\gamepad.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _3284_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net39),
    .D(net208),
    .Q_N(_1539_),
    .Q(\gamepad.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _3285_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net35),
    .D(net205),
    .Q_N(_1538_),
    .Q(\gamepad.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _3286_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net31),
    .D(net197),
    .Q_N(_1537_),
    .Q(\gamepad.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _3287_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net27),
    .D(net187),
    .Q_N(_1536_),
    .Q(\gamepad.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _3288_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net23),
    .D(net179),
    .Q_N(_1535_),
    .Q(\gamepad.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _3289_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net117),
    .D(_0099_),
    .Q_N(_1534_),
    .Q(\gamepad.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _3290_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net115),
    .D(_0100_),
    .Q_N(_1533_),
    .Q(\gamepad.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _3291_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net113),
    .D(_0101_),
    .Q_N(_1532_),
    .Q(\gamepad.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _3292_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net111),
    .D(_0102_),
    .Q_N(_1531_),
    .Q(\gamepad.driver.pmod_clk_sync[1] ));
 sg13g2_dfrbp_1 _3293_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net109),
    .D(_0103_),
    .Q_N(_1530_),
    .Q(\gamepad.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _3294_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net118),
    .D(_0104_),
    .Q_N(_1599_),
    .Q(\gamepad.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _3295_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net106),
    .D(net226),
    .Q_N(_1529_),
    .Q(hsync));
 sg13g2_dfrbp_1 _3296_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net104),
    .D(_0105_),
    .Q_N(_0017_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _3297_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net71),
    .D(_0106_),
    .Q_N(_1528_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _3298_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net53),
    .D(net245),
    .Q_N(_1527_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _3299_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net45),
    .D(_0108_),
    .Q_N(_1526_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _3300_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net37),
    .D(_0109_),
    .Q_N(_1525_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _3301_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net29),
    .D(_0110_),
    .Q_N(_1524_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _3302_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net124),
    .D(_0111_),
    .Q_N(_1523_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _3303_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net57),
    .D(net232),
    .Q_N(_1522_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _3304_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net41),
    .D(_0113_),
    .Q_N(_1521_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _3305_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net120),
    .D(_0114_),
    .Q_N(_1600_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _3306_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net25),
    .D(net238),
    .Q_N(_1520_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _3307_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net121),
    .D(_0115_),
    .Q_N(_1601_),
    .Q(\palette_inst.rrggbb[5] ));
 sg13g2_dfrbp_1 _3308_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net122),
    .D(_0000_),
    .Q_N(_1602_),
    .Q(\palette_inst.rrggbb[0] ));
 sg13g2_dfrbp_1 _3309_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net123),
    .D(_0001_),
    .Q_N(_1603_),
    .Q(\palette_inst.rrggbb[1] ));
 sg13g2_dfrbp_1 _3310_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net75),
    .D(_0002_),
    .Q_N(_1604_),
    .Q(\palette_inst.rrggbb[2] ));
 sg13g2_dfrbp_1 _3311_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net49),
    .D(_0003_),
    .Q_N(_1519_),
    .Q(\palette_inst.rrggbb[3] ));
 sg13g2_dfrbp_1 _3312_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net33),
    .D(_0116_),
    .Q_N(_1518_),
    .Q(\palette_inst.rrggbb[4] ));
 sg13g2_tiehi _3288__23 (.L_HI(net23));
 sg13g2_tiehi _3252__24 (.L_HI(net24));
 sg13g2_tiehi _3306__25 (.L_HI(net25));
 sg13g2_tiehi _3251__26 (.L_HI(net26));
 sg13g2_tiehi _3287__27 (.L_HI(net27));
 sg13g2_tiehi _3250__28 (.L_HI(net28));
 sg13g2_tiehi _3301__29 (.L_HI(net29));
 sg13g2_tiehi _3249__30 (.L_HI(net30));
 sg13g2_tiehi _3286__31 (.L_HI(net31));
 sg13g2_tiehi _3248__32 (.L_HI(net32));
 sg13g2_tiehi _3312__33 (.L_HI(net33));
 sg13g2_tiehi _3247__34 (.L_HI(net34));
 sg13g2_tiehi _3285__35 (.L_HI(net35));
 sg13g2_tiehi _3246__36 (.L_HI(net36));
 sg13g2_tiehi _3300__37 (.L_HI(net37));
 sg13g2_tiehi _3245__38 (.L_HI(net38));
 sg13g2_tiehi _3284__39 (.L_HI(net39));
 sg13g2_tiehi _3244__40 (.L_HI(net40));
 sg13g2_tiehi _3304__41 (.L_HI(net41));
 sg13g2_tiehi _3243__42 (.L_HI(net42));
 sg13g2_tiehi _3283__43 (.L_HI(net43));
 sg13g2_tiehi _3242__44 (.L_HI(net44));
 sg13g2_tiehi _3299__45 (.L_HI(net45));
 sg13g2_tiehi _3241__46 (.L_HI(net46));
 sg13g2_tiehi _3282__47 (.L_HI(net47));
 sg13g2_tiehi _3240__48 (.L_HI(net48));
 sg13g2_tiehi _3311__49 (.L_HI(net49));
 sg13g2_tiehi _3239__50 (.L_HI(net50));
 sg13g2_tiehi _3281__51 (.L_HI(net51));
 sg13g2_tiehi _3238__52 (.L_HI(net52));
 sg13g2_tiehi _3298__53 (.L_HI(net53));
 sg13g2_tiehi _3237__54 (.L_HI(net54));
 sg13g2_tiehi _3280__55 (.L_HI(net55));
 sg13g2_tiehi _3236__56 (.L_HI(net56));
 sg13g2_tiehi _3303__57 (.L_HI(net57));
 sg13g2_tiehi _3235__58 (.L_HI(net58));
 sg13g2_tiehi _3234__59 (.L_HI(net59));
 sg13g2_tiehi _3233__60 (.L_HI(net60));
 sg13g2_tiehi _3232__61 (.L_HI(net61));
 sg13g2_tiehi _3231__62 (.L_HI(net62));
 sg13g2_tiehi _3230__63 (.L_HI(net63));
 sg13g2_tiehi _3229__64 (.L_HI(net64));
 sg13g2_tiehi _3228__65 (.L_HI(net65));
 sg13g2_tiehi _3227__66 (.L_HI(net66));
 sg13g2_tiehi _3226__67 (.L_HI(net67));
 sg13g2_tiehi _3225__68 (.L_HI(net68));
 sg13g2_tiehi _3279__69 (.L_HI(net69));
 sg13g2_tiehi _3224__70 (.L_HI(net70));
 sg13g2_tiehi _3297__71 (.L_HI(net71));
 sg13g2_tiehi _3223__72 (.L_HI(net72));
 sg13g2_tiehi _3278__73 (.L_HI(net73));
 sg13g2_tiehi _3222__74 (.L_HI(net74));
 sg13g2_tiehi _3310__75 (.L_HI(net75));
 sg13g2_tiehi _3221__76 (.L_HI(net76));
 sg13g2_tiehi _3277__77 (.L_HI(net77));
 sg13g2_tiehi _3220__78 (.L_HI(net78));
 sg13g2_tiehi _3276__79 (.L_HI(net79));
 sg13g2_tiehi _3219__80 (.L_HI(net80));
 sg13g2_tiehi _3273__81 (.L_HI(net81));
 sg13g2_tiehi _3218__82 (.L_HI(net82));
 sg13g2_tiehi _3272__83 (.L_HI(net83));
 sg13g2_tiehi _3217__84 (.L_HI(net84));
 sg13g2_tiehi _3271__85 (.L_HI(net85));
 sg13g2_tiehi _3216__86 (.L_HI(net86));
 sg13g2_tiehi _3210__87 (.L_HI(net87));
 sg13g2_tiehi _3274__88 (.L_HI(net88));
 sg13g2_tiehi _3270__89 (.L_HI(net89));
 sg13g2_tiehi _3215__90 (.L_HI(net90));
 sg13g2_tiehi _3269__91 (.L_HI(net91));
 sg13g2_tiehi _3214__92 (.L_HI(net92));
 sg13g2_tiehi _3268__93 (.L_HI(net93));
 sg13g2_tiehi _3213__94 (.L_HI(net94));
 sg13g2_tiehi _3267__95 (.L_HI(net95));
 sg13g2_tiehi _3212__96 (.L_HI(net96));
 sg13g2_tiehi _3211__97 (.L_HI(net97));
 sg13g2_tiehi _3266__98 (.L_HI(net98));
 sg13g2_tiehi _3265__99 (.L_HI(net99));
 sg13g2_tiehi _3264__100 (.L_HI(net100));
 sg13g2_tiehi _3263__101 (.L_HI(net101));
 sg13g2_tiehi _3262__102 (.L_HI(net102));
 sg13g2_tiehi _3261__103 (.L_HI(net103));
 sg13g2_tiehi _3296__104 (.L_HI(net104));
 sg13g2_tiehi _3260__105 (.L_HI(net105));
 sg13g2_tiehi _3295__106 (.L_HI(net106));
 sg13g2_tiehi _3275__107 (.L_HI(net107));
 sg13g2_tiehi _3259__108 (.L_HI(net108));
 sg13g2_tiehi _3293__109 (.L_HI(net109));
 sg13g2_tiehi _3258__110 (.L_HI(net110));
 sg13g2_tiehi _3292__111 (.L_HI(net111));
 sg13g2_tiehi _3257__112 (.L_HI(net112));
 sg13g2_tiehi _3291__113 (.L_HI(net113));
 sg13g2_tiehi _3256__114 (.L_HI(net114));
 sg13g2_tiehi _3290__115 (.L_HI(net115));
 sg13g2_tiehi _3255__116 (.L_HI(net116));
 sg13g2_tiehi _3289__117 (.L_HI(net117));
 sg13g2_tiehi _3294__118 (.L_HI(net118));
 sg13g2_tiehi _3254__119 (.L_HI(net119));
 sg13g2_tiehi _3305__120 (.L_HI(net120));
 sg13g2_tiehi _3307__121 (.L_HI(net121));
 sg13g2_tiehi _3308__122 (.L_HI(net122));
 sg13g2_tiehi _3309__123 (.L_HI(net123));
 sg13g2_tiehi _3302__124 (.L_HI(net124));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_7 (.L_LO(net7));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_8 (.L_LO(net8));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_9 (.L_LO(net9));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_10 (.L_LO(net10));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_11 (.L_LO(net11));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_12 (.L_LO(net12));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_13 (.L_LO(net13));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_14 (.L_LO(net14));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_15 (.L_LO(net15));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_16 (.L_LO(net16));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_17 (.L_LO(net17));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_18 (.L_LO(net18));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_19 (.L_LO(net19));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_20 (.L_LO(net20));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_21 (.L_LO(net21));
 sg13g2_tiehi _3253__22 (.L_HI(net22));
 sg13g2_buf_1 _3432_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _3433_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(_0591_));
 sg13g2_buf_2 fanout612 (.A(_0591_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_0580_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net617),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_0492_),
    .X(net616));
 sg13g2_buf_1 fanout617 (.A(_0492_),
    .X(net617));
 sg13g2_buf_4 fanout618 (.X(net618),
    .A(_1102_));
 sg13g2_buf_1 fanout619 (.A(_1102_),
    .X(net619));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(_0490_));
 sg13g2_buf_2 fanout621 (.A(_0490_),
    .X(net621));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(_1243_));
 sg13g2_buf_2 fanout623 (.A(_1210_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_1304_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_1207_),
    .X(net625));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(_1206_));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(_1123_));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(_1107_));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(_1074_));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(net632));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(net632));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(_1073_));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(_1063_));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(_1062_));
 sg13g2_buf_4 fanout636 (.X(net636),
    .A(_1062_));
 sg13g2_buf_4 fanout637 (.X(net637),
    .A(_1033_));
 sg13g2_buf_2 fanout638 (.A(_1008_),
    .X(net638));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(_1006_));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(net642));
 sg13g2_buf_2 fanout642 (.A(_0994_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_0984_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_0981_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_0981_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(net651),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_0980_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_0980_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_0474_),
    .X(net654));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(_1295_));
 sg13g2_buf_2 fanout656 (.A(_1075_),
    .X(net656));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(net659));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net659));
 sg13g2_buf_4 fanout659 (.X(net659),
    .A(_1052_));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(net661));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(_1051_));
 sg13g2_buf_2 fanout662 (.A(net665),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net665),
    .X(net663));
 sg13g2_buf_4 fanout664 (.X(net664),
    .A(net665));
 sg13g2_buf_2 fanout665 (.A(_1042_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(_1041_));
 sg13g2_buf_2 fanout668 (.A(net669),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_1041_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_1023_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_1023_),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(_1022_));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(_1022_));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(_1020_));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_1002_));
 sg13g2_buf_2 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_1001_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_0979_),
    .X(net678));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_0979_));
 sg13g2_buf_2 fanout680 (.A(_0978_),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_0978_));
 sg13g2_buf_2 fanout682 (.A(_0977_),
    .X(net682));
 sg13g2_buf_1 fanout683 (.A(_0977_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_0977_),
    .X(net684));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(_0976_));
 sg13g2_buf_2 fanout686 (.A(net689),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net689),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_0975_),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(_0974_));
 sg13g2_buf_2 fanout691 (.A(_0964_),
    .X(net691));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(net693));
 sg13g2_buf_2 fanout693 (.A(net694),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(net697),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_0955_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_1 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_0954_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net704),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net704),
    .X(net703));
 sg13g2_buf_1 fanout704 (.A(_0954_),
    .X(net704));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(_0933_));
 sg13g2_buf_1 fanout706 (.A(_0933_),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_1024_));
 sg13g2_buf_2 fanout708 (.A(net709),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_0961_),
    .X(net709));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(_0961_));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(net712));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(_0960_));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_0958_));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(_0958_));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(_0957_));
 sg13g2_buf_2 fanout716 (.A(_0957_),
    .X(net716));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(net718));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(_0930_));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(net722));
 sg13g2_buf_2 fanout720 (.A(net722),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_0930_),
    .X(net722));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(net727));
 sg13g2_buf_2 fanout724 (.A(net727),
    .X(net724));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(net727));
 sg13g2_buf_2 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_0929_),
    .X(net727));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(_1043_));
 sg13g2_buf_2 fanout729 (.A(_1043_),
    .X(net729));
 sg13g2_buf_4 fanout730 (.X(net730),
    .A(net731));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(_1000_));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(_0999_));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(_0999_));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(net736));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net736));
 sg13g2_buf_2 fanout736 (.A(_0993_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(net739),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(_0992_));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net741));
 sg13g2_buf_2 fanout741 (.A(_0932_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(_0932_));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(net747));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(net747));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_0931_),
    .X(net747));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(_0719_));
 sg13g2_buf_2 fanout749 (.A(_0719_),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(_0462_));
 sg13g2_buf_2 fanout751 (.A(_0462_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(net754),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_0991_),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(_0991_));
 sg13g2_buf_2 fanout756 (.A(_0991_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(net759),
    .X(net757));
 sg13g2_buf_1 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(_0990_));
 sg13g2_buf_2 fanout760 (.A(net762),
    .X(net760));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(_0990_));
 sg13g2_buf_1 fanout762 (.A(_0990_),
    .X(net762));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(net765));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(net769));
 sg13g2_buf_2 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_4 fanout767 (.X(net767),
    .A(net768));
 sg13g2_buf_1 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_0988_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(net775),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(net774));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(net775));
 sg13g2_buf_2 fanout775 (.A(_0987_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_0718_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_0718_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_0461_),
    .X(net778));
 sg13g2_buf_1 fanout779 (.A(_0461_),
    .X(net779));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(_0756_));
 sg13g2_buf_1 fanout781 (.A(_0756_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(net237),
    .X(net783));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(net787));
 sg13g2_buf_2 fanout785 (.A(net786),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(manual_mode),
    .X(net787));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(net790));
 sg13g2_buf_1 fanout789 (.A(net790),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net253));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(net792));
 sg13g2_buf_2 fanout792 (.A(dir_x),
    .X(net792));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(net257));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(net265));
 sg13g2_buf_2 fanout795 (.A(net254),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net271),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(net266));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(net264));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(\logo_left[4] ));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net270));
 sg13g2_buf_2 fanout801 (.A(net267),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_1 fanout803 (.A(\logo_left[1] ),
    .X(net803));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(\logo_left[0] ));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_0773_));
 sg13g2_buf_2 fanout806 (.A(net807),
    .X(net806));
 sg13g2_buf_1 fanout807 (.A(ui_in[1]),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net811));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(net1));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_1 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(net815),
    .X(net814));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_tielo tt_um_zerotoasic_logo_screensaver_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad.driver.pmod_latch_sync[1] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad.driver.pmod_clk_sync[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0021_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0017_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0721_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold6 (.A(\gamepad.driver.pmod_latch_sync[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold7 (.A(\gamepad.driver.pmod_data_sync[0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold8 (.A(\gamepad.driver.pmod_clk_sync[0] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0020_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0047_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0004_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0691_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0069_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0019_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0057_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold16 (.A(\gamepad.decoder.data_reg[3] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0027_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold18 (.A(\gamepad.decoder.data_reg[0] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0024_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold20 (.A(\gamepad.decoder.data_reg[11] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0035_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold22 (.A(\color_index[2] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0072_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold24 (.A(\gamepad.decoder.data_reg[2] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0026_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold26 (.A(\gamepad.decoder.data_reg[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0025_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold28 (.A(gamepad_start_prev),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0036_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold30 (.A(\gamepad.decoder.data_reg[10] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0034_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold32 (.A(\palette_inst.rrggbb[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold33 (.A(\prev_y[7] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0080_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold35 (.A(\prev_y[9] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0082_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold37 (.A(\gamepad.decoder.data_reg[9] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0033_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold39 (.A(\prev_y[8] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0081_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold41 (.A(\prev_y[5] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0078_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold43 (.A(\palette_inst.rrggbb[2] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold44 (.A(\palette_inst.rrggbb[5] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold45 (.A(\prev_y[2] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0075_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold47 (.A(\palette_inst.rrggbb[4] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold48 (.A(\prev_y[6] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0079_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold50 (.A(\prev_y[4] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0077_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold52 (.A(\prev_y[3] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0076_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold54 (.A(\gamepad.driver.shift_reg[11] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0098_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold56 (.A(\gamepad.driver.shift_reg[3] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0090_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold58 (.A(\gamepad.decoder.data_reg[8] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0032_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold60 (.A(\prev_y[1] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0074_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold62 (.A(\gamepad.driver.shift_reg[10] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0097_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold64 (.A(\gamepad.driver.shift_reg[5] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0092_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold66 (.A(\prev_y[0] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0073_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold68 (.A(\gamepad.driver.shift_reg[6] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0093_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold70 (.A(\gamepad.decoder.data_reg[7] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0031_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold72 (.A(\gamepad.driver.shift_reg[9] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0096_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold74 (.A(\gamepad.decoder.data_reg[4] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0028_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold76 (.A(\gamepad.driver.shift_reg[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0089_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold78 (.A(\gamepad.driver.shift_reg[0] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0087_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold80 (.A(\gamepad.driver.shift_reg[8] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0095_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold82 (.A(\gamepad.driver.shift_reg[1] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold83 (.A(\gamepad.driver.shift_reg[7] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0094_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold85 (.A(\gamepad.decoder.data_reg[6] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold86 (.A(\gamepad.decoder.data_reg[5] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold87 (.A(\pix_x[2] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0476_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0039_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold90 (.A(\gamepad.driver.shift_reg[4] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold91 (.A(\color_index[1] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0071_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pix_x[6] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0480_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold95 (.A(\palette_inst.rrggbb[3] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0018_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0692_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pix_x[1] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0475_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold100 (.A(\pix_x[9] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0804_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0005_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold103 (.A(\pix_x[3] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0477_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold105 (.A(\palette_inst.rrggbb[1] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold106 (.A(\pix_y[9] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold107 (.A(\pix_y[7] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0112_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold109 (.A(\pix_x[8] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0483_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold111 (.A(\pix_x[4] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold112 (.A(\pix_y[5] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold113 (.A(\pix_y[3] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0006_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold115 (.A(\pix_y[1] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0722_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold117 (.A(\pix_y[4] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold118 (.A(\logo_top[2] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold119 (.A(\pix_x[7] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold120 (.A(\pix_y[0] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0107_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold122 (.A(\pix_x[7] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold123 (.A(\logo_top[3] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold124 (.A(\logo_top[8] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold125 (.A(\pix_x[5] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0015_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold127 (.A(\logo_top[4] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0016_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold129 (.A(dir_y),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold130 (.A(\logo_top[1] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold131 (.A(\logo_top[6] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold132 (.A(\logo_left[8] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold133 (.A(\logo_top[9] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0008_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0051_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold136 (.A(\pix_y[6] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold137 (.A(\pix_y[8] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0741_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold139 (.A(\logo_left[9] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold140 (.A(\logo_left[5] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold141 (.A(\logo_top[7] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold142 (.A(\logo_left[6] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold143 (.A(\logo_left[2] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold144 (.A(dir_x),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold145 (.A(\logo_top[5] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold146 (.A(\logo_left[3] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold147 (.A(\logo_left[7] ),
    .X(net271));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_4 FILLER_0_49 ();
 sg13g2_decap_4 FILLER_0_77 ();
 sg13g2_fill_2 FILLER_0_90 ();
 sg13g2_fill_1 FILLER_0_92 ();
 sg13g2_fill_2 FILLER_0_107 ();
 sg13g2_fill_2 FILLER_0_114 ();
 sg13g2_fill_2 FILLER_0_127 ();
 sg13g2_fill_1 FILLER_0_129 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_4 FILLER_0_141 ();
 sg13g2_fill_2 FILLER_0_163 ();
 sg13g2_fill_1 FILLER_0_177 ();
 sg13g2_fill_1 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_4 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_214 ();
 sg13g2_fill_2 FILLER_0_219 ();
 sg13g2_fill_1 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_4 FILLER_0_237 ();
 sg13g2_fill_1 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_fill_1 FILLER_0_269 ();
 sg13g2_fill_2 FILLER_0_290 ();
 sg13g2_fill_1 FILLER_0_305 ();
 sg13g2_decap_4 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_fill_1 FILLER_1_42 ();
 sg13g2_decap_4 FILLER_1_47 ();
 sg13g2_fill_2 FILLER_1_59 ();
 sg13g2_fill_1 FILLER_1_61 ();
 sg13g2_fill_2 FILLER_1_74 ();
 sg13g2_fill_1 FILLER_1_76 ();
 sg13g2_fill_1 FILLER_1_132 ();
 sg13g2_decap_4 FILLER_1_148 ();
 sg13g2_fill_2 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_169 ();
 sg13g2_fill_2 FILLER_1_176 ();
 sg13g2_fill_1 FILLER_1_178 ();
 sg13g2_fill_1 FILLER_1_199 ();
 sg13g2_fill_2 FILLER_1_214 ();
 sg13g2_fill_2 FILLER_1_274 ();
 sg13g2_fill_2 FILLER_1_284 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_fill_2 FILLER_1_304 ();
 sg13g2_fill_1 FILLER_1_306 ();
 sg13g2_fill_1 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_21 ();
 sg13g2_decap_4 FILLER_2_31 ();
 sg13g2_fill_1 FILLER_2_40 ();
 sg13g2_fill_1 FILLER_2_61 ();
 sg13g2_fill_1 FILLER_2_72 ();
 sg13g2_fill_2 FILLER_2_79 ();
 sg13g2_fill_1 FILLER_2_132 ();
 sg13g2_fill_2 FILLER_2_158 ();
 sg13g2_fill_1 FILLER_2_160 ();
 sg13g2_fill_2 FILLER_2_166 ();
 sg13g2_fill_1 FILLER_2_201 ();
 sg13g2_fill_2 FILLER_2_216 ();
 sg13g2_fill_2 FILLER_2_240 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_fill_2 FILLER_2_289 ();
 sg13g2_fill_1 FILLER_2_291 ();
 sg13g2_fill_2 FILLER_2_319 ();
 sg13g2_decap_4 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_43 ();
 sg13g2_fill_2 FILLER_3_82 ();
 sg13g2_decap_4 FILLER_3_93 ();
 sg13g2_decap_4 FILLER_3_139 ();
 sg13g2_fill_2 FILLER_3_175 ();
 sg13g2_fill_2 FILLER_3_191 ();
 sg13g2_fill_2 FILLER_3_198 ();
 sg13g2_decap_4 FILLER_3_211 ();
 sg13g2_fill_1 FILLER_3_215 ();
 sg13g2_fill_2 FILLER_3_240 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_fill_2 FILLER_3_248 ();
 sg13g2_fill_2 FILLER_3_265 ();
 sg13g2_fill_1 FILLER_3_267 ();
 sg13g2_fill_2 FILLER_3_285 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_1 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_fill_1 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_5 ();
 sg13g2_decap_8 FILLER_4_10 ();
 sg13g2_decap_4 FILLER_4_26 ();
 sg13g2_fill_2 FILLER_4_38 ();
 sg13g2_fill_1 FILLER_4_40 ();
 sg13g2_fill_2 FILLER_4_54 ();
 sg13g2_fill_2 FILLER_4_65 ();
 sg13g2_fill_2 FILLER_4_73 ();
 sg13g2_fill_1 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_decap_4 FILLER_4_106 ();
 sg13g2_fill_2 FILLER_4_123 ();
 sg13g2_fill_1 FILLER_4_125 ();
 sg13g2_fill_2 FILLER_4_151 ();
 sg13g2_decap_4 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_176 ();
 sg13g2_fill_2 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_201 ();
 sg13g2_decap_4 FILLER_4_212 ();
 sg13g2_fill_1 FILLER_4_216 ();
 sg13g2_fill_2 FILLER_4_243 ();
 sg13g2_fill_1 FILLER_4_245 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_fill_2 FILLER_4_262 ();
 sg13g2_fill_2 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_decap_4 FILLER_5_23 ();
 sg13g2_fill_2 FILLER_5_57 ();
 sg13g2_fill_2 FILLER_5_65 ();
 sg13g2_fill_1 FILLER_5_94 ();
 sg13g2_fill_2 FILLER_5_111 ();
 sg13g2_fill_1 FILLER_5_118 ();
 sg13g2_fill_2 FILLER_5_124 ();
 sg13g2_decap_4 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_163 ();
 sg13g2_fill_2 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_2 FILLER_5_190 ();
 sg13g2_fill_1 FILLER_5_192 ();
 sg13g2_fill_1 FILLER_5_215 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_decap_4 FILLER_5_278 ();
 sg13g2_fill_2 FILLER_5_313 ();
 sg13g2_fill_2 FILLER_5_325 ();
 sg13g2_fill_1 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_40 ();
 sg13g2_decap_4 FILLER_6_76 ();
 sg13g2_fill_2 FILLER_6_86 ();
 sg13g2_fill_1 FILLER_6_88 ();
 sg13g2_fill_2 FILLER_6_115 ();
 sg13g2_decap_8 FILLER_6_125 ();
 sg13g2_fill_2 FILLER_6_132 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_fill_2 FILLER_6_177 ();
 sg13g2_fill_1 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_206 ();
 sg13g2_fill_2 FILLER_6_218 ();
 sg13g2_fill_1 FILLER_6_220 ();
 sg13g2_fill_2 FILLER_6_226 ();
 sg13g2_fill_1 FILLER_6_254 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_fill_1 FILLER_6_266 ();
 sg13g2_decap_4 FILLER_6_287 ();
 sg13g2_fill_1 FILLER_6_291 ();
 sg13g2_fill_2 FILLER_6_301 ();
 sg13g2_fill_1 FILLER_6_303 ();
 sg13g2_fill_1 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_16 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_fill_2 FILLER_7_75 ();
 sg13g2_fill_2 FILLER_7_97 ();
 sg13g2_fill_1 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_111 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_decap_4 FILLER_7_148 ();
 sg13g2_fill_1 FILLER_7_152 ();
 sg13g2_fill_2 FILLER_7_169 ();
 sg13g2_decap_4 FILLER_7_224 ();
 sg13g2_decap_4 FILLER_7_248 ();
 sg13g2_fill_1 FILLER_7_256 ();
 sg13g2_fill_2 FILLER_7_262 ();
 sg13g2_fill_1 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_decap_4 FILLER_7_297 ();
 sg13g2_fill_1 FILLER_7_301 ();
 sg13g2_fill_2 FILLER_7_321 ();
 sg13g2_decap_4 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_2 FILLER_8_29 ();
 sg13g2_fill_1 FILLER_8_31 ();
 sg13g2_fill_2 FILLER_8_48 ();
 sg13g2_fill_1 FILLER_8_50 ();
 sg13g2_fill_2 FILLER_8_73 ();
 sg13g2_fill_2 FILLER_8_97 ();
 sg13g2_fill_1 FILLER_8_99 ();
 sg13g2_fill_1 FILLER_8_106 ();
 sg13g2_fill_2 FILLER_8_134 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_189 ();
 sg13g2_fill_2 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_218 ();
 sg13g2_decap_4 FILLER_8_224 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_fill_2 FILLER_8_261 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_decap_4 FILLER_8_293 ();
 sg13g2_decap_4 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_4 FILLER_8_397 ();
 sg13g2_fill_2 FILLER_8_401 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_fill_2 FILLER_9_71 ();
 sg13g2_fill_1 FILLER_9_104 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_1 FILLER_9_132 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_149 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_168 ();
 sg13g2_fill_2 FILLER_9_177 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_2 FILLER_9_221 ();
 sg13g2_fill_2 FILLER_9_254 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_fill_2 FILLER_9_299 ();
 sg13g2_fill_1 FILLER_9_318 ();
 sg13g2_fill_2 FILLER_9_344 ();
 sg13g2_fill_1 FILLER_9_346 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_fill_2 FILLER_9_390 ();
 sg13g2_fill_1 FILLER_9_392 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_23 ();
 sg13g2_fill_2 FILLER_10_36 ();
 sg13g2_fill_2 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_57 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_fill_1 FILLER_10_78 ();
 sg13g2_fill_1 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_121 ();
 sg13g2_fill_1 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_129 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_166 ();
 sg13g2_decap_4 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_192 ();
 sg13g2_decap_4 FILLER_10_220 ();
 sg13g2_decap_4 FILLER_10_232 ();
 sg13g2_fill_2 FILLER_10_265 ();
 sg13g2_fill_1 FILLER_10_267 ();
 sg13g2_fill_2 FILLER_10_279 ();
 sg13g2_fill_1 FILLER_10_281 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_decap_4 FILLER_10_318 ();
 sg13g2_fill_2 FILLER_10_345 ();
 sg13g2_fill_2 FILLER_10_372 ();
 sg13g2_decap_4 FILLER_10_380 ();
 sg13g2_fill_1 FILLER_10_384 ();
 sg13g2_fill_1 FILLER_10_388 ();
 sg13g2_fill_2 FILLER_10_398 ();
 sg13g2_fill_1 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_56 ();
 sg13g2_fill_2 FILLER_11_134 ();
 sg13g2_fill_2 FILLER_11_150 ();
 sg13g2_fill_2 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_159 ();
 sg13g2_fill_2 FILLER_11_169 ();
 sg13g2_decap_4 FILLER_11_200 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_fill_2 FILLER_11_253 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_fill_1 FILLER_11_313 ();
 sg13g2_fill_2 FILLER_11_387 ();
 sg13g2_fill_1 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_12_51 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_113 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_154 ();
 sg13g2_decap_4 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_decap_4 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_249 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_decap_4 FILLER_12_292 ();
 sg13g2_fill_2 FILLER_12_296 ();
 sg13g2_decap_4 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_307 ();
 sg13g2_fill_2 FILLER_12_314 ();
 sg13g2_fill_2 FILLER_12_357 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_41 ();
 sg13g2_fill_2 FILLER_13_57 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_2 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_90 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_162 ();
 sg13g2_fill_2 FILLER_13_180 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_211 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_fill_1 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_272 ();
 sg13g2_fill_1 FILLER_13_274 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_fill_2 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_322 ();
 sg13g2_fill_2 FILLER_13_364 ();
 sg13g2_fill_1 FILLER_13_370 ();
 sg13g2_fill_1 FILLER_13_383 ();
 sg13g2_fill_2 FILLER_13_394 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_44 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_135 ();
 sg13g2_fill_1 FILLER_14_137 ();
 sg13g2_fill_2 FILLER_14_165 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_272 ();
 sg13g2_fill_2 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_389 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_31 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_fill_2 FILLER_15_87 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_143 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_1 FILLER_15_177 ();
 sg13g2_fill_2 FILLER_15_198 ();
 sg13g2_fill_1 FILLER_15_200 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_2 FILLER_15_246 ();
 sg13g2_fill_1 FILLER_15_272 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_fill_2 FILLER_15_354 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_fill_1 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_fill_2 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_248 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_373 ();
 sg13g2_fill_2 FILLER_17_50 ();
 sg13g2_fill_2 FILLER_17_57 ();
 sg13g2_fill_2 FILLER_17_67 ();
 sg13g2_fill_1 FILLER_17_69 ();
 sg13g2_fill_2 FILLER_17_74 ();
 sg13g2_fill_2 FILLER_17_89 ();
 sg13g2_fill_2 FILLER_17_102 ();
 sg13g2_fill_2 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_fill_2 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_194 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_fill_2 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_325 ();
 sg13g2_fill_1 FILLER_17_358 ();
 sg13g2_fill_1 FILLER_17_368 ();
 sg13g2_fill_2 FILLER_18_24 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_2 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_181 ();
 sg13g2_fill_1 FILLER_18_183 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_fill_2 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_73 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_103 ();
 sg13g2_fill_2 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_279 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_2 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_61 ();
 sg13g2_fill_1 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_81 ();
 sg13g2_fill_2 FILLER_21_109 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_fill_1 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_fill_2 FILLER_22_61 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_2 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_fill_2 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_290 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_385 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_22 ();
 sg13g2_fill_1 FILLER_23_66 ();
 sg13g2_fill_1 FILLER_23_76 ();
 sg13g2_fill_2 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_2 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_fill_2 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_395 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_2 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_fill_2 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_287 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_fill_2 FILLER_28_245 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_29_78 ();
 sg13g2_fill_1 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_197 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_30_13 ();
 sg13g2_fill_2 FILLER_30_24 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_239 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_333 ();
 sg13g2_fill_2 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_58 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_fill_1 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_fill_2 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_360 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_299 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_31 ();
 sg13g2_fill_2 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_362 ();
 sg13g2_fill_1 FILLER_38_372 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule
