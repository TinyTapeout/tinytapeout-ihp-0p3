module tt_um_calonso88_spi_test (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire \config_regs[0] ;
 wire \config_regs[10] ;
 wire \config_regs[11] ;
 wire \config_regs[12] ;
 wire \config_regs[13] ;
 wire \config_regs[14] ;
 wire \config_regs[15] ;
 wire \config_regs[16] ;
 wire \config_regs[17] ;
 wire \config_regs[18] ;
 wire \config_regs[19] ;
 wire \config_regs[1] ;
 wire \config_regs[20] ;
 wire \config_regs[21] ;
 wire \config_regs[22] ;
 wire \config_regs[23] ;
 wire \config_regs[24] ;
 wire \config_regs[25] ;
 wire \config_regs[26] ;
 wire \config_regs[27] ;
 wire \config_regs[28] ;
 wire \config_regs[29] ;
 wire \config_regs[2] ;
 wire \config_regs[30] ;
 wire \config_regs[31] ;
 wire \config_regs[32] ;
 wire \config_regs[33] ;
 wire \config_regs[34] ;
 wire \config_regs[35] ;
 wire \config_regs[36] ;
 wire \config_regs[37] ;
 wire \config_regs[38] ;
 wire \config_regs[39] ;
 wire \config_regs[3] ;
 wire \config_regs[40] ;
 wire \config_regs[41] ;
 wire \config_regs[42] ;
 wire \config_regs[43] ;
 wire \config_regs[44] ;
 wire \config_regs[45] ;
 wire \config_regs[46] ;
 wire \config_regs[47] ;
 wire \config_regs[48] ;
 wire \config_regs[49] ;
 wire \config_regs[4] ;
 wire \config_regs[50] ;
 wire \config_regs[51] ;
 wire \config_regs[52] ;
 wire \config_regs[53] ;
 wire \config_regs[54] ;
 wire \config_regs[55] ;
 wire \config_regs[56] ;
 wire \config_regs[57] ;
 wire \config_regs[58] ;
 wire \config_regs[59] ;
 wire \config_regs[5] ;
 wire \config_regs[60] ;
 wire \config_regs[61] ;
 wire \config_regs[62] ;
 wire \config_regs[63] ;
 wire \config_regs[6] ;
 wire \config_regs[7] ;
 wire \config_regs[8] ;
 wire \config_regs[9] ;
 wire cpha_sync;
 wire cpol_sync;
 wire spi_clk_sync;
 wire spi_cs_n_sync;
 wire spi_miso;
 wire spi_mosi_sync;
 wire \spi_wrapper_i.reg_addr[0] ;
 wire \spi_wrapper_i.reg_addr[1] ;
 wire \spi_wrapper_i.reg_addr[2] ;
 wire \spi_wrapper_i.reg_addr[3] ;
 wire \spi_wrapper_i.reg_data_o[0] ;
 wire \spi_wrapper_i.reg_data_o[1] ;
 wire \spi_wrapper_i.reg_data_o[2] ;
 wire \spi_wrapper_i.reg_data_o[3] ;
 wire \spi_wrapper_i.reg_data_o[4] ;
 wire \spi_wrapper_i.reg_data_o[5] ;
 wire \spi_wrapper_i.reg_data_o[6] ;
 wire \spi_wrapper_i.reg_data_o[7] ;
 wire \spi_wrapper_i.reg_data_o_vld ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[3] ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.reg_rw ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[7] ;
 wire \spi_wrapper_i.spi_reg_inst.state[0] ;
 wire \spi_wrapper_i.spi_reg_inst.state[1] ;
 wire \spi_wrapper_i.spi_reg_inst.state[2] ;
 wire \spi_wrapper_i.spi_reg_inst.state[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[6] ;
 wire \synchronizer_spi_clk_inst.data_sync[1] ;
 wire \synchronizer_spi_cs_n_inst.data_sync[1] ;
 wire \synchronizer_spi_mode_cpha.data_sync[1] ;
 wire \synchronizer_spi_mode_cpol.data_sync[1] ;
 wire \synchronizer_spi_mosi_inst.data_sync[1] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;

 sg13g2_inv_1 _383_ (.Y(_132_),
    .A(\spi_wrapper_i.reg_addr[2] ));
 sg13g2_inv_1 _384_ (.Y(_133_),
    .A(_004_));
 sg13g2_inv_1 _385_ (.Y(_134_),
    .A(net37));
 sg13g2_inv_1 _386_ (.Y(_135_),
    .A(net44));
 sg13g2_inv_1 _387_ (.Y(_136_),
    .A(net232));
 sg13g2_inv_1 _388_ (.Y(_137_),
    .A(net20));
 sg13g2_inv_1 _389_ (.Y(_138_),
    .A(net242));
 sg13g2_nor3_1 _390_ (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ),
    .B(\spi_wrapper_i.spi_reg_inst.buffer_counter[0] ),
    .C(\spi_wrapper_i.spi_reg_inst.buffer_counter[2] ),
    .Y(_139_));
 sg13g2_nor2b_2 _391_ (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ),
    .B_N(_139_),
    .Y(_140_));
 sg13g2_nand2b_1 _392_ (.Y(_141_),
    .B(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .A_N(_140_));
 sg13g2_nand2_1 _393_ (.Y(_142_),
    .A(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ),
    .B(_139_));
 sg13g2_o21ai_1 _394_ (.B1(_142_),
    .Y(_143_),
    .A1(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .A2(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_and3_2 _395_ (.X(_144_),
    .A(net164),
    .B(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ),
    .C(_139_));
 sg13g2_nand2_1 _396_ (.Y(_145_),
    .A(net165),
    .B(net206));
 sg13g2_nor2_1 _397_ (.A(net232),
    .B(_145_),
    .Y(_146_));
 sg13g2_nor2_2 _398_ (.A(_144_),
    .B(_146_),
    .Y(_147_));
 sg13g2_a21oi_1 _399_ (.A1(_141_),
    .A2(_143_),
    .Y(_148_),
    .B1(_147_));
 sg13g2_nand2_1 _400_ (.Y(_149_),
    .A(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .B(_144_));
 sg13g2_nand2b_1 _401_ (.Y(_150_),
    .B(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .A_N(spi_cs_n_sync));
 sg13g2_nand3b_1 _402_ (.B(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .C(net165),
    .Y(_151_),
    .A_N(spi_cs_n_sync));
 sg13g2_a221oi_1 _403_ (.B2(net20),
    .C1(_148_),
    .B1(_151_),
    .A1(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .Y(_021_),
    .A2(_144_));
 sg13g2_nand2_1 _404_ (.Y(_152_),
    .A(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_140_));
 sg13g2_nand2_1 _405_ (.Y(_153_),
    .A(net164),
    .B(net44));
 sg13g2_o21ai_1 _406_ (.B1(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .Y(_154_),
    .A1(_140_),
    .A2(_147_));
 sg13g2_o21ai_1 _407_ (.B1(_154_),
    .Y(_000_),
    .A1(net37),
    .A2(_153_));
 sg13g2_nand2_1 _408_ (.Y(_155_),
    .A(net30),
    .B(_144_));
 sg13g2_o21ai_1 _409_ (.B1(net125),
    .Y(_001_),
    .A1(net164),
    .A2(_135_));
 sg13g2_nand2_1 _410_ (.Y(_156_),
    .A(net30),
    .B(_147_));
 sg13g2_o21ai_1 _411_ (.B1(net31),
    .Y(_002_),
    .A1(_137_),
    .A2(_151_));
 sg13g2_nand2_1 _412_ (.Y(_157_),
    .A(net233),
    .B(_147_));
 sg13g2_o21ai_1 _413_ (.B1(_157_),
    .Y(_003_),
    .A1(_134_),
    .A2(_153_));
 sg13g2_xor2_1 _414_ (.B(cpol_sync),
    .A(cpha_sync),
    .X(_158_));
 sg13g2_nand3b_1 _415_ (.B(uio_oe[3]),
    .C(spi_clk_sync),
    .Y(_159_),
    .A_N(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_nand2b_1 _416_ (.Y(_160_),
    .B(_159_),
    .A_N(_158_));
 sg13g2_nand3b_1 _417_ (.B(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .C(uio_oe[3]),
    .Y(_161_),
    .A_N(spi_clk_sync));
 sg13g2_nand2_1 _418_ (.Y(_162_),
    .A(_158_),
    .B(_161_));
 sg13g2_and3_2 _419_ (.X(_163_),
    .A(net164),
    .B(_160_),
    .C(_162_));
 sg13g2_nand3_1 _420_ (.B(_160_),
    .C(_162_),
    .A(net164),
    .Y(_164_));
 sg13g2_nand2_1 _421_ (.Y(_165_),
    .A(_142_),
    .B(_163_));
 sg13g2_a21oi_1 _422_ (.A1(_142_),
    .A2(_163_),
    .Y(_166_),
    .B1(net240));
 sg13g2_a21oi_1 _423_ (.A1(net240),
    .A2(_163_),
    .Y(_022_),
    .B1(net241));
 sg13g2_nand3_1 _424_ (.B(net240),
    .C(_163_),
    .A(net246),
    .Y(_167_));
 sg13g2_a21o_1 _425_ (.A2(_163_),
    .A1(net240),
    .B1(net246),
    .X(_168_));
 sg13g2_and2_1 _426_ (.A(_167_),
    .B(_168_),
    .X(_023_));
 sg13g2_nand3_1 _427_ (.B(net240),
    .C(net181),
    .A(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ),
    .Y(_169_));
 sg13g2_xnor2_1 _428_ (.Y(_024_),
    .A(net181),
    .B(_167_));
 sg13g2_nand3b_1 _429_ (.B(_164_),
    .C(net244),
    .Y(_170_),
    .A_N(_144_));
 sg13g2_xor2_1 _430_ (.B(_169_),
    .A(net244),
    .X(_171_));
 sg13g2_o21ai_1 _431_ (.B1(_170_),
    .Y(_025_),
    .A1(_165_),
    .A2(_171_));
 sg13g2_nor2_1 _432_ (.A(net43),
    .B(net125),
    .Y(_172_));
 sg13g2_a21oi_1 _433_ (.A1(_134_),
    .A2(net125),
    .Y(_026_),
    .B1(_172_));
 sg13g2_mux2_1 _434_ (.A0(net185),
    .A1(net222),
    .S(net125),
    .X(_027_));
 sg13g2_mux2_1 _435_ (.A0(net210),
    .A1(net226),
    .S(_155_),
    .X(_028_));
 sg13g2_nor2_1 _436_ (.A(net209),
    .B(net125),
    .Y(_173_));
 sg13g2_a21oi_1 _437_ (.A1(_132_),
    .A2(net125),
    .Y(_029_),
    .B1(_173_));
 sg13g2_nor2_1 _438_ (.A(net215),
    .B(net125),
    .Y(_174_));
 sg13g2_a21oi_1 _439_ (.A1(_138_),
    .A2(net125),
    .Y(_030_),
    .B1(_174_));
 sg13g2_nand2b_1 _440_ (.Y(_175_),
    .B(net234),
    .A_N(net164));
 sg13g2_o21ai_1 _441_ (.B1(_175_),
    .Y(_031_),
    .A1(_134_),
    .A2(net129));
 sg13g2_mux2_1 _442_ (.A0(net185),
    .A1(net141),
    .S(net129),
    .X(_032_));
 sg13g2_mux2_1 _443_ (.A0(net210),
    .A1(net140),
    .S(net129),
    .X(_033_));
 sg13g2_mux2_1 _444_ (.A0(net209),
    .A1(net139),
    .S(net129),
    .X(_034_));
 sg13g2_mux2_1 _445_ (.A0(net215),
    .A1(net138),
    .S(net129),
    .X(_035_));
 sg13g2_mux2_1 _446_ (.A0(net121),
    .A1(net137),
    .S(net129),
    .X(_036_));
 sg13g2_mux2_1 _447_ (.A0(net199),
    .A1(net136),
    .S(net129),
    .X(_037_));
 sg13g2_mux2_1 _448_ (.A0(net224),
    .A1(net135),
    .S(net129),
    .X(_038_));
 sg13g2_mux2_1 _449_ (.A0(net43),
    .A1(net134),
    .S(_149_),
    .X(_039_));
 sg13g2_mux2_1 _450_ (.A0(_161_),
    .A1(_159_),
    .S(_158_),
    .X(_176_));
 sg13g2_nand3_1 _451_ (.B(net128),
    .C(_176_),
    .A(_150_),
    .Y(_177_));
 sg13g2_nand2_2 _452_ (.Y(_178_),
    .A(net166),
    .B(_177_));
 sg13g2_nand2_1 _453_ (.Y(_179_),
    .A(net35),
    .B(_178_));
 sg13g2_or2_1 _454_ (.X(_180_),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .A(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_a21oi_2 _455_ (.B1(_133_),
    .Y(_181_),
    .A2(_180_),
    .A1(_132_));
 sg13g2_a21o_1 _456_ (.A2(_180_),
    .A1(_132_),
    .B1(_133_),
    .X(_182_));
 sg13g2_nand2_1 _457_ (.Y(_183_),
    .A(_005_),
    .B(_181_));
 sg13g2_nand2b_2 _458_ (.Y(_184_),
    .B(\spi_wrapper_i.reg_addr[1] ),
    .A_N(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_nor2_2 _459_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_184_),
    .Y(_185_));
 sg13g2_nand2_1 _460_ (.Y(_186_),
    .A(\config_regs[16] ),
    .B(net132));
 sg13g2_nand2_2 _461_ (.Y(_187_),
    .A(\spi_wrapper_i.reg_addr[1] ),
    .B(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_nor2_2 _462_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_187_),
    .Y(_188_));
 sg13g2_nand2b_2 _463_ (.Y(_189_),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .A_N(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_nor2_2 _464_ (.A(net142),
    .B(_189_),
    .Y(_190_));
 sg13g2_a22oi_1 _465_ (.Y(_191_),
    .B1(_190_),
    .B2(\config_regs[40] ),
    .A2(net131),
    .A1(\config_regs[24] ));
 sg13g2_nor2_2 _466_ (.A(net142),
    .B(_187_),
    .Y(_192_));
 sg13g2_nor2_1 _467_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_189_),
    .Y(_193_));
 sg13g2_a22oi_1 _468_ (.Y(_194_),
    .B1(_193_),
    .B2(\config_regs[8] ),
    .A2(_192_),
    .A1(\config_regs[56] ));
 sg13g2_nor2_2 _469_ (.A(net142),
    .B(_184_),
    .Y(_195_));
 sg13g2_a21oi_1 _470_ (.A1(\config_regs[48] ),
    .A2(_195_),
    .Y(_196_),
    .B1(_181_));
 sg13g2_nand4_1 _471_ (.B(_191_),
    .C(_194_),
    .A(_186_),
    .Y(_197_),
    .D(_196_));
 sg13g2_nor3_2 _472_ (.A(\spi_wrapper_i.reg_addr[1] ),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .C(net142),
    .Y(_198_));
 sg13g2_a221oi_1 _473_ (.B2(\config_regs[32] ),
    .C1(\spi_wrapper_i.reg_addr[3] ),
    .B1(net133),
    .A1(_183_),
    .Y(_199_),
    .A2(_197_));
 sg13g2_o21ai_1 _474_ (.B1(\spi_wrapper_i.reg_addr[3] ),
    .Y(_200_),
    .A1(\spi_wrapper_i.reg_addr[0] ),
    .A2(_004_));
 sg13g2_nor2_1 _475_ (.A(net131),
    .B(_200_),
    .Y(_201_));
 sg13g2_nand4_1 _476_ (.B(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .C(_140_),
    .A(net166),
    .Y(_202_),
    .D(_150_));
 sg13g2_or2_1 _477_ (.X(_203_),
    .B(_202_),
    .A(_201_));
 sg13g2_o21ai_1 _478_ (.B1(_179_),
    .Y(_040_),
    .A1(_199_),
    .A2(_203_));
 sg13g2_nand2_1 _479_ (.Y(_204_),
    .A(net28),
    .B(_178_));
 sg13g2_and2_1 _480_ (.A(\config_regs[33] ),
    .B(net133),
    .X(_205_));
 sg13g2_a22oi_1 _481_ (.Y(_206_),
    .B1(net130),
    .B2(\config_regs[9] ),
    .A2(net131),
    .A1(\config_regs[25] ));
 sg13g2_nor2_2 _482_ (.A(\spi_wrapper_i.reg_addr[3] ),
    .B(_181_),
    .Y(_207_));
 sg13g2_a221oi_1 _483_ (.B2(\config_regs[41] ),
    .C1(_205_),
    .B1(_190_),
    .A1(\config_regs[17] ),
    .Y(_208_),
    .A2(net132));
 sg13g2_a22oi_1 _484_ (.Y(_209_),
    .B1(_195_),
    .B2(\config_regs[49] ),
    .A2(_192_),
    .A1(\config_regs[57] ));
 sg13g2_nand4_1 _485_ (.B(_207_),
    .C(_208_),
    .A(_206_),
    .Y(_210_),
    .D(_209_));
 sg13g2_xor2_1 _486_ (.B(\spi_wrapper_i.reg_addr[0] ),
    .A(\spi_wrapper_i.reg_addr[1] ),
    .X(_211_));
 sg13g2_nor2_1 _487_ (.A(net142),
    .B(_211_),
    .Y(_212_));
 sg13g2_nor4_1 _488_ (.A(_138_),
    .B(_181_),
    .C(net132),
    .D(_212_),
    .Y(_213_));
 sg13g2_nor2_2 _489_ (.A(\spi_wrapper_i.reg_addr[3] ),
    .B(_182_),
    .Y(_214_));
 sg13g2_a21oi_1 _490_ (.A1(_007_),
    .A2(_214_),
    .Y(_215_),
    .B1(_213_));
 sg13g2_a21oi_1 _491_ (.A1(_210_),
    .A2(_215_),
    .Y(_216_),
    .B1(net127));
 sg13g2_nand3_1 _492_ (.B(_150_),
    .C(_177_),
    .A(net166),
    .Y(_217_));
 sg13g2_a21o_1 _493_ (.A2(net127),
    .A1(_006_),
    .B1(_216_),
    .X(_218_));
 sg13g2_o21ai_1 _494_ (.B1(_204_),
    .Y(_041_),
    .A1(_217_),
    .A2(_218_));
 sg13g2_and2_1 _495_ (.A(\config_regs[34] ),
    .B(net133),
    .X(_219_));
 sg13g2_a22oi_1 _496_ (.Y(_220_),
    .B1(_188_),
    .B2(\config_regs[26] ),
    .A2(_185_),
    .A1(\config_regs[18] ));
 sg13g2_a221oi_1 _497_ (.B2(\config_regs[10] ),
    .C1(_219_),
    .B1(net130),
    .A1(\config_regs[42] ),
    .Y(_221_),
    .A2(_190_));
 sg13g2_a22oi_1 _498_ (.Y(_222_),
    .B1(_195_),
    .B2(\config_regs[50] ),
    .A2(_192_),
    .A1(\config_regs[58] ));
 sg13g2_nand4_1 _499_ (.B(_220_),
    .C(_221_),
    .A(_207_),
    .Y(_223_),
    .D(_222_));
 sg13g2_a21oi_1 _500_ (.A1(_009_),
    .A2(_214_),
    .Y(_224_),
    .B1(_201_));
 sg13g2_a21oi_1 _501_ (.A1(_223_),
    .A2(_224_),
    .Y(_225_),
    .B1(net127));
 sg13g2_a21o_1 _502_ (.A2(net127),
    .A1(_008_),
    .B1(_225_),
    .X(_226_));
 sg13g2_nand2_1 _503_ (.Y(_227_),
    .A(net24),
    .B(_178_));
 sg13g2_o21ai_1 _504_ (.B1(_227_),
    .Y(_042_),
    .A1(_217_),
    .A2(_226_));
 sg13g2_nand2_1 _505_ (.Y(_228_),
    .A(\config_regs[11] ),
    .B(net130));
 sg13g2_a22oi_1 _506_ (.Y(_229_),
    .B1(_195_),
    .B2(\config_regs[51] ),
    .A2(_192_),
    .A1(\config_regs[59] ));
 sg13g2_a22oi_1 _507_ (.Y(_230_),
    .B1(_198_),
    .B2(\config_regs[35] ),
    .A2(_185_),
    .A1(\config_regs[19] ));
 sg13g2_a22oi_1 _508_ (.Y(_231_),
    .B1(_190_),
    .B2(\config_regs[43] ),
    .A2(_188_),
    .A1(\config_regs[27] ));
 sg13g2_and4_1 _509_ (.A(_228_),
    .B(_229_),
    .C(_230_),
    .D(_231_),
    .X(_232_));
 sg13g2_a221oi_1 _510_ (.B2(_207_),
    .C1(_213_),
    .B1(_232_),
    .A1(_011_),
    .Y(_233_),
    .A2(_214_));
 sg13g2_nand2_1 _511_ (.Y(_234_),
    .A(_010_),
    .B(net126));
 sg13g2_o21ai_1 _512_ (.B1(_234_),
    .Y(_235_),
    .A1(net126),
    .A2(_233_));
 sg13g2_nand2_1 _513_ (.Y(_236_),
    .A(net33),
    .B(_178_));
 sg13g2_o21ai_1 _514_ (.B1(_236_),
    .Y(_043_),
    .A1(_217_),
    .A2(_235_));
 sg13g2_nand2_1 _515_ (.Y(_237_),
    .A(net26),
    .B(_178_));
 sg13g2_and2_1 _516_ (.A(\config_regs[60] ),
    .B(_192_),
    .X(_238_));
 sg13g2_a221oi_1 _517_ (.B2(\config_regs[12] ),
    .C1(_238_),
    .B1(net130),
    .A1(\config_regs[20] ),
    .Y(_239_),
    .A2(net132));
 sg13g2_a22oi_1 _518_ (.Y(_240_),
    .B1(_195_),
    .B2(\config_regs[52] ),
    .A2(net131),
    .A1(\config_regs[28] ));
 sg13g2_a22oi_1 _519_ (.Y(_241_),
    .B1(net133),
    .B2(\config_regs[36] ),
    .A2(_190_),
    .A1(\config_regs[44] ));
 sg13g2_nand4_1 _520_ (.B(_239_),
    .C(_240_),
    .A(_207_),
    .Y(_242_),
    .D(_241_));
 sg13g2_nor4_1 _521_ (.A(_138_),
    .B(net131),
    .C(net130),
    .D(_212_),
    .Y(_243_));
 sg13g2_a21oi_1 _522_ (.A1(_013_),
    .A2(_214_),
    .Y(_244_),
    .B1(_243_));
 sg13g2_a21oi_1 _523_ (.A1(_242_),
    .A2(_244_),
    .Y(_245_),
    .B1(net126));
 sg13g2_a21o_1 _524_ (.A2(net126),
    .A1(_012_),
    .B1(_217_),
    .X(_246_));
 sg13g2_o21ai_1 _525_ (.B1(_237_),
    .Y(_044_),
    .A1(_245_),
    .A2(_246_));
 sg13g2_nand2_1 _526_ (.Y(_247_),
    .A(\config_regs[61] ),
    .B(_192_));
 sg13g2_a22oi_1 _527_ (.Y(_248_),
    .B1(_195_),
    .B2(\config_regs[53] ),
    .A2(net131),
    .A1(\config_regs[29] ));
 sg13g2_a22oi_1 _528_ (.Y(_249_),
    .B1(_190_),
    .B2(\config_regs[45] ),
    .A2(net132),
    .A1(\config_regs[21] ));
 sg13g2_a22oi_1 _529_ (.Y(_250_),
    .B1(net133),
    .B2(\config_regs[37] ),
    .A2(net130),
    .A1(\config_regs[13] ));
 sg13g2_and4_1 _530_ (.A(_247_),
    .B(_248_),
    .C(_249_),
    .D(_250_),
    .X(_251_));
 sg13g2_nor2_1 _531_ (.A(net132),
    .B(_200_),
    .Y(_252_));
 sg13g2_a221oi_1 _532_ (.B2(_207_),
    .C1(_252_),
    .B1(_251_),
    .A1(_015_),
    .Y(_253_),
    .A2(_214_));
 sg13g2_nand2_1 _533_ (.Y(_254_),
    .A(_014_),
    .B(net126));
 sg13g2_o21ai_1 _534_ (.B1(_254_),
    .Y(_255_),
    .A1(net126),
    .A2(_253_));
 sg13g2_nand2_1 _535_ (.Y(_256_),
    .A(net22),
    .B(_178_));
 sg13g2_o21ai_1 _536_ (.B1(_256_),
    .Y(_045_),
    .A1(_217_),
    .A2(_255_));
 sg13g2_and2_1 _537_ (.A(\config_regs[38] ),
    .B(net133),
    .X(_257_));
 sg13g2_a22oi_1 _538_ (.Y(_258_),
    .B1(net130),
    .B2(\config_regs[14] ),
    .A2(_190_),
    .A1(\config_regs[46] ));
 sg13g2_a22oi_1 _539_ (.Y(_259_),
    .B1(_195_),
    .B2(\config_regs[54] ),
    .A2(net131),
    .A1(\config_regs[30] ));
 sg13g2_a221oi_1 _540_ (.B2(\config_regs[62] ),
    .C1(_257_),
    .B1(_192_),
    .A1(\config_regs[22] ),
    .Y(_260_),
    .A2(net132));
 sg13g2_nand3_1 _541_ (.B(_259_),
    .C(_260_),
    .A(_258_),
    .Y(_261_));
 sg13g2_nand2_1 _542_ (.Y(_262_),
    .A(_207_),
    .B(_261_));
 sg13g2_nor3_1 _543_ (.A(\spi_wrapper_i.reg_addr[3] ),
    .B(_017_),
    .C(_182_),
    .Y(_263_));
 sg13g2_nor2_1 _544_ (.A(_138_),
    .B(_211_),
    .Y(_264_));
 sg13g2_nor3_1 _545_ (.A(net128),
    .B(_263_),
    .C(_264_),
    .Y(_265_));
 sg13g2_a221oi_1 _546_ (.B2(_265_),
    .C1(_217_),
    .B1(_262_),
    .A1(_016_),
    .Y(_266_),
    .A2(net126));
 sg13g2_a21o_1 _547_ (.A2(_178_),
    .A1(net41),
    .B1(_266_),
    .X(_046_));
 sg13g2_a22oi_1 _548_ (.Y(_267_),
    .B1(_192_),
    .B2(\config_regs[63] ),
    .A2(net132),
    .A1(\config_regs[23] ));
 sg13g2_a22oi_1 _549_ (.Y(_268_),
    .B1(_195_),
    .B2(\config_regs[55] ),
    .A2(net130),
    .A1(\config_regs[15] ));
 sg13g2_a22oi_1 _550_ (.Y(_269_),
    .B1(_190_),
    .B2(\config_regs[47] ),
    .A2(net131),
    .A1(\config_regs[31] ));
 sg13g2_a21oi_1 _551_ (.A1(\config_regs[39] ),
    .A2(net133),
    .Y(_270_),
    .B1(\spi_wrapper_i.reg_addr[3] ));
 sg13g2_and4_1 _552_ (.A(_267_),
    .B(_268_),
    .C(_269_),
    .D(_270_),
    .X(_271_));
 sg13g2_o21ai_1 _553_ (.B1(_182_),
    .Y(_272_),
    .A1(_252_),
    .A2(_271_));
 sg13g2_nand2_1 _554_ (.Y(_273_),
    .A(_019_),
    .B(_214_));
 sg13g2_a21oi_1 _555_ (.A1(_272_),
    .A2(_273_),
    .Y(_274_),
    .B1(net128));
 sg13g2_a21o_1 _556_ (.A2(net126),
    .A1(_018_),
    .B1(_217_),
    .X(_275_));
 sg13g2_nand2_1 _557_ (.Y(_276_),
    .A(net39),
    .B(_178_));
 sg13g2_o21ai_1 _558_ (.B1(_276_),
    .Y(_047_),
    .A1(_274_),
    .A2(_275_));
 sg13g2_nand2_2 _559_ (.Y(_277_),
    .A(\spi_wrapper_i.reg_data_o_vld ),
    .B(net166));
 sg13g2_nor3_2 _560_ (.A(net142),
    .B(_187_),
    .C(_277_),
    .Y(_278_));
 sg13g2_mux2_1 _561_ (.A0(net100),
    .A1(\spi_wrapper_i.reg_data_o[0] ),
    .S(_278_),
    .X(_048_));
 sg13g2_mux2_1 _562_ (.A0(net102),
    .A1(\spi_wrapper_i.reg_data_o[1] ),
    .S(_278_),
    .X(_049_));
 sg13g2_mux2_1 _563_ (.A0(net51),
    .A1(\spi_wrapper_i.reg_data_o[2] ),
    .S(_278_),
    .X(_050_));
 sg13g2_mux2_1 _564_ (.A0(net45),
    .A1(\spi_wrapper_i.reg_data_o[3] ),
    .S(_278_),
    .X(_051_));
 sg13g2_mux2_1 _565_ (.A0(net106),
    .A1(net137),
    .S(_278_),
    .X(_052_));
 sg13g2_mux2_1 _566_ (.A0(net191),
    .A1(net136),
    .S(_278_),
    .X(_053_));
 sg13g2_mux2_1 _567_ (.A0(net96),
    .A1(\spi_wrapper_i.reg_data_o[6] ),
    .S(_278_),
    .X(_054_));
 sg13g2_mux2_1 _568_ (.A0(net172),
    .A1(\spi_wrapper_i.reg_data_o[7] ),
    .S(_278_),
    .X(_055_));
 sg13g2_mux2_1 _569_ (.A0(net203),
    .A1(net196),
    .S(net165),
    .X(_056_));
 sg13g2_mux2_1 _570_ (.A0(net185),
    .A1(net203),
    .S(_163_),
    .X(_057_));
 sg13g2_mux2_1 _571_ (.A0(net185),
    .A1(net210),
    .S(_164_),
    .X(_058_));
 sg13g2_mux2_1 _572_ (.A0(net210),
    .A1(net209),
    .S(_164_),
    .X(_059_));
 sg13g2_mux2_1 _573_ (.A0(net209),
    .A1(net215),
    .S(_164_),
    .X(_060_));
 sg13g2_mux2_1 _574_ (.A0(net215),
    .A1(net121),
    .S(_164_),
    .X(_061_));
 sg13g2_mux2_1 _575_ (.A0(net121),
    .A1(net199),
    .S(_164_),
    .X(_062_));
 sg13g2_mux2_1 _576_ (.A0(net199),
    .A1(net224),
    .S(_164_),
    .X(_063_));
 sg13g2_mux2_1 _577_ (.A0(net43),
    .A1(net224),
    .S(_163_),
    .X(_064_));
 sg13g2_o21ai_1 _578_ (.B1(_145_),
    .Y(_065_),
    .A1(net165),
    .A2(_136_));
 sg13g2_nand3_1 _579_ (.B(net166),
    .C(net133),
    .A(\spi_wrapper_i.reg_data_o_vld ),
    .Y(_279_));
 sg13g2_mux2_1 _580_ (.A0(net141),
    .A1(net228),
    .S(_279_),
    .X(_066_));
 sg13g2_mux2_1 _581_ (.A0(net140),
    .A1(net237),
    .S(_279_),
    .X(_067_));
 sg13g2_mux2_1 _582_ (.A0(net139),
    .A1(net220),
    .S(_279_),
    .X(_068_));
 sg13g2_mux2_1 _583_ (.A0(net138),
    .A1(net230),
    .S(_279_),
    .X(_069_));
 sg13g2_mux2_1 _584_ (.A0(net65),
    .A1(\config_regs[36] ),
    .S(_279_),
    .X(_070_));
 sg13g2_mux2_1 _585_ (.A0(net136),
    .A1(net235),
    .S(_279_),
    .X(_071_));
 sg13g2_mux2_1 _586_ (.A0(net135),
    .A1(net218),
    .S(_279_),
    .X(_072_));
 sg13g2_mux2_1 _587_ (.A0(net134),
    .A1(net225),
    .S(_279_),
    .X(_073_));
 sg13g2_nor3_2 _588_ (.A(net142),
    .B(_189_),
    .C(_277_),
    .Y(_280_));
 sg13g2_mux2_1 _589_ (.A0(net216),
    .A1(net141),
    .S(_280_),
    .X(_074_));
 sg13g2_mux2_1 _590_ (.A0(net81),
    .A1(net140),
    .S(_280_),
    .X(_075_));
 sg13g2_mux2_1 _591_ (.A0(net197),
    .A1(net139),
    .S(_280_),
    .X(_076_));
 sg13g2_mux2_1 _592_ (.A0(net187),
    .A1(net138),
    .S(_280_),
    .X(_077_));
 sg13g2_mux2_1 _593_ (.A0(net70),
    .A1(net137),
    .S(_280_),
    .X(_078_));
 sg13g2_mux2_1 _594_ (.A0(net75),
    .A1(net136),
    .S(_280_),
    .X(_079_));
 sg13g2_mux2_1 _595_ (.A0(net49),
    .A1(net135),
    .S(_280_),
    .X(_080_));
 sg13g2_mux2_1 _596_ (.A0(net86),
    .A1(net134),
    .S(_280_),
    .X(_081_));
 sg13g2_nor3_2 _597_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_187_),
    .C(_277_),
    .Y(_281_));
 sg13g2_mux2_1 _598_ (.A0(net47),
    .A1(net141),
    .S(_281_),
    .X(_082_));
 sg13g2_mux2_1 _599_ (.A0(net53),
    .A1(net140),
    .S(_281_),
    .X(_083_));
 sg13g2_mux2_1 _600_ (.A0(net174),
    .A1(net139),
    .S(_281_),
    .X(_084_));
 sg13g2_mux2_1 _601_ (.A0(net90),
    .A1(net138),
    .S(_281_),
    .X(_085_));
 sg13g2_mux2_1 _602_ (.A0(net69),
    .A1(net137),
    .S(_281_),
    .X(_086_));
 sg13g2_mux2_1 _603_ (.A0(net59),
    .A1(net136),
    .S(_281_),
    .X(_087_));
 sg13g2_mux2_1 _604_ (.A0(net55),
    .A1(net135),
    .S(_281_),
    .X(_088_));
 sg13g2_mux2_1 _605_ (.A0(net94),
    .A1(net134),
    .S(_281_),
    .X(_089_));
 sg13g2_nor3_2 _606_ (.A(net142),
    .B(_184_),
    .C(_277_),
    .Y(_282_));
 sg13g2_mux2_1 _607_ (.A0(net104),
    .A1(net141),
    .S(_282_),
    .X(_090_));
 sg13g2_mux2_1 _608_ (.A0(net122),
    .A1(net140),
    .S(_282_),
    .X(_091_));
 sg13g2_mux2_1 _609_ (.A0(net189),
    .A1(net139),
    .S(_282_),
    .X(_092_));
 sg13g2_mux2_1 _610_ (.A0(net111),
    .A1(net138),
    .S(_282_),
    .X(_093_));
 sg13g2_mux2_1 _611_ (.A0(net114),
    .A1(net137),
    .S(_282_),
    .X(_094_));
 sg13g2_mux2_1 _612_ (.A0(net194),
    .A1(net136),
    .S(_282_),
    .X(_095_));
 sg13g2_mux2_1 _613_ (.A0(net98),
    .A1(net135),
    .S(_282_),
    .X(_096_));
 sg13g2_mux2_1 _614_ (.A0(net183),
    .A1(net134),
    .S(_282_),
    .X(_097_));
 sg13g2_nor3_2 _615_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_184_),
    .C(_277_),
    .Y(_283_));
 sg13g2_mux2_1 _616_ (.A0(net88),
    .A1(net141),
    .S(_283_),
    .X(_098_));
 sg13g2_mux2_1 _617_ (.A0(net170),
    .A1(net140),
    .S(_283_),
    .X(_099_));
 sg13g2_mux2_1 _618_ (.A0(net61),
    .A1(net139),
    .S(_283_),
    .X(_100_));
 sg13g2_mux2_1 _619_ (.A0(net71),
    .A1(net138),
    .S(_283_),
    .X(_101_));
 sg13g2_mux2_1 _620_ (.A0(net124),
    .A1(net137),
    .S(_283_),
    .X(_102_));
 sg13g2_mux2_1 _621_ (.A0(net109),
    .A1(net136),
    .S(_283_),
    .X(_103_));
 sg13g2_mux2_1 _622_ (.A0(net176),
    .A1(net135),
    .S(_283_),
    .X(_104_));
 sg13g2_mux2_1 _623_ (.A0(net73),
    .A1(net134),
    .S(_283_),
    .X(_105_));
 sg13g2_nor3_2 _624_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_189_),
    .C(_277_),
    .Y(_284_));
 sg13g2_mux2_1 _625_ (.A0(net115),
    .A1(net141),
    .S(_284_),
    .X(_106_));
 sg13g2_mux2_1 _626_ (.A0(net92),
    .A1(net140),
    .S(_284_),
    .X(_107_));
 sg13g2_mux2_1 _627_ (.A0(net178),
    .A1(net139),
    .S(_284_),
    .X(_108_));
 sg13g2_mux2_1 _628_ (.A0(net201),
    .A1(net138),
    .S(_284_),
    .X(_109_));
 sg13g2_mux2_1 _629_ (.A0(net83),
    .A1(net137),
    .S(_284_),
    .X(_110_));
 sg13g2_mux2_1 _630_ (.A0(net213),
    .A1(net136),
    .S(_284_),
    .X(_111_));
 sg13g2_mux2_1 _631_ (.A0(net207),
    .A1(net135),
    .S(_284_),
    .X(_112_));
 sg13g2_mux2_1 _632_ (.A0(net79),
    .A1(net134),
    .S(_284_),
    .X(_113_));
 sg13g2_nor3_2 _633_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(_180_),
    .C(_277_),
    .Y(_285_));
 sg13g2_mux2_1 _634_ (.A0(net84),
    .A1(net141),
    .S(_285_),
    .X(_114_));
 sg13g2_mux2_1 _635_ (.A0(net119),
    .A1(net140),
    .S(_285_),
    .X(_115_));
 sg13g2_mux2_1 _636_ (.A0(net67),
    .A1(net139),
    .S(_285_),
    .X(_116_));
 sg13g2_mux2_1 _637_ (.A0(net107),
    .A1(net138),
    .S(_285_),
    .X(_117_));
 sg13g2_mux2_1 _638_ (.A0(net180),
    .A1(net137),
    .S(_285_),
    .X(_118_));
 sg13g2_mux2_1 _639_ (.A0(net57),
    .A1(\spi_wrapper_i.reg_data_o[5] ),
    .S(_285_),
    .X(_119_));
 sg13g2_mux2_1 _640_ (.A0(net77),
    .A1(net135),
    .S(_285_),
    .X(_120_));
 sg13g2_mux2_1 _641_ (.A0(net63),
    .A1(net134),
    .S(_285_),
    .X(_121_));
 sg13g2_mux2_1 _642_ (.A0(net117),
    .A1(net1),
    .S(net167),
    .X(_122_));
 sg13g2_mux2_1 _643_ (.A0(net223),
    .A1(net113),
    .S(net167),
    .X(_123_));
 sg13g2_mux2_1 _644_ (.A0(net113),
    .A1(net2),
    .S(net167),
    .X(_124_));
 sg13g2_mux2_1 _645_ (.A0(net206),
    .A1(net193),
    .S(net164),
    .X(_125_));
 sg13g2_mux2_1 _646_ (.A0(net193),
    .A1(net3),
    .S(net166),
    .X(_126_));
 sg13g2_mux2_1 _647_ (.A0(spi_clk_sync),
    .A1(net168),
    .S(net167),
    .X(_127_));
 sg13g2_mux2_1 _648_ (.A0(net168),
    .A1(net4),
    .S(net167),
    .X(_128_));
 sg13g2_mux2_1 _649_ (.A0(net204),
    .A1(spi_clk_sync),
    .S(net164),
    .X(_129_));
 sg13g2_mux2_1 _650_ (.A0(net196),
    .A1(net5),
    .S(net167),
    .X(_130_));
 sg13g2_mux2_1 _651_ (.A0(cpol_sync),
    .A1(net117),
    .S(net167),
    .X(_131_));
 sg13g2_dfrbp_1 _652_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net147),
    .D(_022_),
    .Q_N(_379_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[0] ));
 sg13g2_dfrbp_1 _653_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net147),
    .D(_023_),
    .Q_N(_378_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ));
 sg13g2_dfrbp_1 _654_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net147),
    .D(net182),
    .Q_N(_377_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[2] ));
 sg13g2_dfrbp_1 _655_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net147),
    .D(net245),
    .Q_N(_376_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ));
 sg13g2_dfrbp_1 _656_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net148),
    .D(_026_),
    .Q_N(_375_),
    .Q(\spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_dfrbp_1 _657_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net149),
    .D(_027_),
    .Q_N(_374_),
    .Q(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_dfrbp_1 _658_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net145),
    .D(_028_),
    .Q_N(_373_),
    .Q(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_dfrbp_1 _659_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net145),
    .D(_029_),
    .Q_N(_004_),
    .Q(\spi_wrapper_i.reg_addr[2] ));
 sg13g2_dfrbp_1 _660_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net149),
    .D(_030_),
    .Q_N(_372_),
    .Q(\spi_wrapper_i.reg_addr[3] ));
 sg13g2_dfrbp_1 _661_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net149),
    .D(_031_),
    .Q_N(_371_),
    .Q(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_dfrbp_1 _662_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net149),
    .D(net186),
    .Q_N(_370_),
    .Q(\spi_wrapper_i.reg_data_o[0] ));
 sg13g2_dfrbp_1 _663_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net146),
    .D(_033_),
    .Q_N(_369_),
    .Q(\spi_wrapper_i.reg_data_o[1] ));
 sg13g2_dfrbp_1 _664_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net145),
    .D(_034_),
    .Q_N(_368_),
    .Q(\spi_wrapper_i.reg_data_o[2] ));
 sg13g2_dfrbp_1 _665_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net144),
    .D(_035_),
    .Q_N(_367_),
    .Q(\spi_wrapper_i.reg_data_o[3] ));
 sg13g2_dfrbp_1 _666_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net144),
    .D(_036_),
    .Q_N(_366_),
    .Q(\spi_wrapper_i.reg_data_o[4] ));
 sg13g2_dfrbp_1 _667_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net144),
    .D(net200),
    .Q_N(_365_),
    .Q(\spi_wrapper_i.reg_data_o[5] ));
 sg13g2_dfrbp_1 _668_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net143),
    .D(_038_),
    .Q_N(_364_),
    .Q(\spi_wrapper_i.reg_data_o[6] ));
 sg13g2_dfrbp_1 _669_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net145),
    .D(net212),
    .Q_N(_363_),
    .Q(\spi_wrapper_i.reg_data_o[7] ));
 sg13g2_dfrbp_1 _670_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net159),
    .D(net36),
    .Q_N(_006_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ));
 sg13g2_dfrbp_1 _671_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net159),
    .D(net29),
    .Q_N(_008_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ));
 sg13g2_dfrbp_1 _672_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net159),
    .D(net25),
    .Q_N(_010_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ));
 sg13g2_dfrbp_1 _673_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net159),
    .D(net34),
    .Q_N(_012_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_dfrbp_1 _674_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net158),
    .D(net27),
    .Q_N(_014_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_dfrbp_1 _675_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net158),
    .D(net23),
    .Q_N(_016_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ));
 sg13g2_dfrbp_1 _676_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net158),
    .D(net42),
    .Q_N(_018_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_dfrbp_1 _677_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net149),
    .D(net40),
    .Q_N(_362_),
    .Q(spi_miso));
 sg13g2_dfrbp_1 _678_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net160),
    .D(net101),
    .Q_N(_361_),
    .Q(\config_regs[56] ));
 sg13g2_dfrbp_1 _679_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net156),
    .D(net103),
    .Q_N(_360_),
    .Q(\config_regs[57] ));
 sg13g2_dfrbp_1 _680_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net156),
    .D(net52),
    .Q_N(_359_),
    .Q(\config_regs[58] ));
 sg13g2_dfrbp_1 _681_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net154),
    .D(net46),
    .Q_N(_358_),
    .Q(\config_regs[59] ));
 sg13g2_dfrbp_1 _682_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net144),
    .D(_052_),
    .Q_N(_357_),
    .Q(\config_regs[60] ));
 sg13g2_dfrbp_1 _683_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net144),
    .D(net192),
    .Q_N(_356_),
    .Q(\config_regs[61] ));
 sg13g2_dfrbp_1 _684_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net154),
    .D(net97),
    .Q_N(_355_),
    .Q(\config_regs[62] ));
 sg13g2_dfrbp_1 _685_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net145),
    .D(net173),
    .Q_N(_354_),
    .Q(\config_regs[63] ));
 sg13g2_dfrbp_1 _686_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net150),
    .D(_056_),
    .Q_N(_353_),
    .Q(spi_mosi_sync));
 sg13g2_dfrbp_1 _687_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net147),
    .D(_057_),
    .Q_N(_352_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ));
 sg13g2_dfrbp_1 _688_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net143),
    .D(_058_),
    .Q_N(_351_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ));
 sg13g2_dfrbp_1 _689_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net143),
    .D(_059_),
    .Q_N(_350_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ));
 sg13g2_dfrbp_1 _690_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net143),
    .D(_060_),
    .Q_N(_349_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ));
 sg13g2_dfrbp_1 _691_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net143),
    .D(_061_),
    .Q_N(_348_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ));
 sg13g2_dfrbp_1 _692_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net143),
    .D(_062_),
    .Q_N(_347_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ));
 sg13g2_dfrbp_1 _693_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net143),
    .D(_063_),
    .Q_N(_346_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ));
 sg13g2_dfrbp_1 _694_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net143),
    .D(_064_),
    .Q_N(_345_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ));
 sg13g2_dfrbp_1 _695_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net148),
    .D(_065_),
    .Q_N(_344_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_dfrbp_1 _696_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net162),
    .D(net229),
    .Q_N(_343_),
    .Q(\config_regs[32] ));
 sg13g2_dfrbp_1 _697_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net160),
    .D(_067_),
    .Q_N(_342_),
    .Q(\config_regs[33] ));
 sg13g2_dfrbp_1 _698_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net156),
    .D(net221),
    .Q_N(_341_),
    .Q(\config_regs[34] ));
 sg13g2_dfrbp_1 _699_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net155),
    .D(net231),
    .Q_N(_340_),
    .Q(\config_regs[35] ));
 sg13g2_dfrbp_1 _700_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net163),
    .D(net66),
    .Q_N(_339_),
    .Q(\config_regs[36] ));
 sg13g2_dfrbp_1 _701_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net152),
    .D(net236),
    .Q_N(_338_),
    .Q(\config_regs[37] ));
 sg13g2_dfrbp_1 _702_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net154),
    .D(net219),
    .Q_N(_337_),
    .Q(\config_regs[38] ));
 sg13g2_dfrbp_1 _703_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net153),
    .D(_073_),
    .Q_N(_336_),
    .Q(\config_regs[39] ));
 sg13g2_dfrbp_1 _704_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net160),
    .D(net217),
    .Q_N(_335_),
    .Q(\config_regs[40] ));
 sg13g2_dfrbp_1 _705_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net160),
    .D(net82),
    .Q_N(_334_),
    .Q(\config_regs[41] ));
 sg13g2_dfrbp_1 _706_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net156),
    .D(net198),
    .Q_N(_333_),
    .Q(\config_regs[42] ));
 sg13g2_dfrbp_1 _707_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net155),
    .D(net188),
    .Q_N(_332_),
    .Q(\config_regs[43] ));
 sg13g2_dfrbp_1 _708_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net153),
    .D(_078_),
    .Q_N(_331_),
    .Q(\config_regs[44] ));
 sg13g2_dfrbp_1 _709_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net144),
    .D(net76),
    .Q_N(_330_),
    .Q(\config_regs[45] ));
 sg13g2_dfrbp_1 _710_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net154),
    .D(net50),
    .Q_N(_329_),
    .Q(\config_regs[46] ));
 sg13g2_dfrbp_1 _711_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net153),
    .D(net87),
    .Q_N(_328_),
    .Q(\config_regs[47] ));
 sg13g2_dfrbp_1 _712_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net160),
    .D(net48),
    .Q_N(_327_),
    .Q(\config_regs[24] ));
 sg13g2_dfrbp_1 _713_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net160),
    .D(net54),
    .Q_N(_326_),
    .Q(\config_regs[25] ));
 sg13g2_dfrbp_1 _714_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net156),
    .D(net175),
    .Q_N(_325_),
    .Q(\config_regs[26] ));
 sg13g2_dfrbp_1 _715_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net155),
    .D(net91),
    .Q_N(_324_),
    .Q(\config_regs[27] ));
 sg13g2_dfrbp_1 _716_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net153),
    .D(_086_),
    .Q_N(_323_),
    .Q(\config_regs[28] ));
 sg13g2_dfrbp_1 _717_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net152),
    .D(net60),
    .Q_N(_322_),
    .Q(\config_regs[29] ));
 sg13g2_dfrbp_1 _718_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net154),
    .D(net56),
    .Q_N(_321_),
    .Q(\config_regs[30] ));
 sg13g2_dfrbp_1 _719_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net144),
    .D(net95),
    .Q_N(_320_),
    .Q(\config_regs[31] ));
 sg13g2_dfrbp_1 _720_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net153),
    .D(net105),
    .Q_N(_319_),
    .Q(\config_regs[48] ));
 sg13g2_dfrbp_1 _721_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net156),
    .D(net123),
    .Q_N(_318_),
    .Q(\config_regs[49] ));
 sg13g2_dfrbp_1 _722_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net156),
    .D(net190),
    .Q_N(_317_),
    .Q(\config_regs[50] ));
 sg13g2_dfrbp_1 _723_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net154),
    .D(net112),
    .Q_N(_316_),
    .Q(\config_regs[51] ));
 sg13g2_dfrbp_1 _724_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net152),
    .D(_094_),
    .Q_N(_315_),
    .Q(\config_regs[52] ));
 sg13g2_dfrbp_1 _725_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net152),
    .D(net195),
    .Q_N(_314_),
    .Q(\config_regs[53] ));
 sg13g2_dfrbp_1 _726_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net152),
    .D(net99),
    .Q_N(_313_),
    .Q(\config_regs[54] ));
 sg13g2_dfrbp_1 _727_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net153),
    .D(net184),
    .Q_N(_312_),
    .Q(\config_regs[55] ));
 sg13g2_dfrbp_1 _728_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net160),
    .D(net89),
    .Q_N(_311_),
    .Q(\config_regs[16] ));
 sg13g2_dfrbp_1 _729_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net161),
    .D(net171),
    .Q_N(_310_),
    .Q(\config_regs[17] ));
 sg13g2_dfrbp_1 _730_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net157),
    .D(net62),
    .Q_N(_309_),
    .Q(\config_regs[18] ));
 sg13g2_dfrbp_1 _731_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net155),
    .D(net72),
    .Q_N(_308_),
    .Q(\config_regs[19] ));
 sg13g2_dfrbp_1 _732_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net152),
    .D(_102_),
    .Q_N(_307_),
    .Q(\config_regs[20] ));
 sg13g2_dfrbp_1 _733_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net144),
    .D(net110),
    .Q_N(_306_),
    .Q(\config_regs[21] ));
 sg13g2_dfrbp_1 _734_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net154),
    .D(net177),
    .Q_N(_305_),
    .Q(\config_regs[22] ));
 sg13g2_dfrbp_1 _735_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net145),
    .D(net74),
    .Q_N(_304_),
    .Q(\config_regs[23] ));
 sg13g2_dfrbp_1 _736_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net160),
    .D(net116),
    .Q_N(_303_),
    .Q(\config_regs[8] ));
 sg13g2_dfrbp_1 _737_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net157),
    .D(net93),
    .Q_N(_302_),
    .Q(\config_regs[9] ));
 sg13g2_dfrbp_1 _738_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net156),
    .D(net179),
    .Q_N(_301_),
    .Q(\config_regs[10] ));
 sg13g2_dfrbp_1 _739_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net155),
    .D(net202),
    .Q_N(_300_),
    .Q(\config_regs[11] ));
 sg13g2_dfrbp_1 _740_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net152),
    .D(_110_),
    .Q_N(_299_),
    .Q(\config_regs[12] ));
 sg13g2_dfrbp_1 _741_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net152),
    .D(net214),
    .Q_N(_298_),
    .Q(\config_regs[13] ));
 sg13g2_dfrbp_1 _742_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net154),
    .D(net208),
    .Q_N(_297_),
    .Q(\config_regs[14] ));
 sg13g2_dfrbp_1 _743_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net153),
    .D(net80),
    .Q_N(_296_),
    .Q(\config_regs[15] ));
 sg13g2_dfrbp_1 _744_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net158),
    .D(net85),
    .Q_N(_005_),
    .Q(\config_regs[0] ));
 sg13g2_dfrbp_1 _745_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net158),
    .D(net120),
    .Q_N(_007_),
    .Q(\config_regs[1] ));
 sg13g2_dfrbp_1 _746_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net158),
    .D(net68),
    .Q_N(_009_),
    .Q(\config_regs[2] ));
 sg13g2_dfrbp_1 _747_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net158),
    .D(net108),
    .Q_N(_011_),
    .Q(\config_regs[3] ));
 sg13g2_dfrbp_1 _748_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net150),
    .D(_118_),
    .Q_N(_013_),
    .Q(\config_regs[4] ));
 sg13g2_dfrbp_1 _749_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net149),
    .D(net58),
    .Q_N(_015_),
    .Q(\config_regs[5] ));
 sg13g2_dfrbp_1 _750_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net150),
    .D(net78),
    .Q_N(_017_),
    .Q(\config_regs[6] ));
 sg13g2_dfrbp_1 _751_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net150),
    .D(net64),
    .Q_N(_019_),
    .Q(\config_regs[7] ));
 sg13g2_dfrbp_1 _752_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net161),
    .D(_122_),
    .Q_N(_295_),
    .Q(\synchronizer_spi_mode_cpol.data_sync[1] ));
 sg13g2_dfrbp_1 _753_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net161),
    .D(_123_),
    .Q_N(_294_),
    .Q(cpha_sync));
 sg13g2_dfrbp_1 _754_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net161),
    .D(_124_),
    .Q_N(_293_),
    .Q(\synchronizer_spi_mode_cpha.data_sync[1] ));
 sg13g2_dfrbp_1 _755_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net148),
    .D(_125_),
    .Q_N(uio_oe[3]),
    .Q(spi_cs_n_sync));
 sg13g2_dfrbp_1 _756_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net149),
    .D(_126_),
    .Q_N(_292_),
    .Q(\synchronizer_spi_cs_n_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _757_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net158),
    .D(net169),
    .Q_N(_291_),
    .Q(spi_clk_sync));
 sg13g2_dfrbp_1 _758_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net159),
    .D(_128_),
    .Q_N(_290_),
    .Q(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _759_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net148),
    .D(net205),
    .Q_N(_289_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_dfrbp_1 _760_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net149),
    .D(_130_),
    .Q_N(_288_),
    .Q(\synchronizer_spi_mosi_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _761_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net161),
    .D(net118),
    .Q_N(_287_),
    .Q(cpol_sync));
 sg13g2_dfrbp_1 _762_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net148),
    .D(net21),
    .Q_N(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .Q(_020_));
 sg13g2_dfrbp_1 _763_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net147),
    .D(net38),
    .Q_N(_380_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[1] ));
 sg13g2_dfrbp_1 _764_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net147),
    .D(_001_),
    .Q_N(_381_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_dfrbp_1 _765_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net148),
    .D(net32),
    .Q_N(_382_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_dfrbp_1 _766_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net147),
    .D(_003_),
    .Q_N(_286_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_tielo tt_um_calonso88_spi_test_7 (.L_LO(net7));
 sg13g2_tielo tt_um_calonso88_spi_test_8 (.L_LO(net8));
 sg13g2_tielo tt_um_calonso88_spi_test_9 (.L_LO(net9));
 sg13g2_tielo tt_um_calonso88_spi_test_10 (.L_LO(net10));
 sg13g2_tielo tt_um_calonso88_spi_test_11 (.L_LO(net11));
 sg13g2_tielo tt_um_calonso88_spi_test_12 (.L_LO(net12));
 sg13g2_tielo tt_um_calonso88_spi_test_13 (.L_LO(net13));
 sg13g2_tielo tt_um_calonso88_spi_test_14 (.L_LO(net14));
 sg13g2_tielo tt_um_calonso88_spi_test_15 (.L_LO(net15));
 sg13g2_tielo tt_um_calonso88_spi_test_16 (.L_LO(net16));
 sg13g2_tielo tt_um_calonso88_spi_test_17 (.L_LO(net17));
 sg13g2_tielo tt_um_calonso88_spi_test_18 (.L_LO(net18));
 sg13g2_tielo tt_um_calonso88_spi_test_19 (.L_LO(net19));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _781_ (.A(spi_miso),
    .X(uio_out[3]));
 sg13g2_buf_1 _782_ (.A(\config_regs[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _783_ (.A(\config_regs[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _784_ (.A(\config_regs[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _785_ (.A(\config_regs[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _786_ (.A(\config_regs[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _787_ (.A(\config_regs[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _788_ (.A(\config_regs[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _789_ (.A(\config_regs[7] ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout125 (.A(_155_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net128),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_152_),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_149_));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_193_));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(_188_));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_185_));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(_198_));
 sg13g2_buf_2 fanout134 (.A(net211),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net239));
 sg13g2_buf_2 fanout136 (.A(\spi_wrapper_i.reg_data_o[5] ),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net65));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net243));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net238));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(net227));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(\spi_wrapper_i.reg_data_o[0] ));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_004_));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(net146));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net146));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net146));
 sg13g2_buf_2 fanout146 (.A(net151),
    .X(net146));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(net148));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net151));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net151));
 sg13g2_buf_2 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(rst_n),
    .X(net151));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(net153));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(net163));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(net157));
 sg13g2_buf_2 fanout155 (.A(net157),
    .X(net155));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net157));
 sg13g2_buf_2 fanout157 (.A(net163),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net162));
 sg13g2_buf_2 fanout159 (.A(net162),
    .X(net159));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net161));
 sg13g2_buf_2 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(rst_n),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net166),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net167));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(ena));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[6]),
    .X(net5));
 sg13g2_tielo tt_um_calonso88_spi_test_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold2 (.A(_021_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold3 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold4 (.A(_045_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold5 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold6 (.A(_042_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold7 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold8 (.A(_044_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold9 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold10 (.A(_041_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold11 (.A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold12 (.A(_156_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold13 (.A(_002_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold14 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold15 (.A(_043_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold16 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold17 (.A(_040_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold18 (.A(\spi_wrapper_i.spi_reg_inst.reg_rw ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold19 (.A(_000_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold20 (.A(spi_miso),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold21 (.A(_047_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold22 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold23 (.A(_046_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold24 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold25 (.A(\spi_wrapper_i.spi_reg_inst.state[2] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold26 (.A(\config_regs[59] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold27 (.A(_051_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold28 (.A(\config_regs[24] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold29 (.A(_082_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold30 (.A(\config_regs[46] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold31 (.A(_080_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold32 (.A(\config_regs[58] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold33 (.A(_050_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold34 (.A(\config_regs[25] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold35 (.A(_083_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold36 (.A(\config_regs[30] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold37 (.A(_088_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold38 (.A(\config_regs[5] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold39 (.A(_119_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold40 (.A(\config_regs[29] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold41 (.A(_087_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold42 (.A(\config_regs[18] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold43 (.A(_100_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold44 (.A(\config_regs[7] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold45 (.A(_121_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold46 (.A(\spi_wrapper_i.reg_data_o[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold47 (.A(_070_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold48 (.A(\config_regs[2] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold49 (.A(_116_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold50 (.A(\config_regs[28] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold51 (.A(\config_regs[44] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold52 (.A(\config_regs[19] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold53 (.A(_101_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold54 (.A(\config_regs[23] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold55 (.A(_105_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold56 (.A(\config_regs[45] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold57 (.A(_079_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold58 (.A(\config_regs[6] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold59 (.A(_120_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold60 (.A(\config_regs[15] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold61 (.A(_113_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold62 (.A(\config_regs[41] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold63 (.A(_075_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold64 (.A(\config_regs[12] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold65 (.A(\config_regs[0] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold66 (.A(_114_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold67 (.A(\config_regs[47] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold68 (.A(_081_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold69 (.A(\config_regs[16] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold70 (.A(_098_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold71 (.A(\config_regs[27] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold72 (.A(_085_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold73 (.A(\config_regs[9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold74 (.A(_107_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold75 (.A(\config_regs[31] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold76 (.A(_089_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold77 (.A(\config_regs[62] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold78 (.A(_054_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold79 (.A(\config_regs[54] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold80 (.A(_096_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold81 (.A(\config_regs[56] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold82 (.A(_048_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold83 (.A(\config_regs[57] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold84 (.A(_049_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold85 (.A(\config_regs[48] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold86 (.A(_090_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold87 (.A(\config_regs[60] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold88 (.A(\config_regs[3] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold89 (.A(_117_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold90 (.A(\config_regs[21] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold91 (.A(_103_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold92 (.A(\config_regs[51] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold93 (.A(_093_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold94 (.A(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold95 (.A(\config_regs[52] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold96 (.A(\config_regs[8] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold97 (.A(_106_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold98 (.A(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold99 (.A(_131_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold100 (.A(\config_regs[1] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold101 (.A(_115_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold102 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold103 (.A(\config_regs[49] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold104 (.A(_091_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold105 (.A(\config_regs[20] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold106 (.A(\synchronizer_spi_clk_inst.data_sync[1] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold107 (.A(_127_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold108 (.A(\config_regs[17] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold109 (.A(_099_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold110 (.A(\config_regs[63] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold111 (.A(_055_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold112 (.A(\config_regs[26] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold113 (.A(_084_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold114 (.A(\config_regs[22] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold115 (.A(_104_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold116 (.A(\config_regs[10] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold117 (.A(_108_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold118 (.A(\config_regs[4] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold119 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[2] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold120 (.A(_024_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold121 (.A(\config_regs[55] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold122 (.A(_097_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold123 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold124 (.A(_032_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold125 (.A(\config_regs[43] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold126 (.A(_077_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold127 (.A(\config_regs[50] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold128 (.A(_092_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold129 (.A(\config_regs[61] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold130 (.A(_053_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold131 (.A(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold132 (.A(\config_regs[53] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold133 (.A(_095_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold134 (.A(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold135 (.A(\config_regs[42] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold136 (.A(_076_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold137 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold138 (.A(_037_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold139 (.A(\config_regs[11] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold140 (.A(_109_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold141 (.A(spi_mosi_sync),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold142 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold143 (.A(_129_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold144 (.A(spi_cs_n_sync),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold145 (.A(\config_regs[14] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold146 (.A(_112_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold147 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold148 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold149 (.A(\spi_wrapper_i.reg_data_o[7] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold150 (.A(_039_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold151 (.A(\config_regs[13] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold152 (.A(_111_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold153 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold154 (.A(\config_regs[40] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold155 (.A(_074_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold156 (.A(\config_regs[38] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold157 (.A(_072_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold158 (.A(\config_regs[34] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold159 (.A(_068_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold160 (.A(\spi_wrapper_i.reg_addr[0] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold161 (.A(cpha_sync),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold162 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold163 (.A(\config_regs[39] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold164 (.A(\spi_wrapper_i.reg_addr[1] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold165 (.A(\spi_wrapper_i.reg_data_o[1] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold166 (.A(\config_regs[32] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold167 (.A(_066_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold168 (.A(\config_regs[35] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold169 (.A(_069_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold170 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold171 (.A(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold172 (.A(\spi_wrapper_i.reg_data_o_vld ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold173 (.A(\config_regs[37] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold174 (.A(_071_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold175 (.A(\config_regs[33] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold176 (.A(\spi_wrapper_i.reg_data_o[2] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold177 (.A(\spi_wrapper_i.reg_data_o[6] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold178 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[0] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold179 (.A(_166_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold180 (.A(\spi_wrapper_i.reg_addr[3] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold181 (.A(\spi_wrapper_i.reg_data_o[3] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold182 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold183 (.A(_025_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold184 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ),
    .X(net246));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_4 FILLER_12_266 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_278 ();
 sg13g2_fill_2 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_4 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_decap_4 FILLER_13_300 ();
 sg13g2_fill_2 FILLER_13_304 ();
 sg13g2_decap_4 FILLER_13_315 ();
 sg13g2_fill_2 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_4 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_193 ();
 sg13g2_fill_1 FILLER_14_195 ();
 sg13g2_decap_4 FILLER_14_259 ();
 sg13g2_decap_4 FILLER_14_315 ();
 sg13g2_decap_4 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_177 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_decap_4 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_4 FILLER_16_140 ();
 sg13g2_decap_4 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_184 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_1 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_167 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_fill_2 FILLER_17_371 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_4 FILLER_18_98 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_decap_8 FILLER_18_121 ();
 sg13g2_decap_4 FILLER_18_128 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_decap_4 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_349 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_77 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_fill_2 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_decap_4 FILLER_19_339 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_359 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_decap_4 FILLER_20_167 ();
 sg13g2_decap_4 FILLER_20_202 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_287 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_decap_4 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_decap_4 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_192 ();
 sg13g2_decap_4 FILLER_21_246 ();
 sg13g2_decap_4 FILLER_21_295 ();
 sg13g2_decap_4 FILLER_21_308 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_4 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_85 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_fill_2 FILLER_22_99 ();
 sg13g2_fill_1 FILLER_22_101 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_decap_4 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_decap_8 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_285 ();
 sg13g2_decap_4 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_fill_2 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_decap_4 FILLER_23_93 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_152 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_1 FILLER_23_251 ();
 sg13g2_decap_4 FILLER_23_276 ();
 sg13g2_decap_4 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_351 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_106 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_decap_4 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_decap_4 FILLER_25_97 ();
 sg13g2_fill_2 FILLER_25_111 ();
 sg13g2_fill_1 FILLER_25_113 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_decap_4 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_309 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_decap_4 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_101 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_228 ();
 sg13g2_decap_4 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_2 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_decap_4 FILLER_27_106 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_decap_8 FILLER_28_155 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_243 ();
 sg13g2_decap_4 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_47 ();
 sg13g2_fill_1 FILLER_29_51 ();
 sg13g2_decap_4 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_337 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_4 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_decap_4 FILLER_30_249 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_155 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_312 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_87 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_183 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_2 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_decap_8 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_181 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_332 ();
 sg13g2_fill_2 FILLER_33_355 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_32 ();
 sg13g2_decap_8 FILLER_34_48 ();
 sg13g2_decap_8 FILLER_34_55 ();
 sg13g2_decap_4 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_151 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_decap_8 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_4 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_decap_4 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_153 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_decap_4 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_decap_4 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_163 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_170 ();
 sg13g2_decap_4 FILLER_37_207 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule
