module tt_um_digital_clock_example (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire net25;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire \desk_clock.clk_gen_inst.i_refclk ;
 wire \desk_clock.clk_gen_inst.refclk_div[0] ;
 wire \desk_clock.clk_gen_inst.refclk_div[10] ;
 wire \desk_clock.clk_gen_inst.refclk_div[11] ;
 wire \desk_clock.clk_gen_inst.refclk_div[12] ;
 wire \desk_clock.clk_gen_inst.refclk_div[13] ;
 wire \desk_clock.clk_gen_inst.refclk_div[14] ;
 wire \desk_clock.clk_gen_inst.refclk_div[1] ;
 wire \desk_clock.clk_gen_inst.refclk_div[2] ;
 wire \desk_clock.clk_gen_inst.refclk_div[3] ;
 wire \desk_clock.clk_gen_inst.refclk_div[4] ;
 wire \desk_clock.clk_gen_inst.refclk_div[5] ;
 wire \desk_clock.clk_gen_inst.refclk_div[6] ;
 wire \desk_clock.clk_gen_inst.refclk_div[7] ;
 wire \desk_clock.clk_gen_inst.refclk_div[8] ;
 wire \desk_clock.clk_gen_inst.refclk_div[9] ;
 wire \desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold ;
 wire \desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold ;
 wire \desk_clock.clk_hours[0] ;
 wire \desk_clock.clk_hours[1] ;
 wire \desk_clock.clk_hours[2] ;
 wire \desk_clock.clk_hours[3] ;
 wire \desk_clock.clk_hours[4] ;
 wire \desk_clock.clk_minutes[0] ;
 wire \desk_clock.clk_minutes[1] ;
 wire \desk_clock.clk_minutes[2] ;
 wire \desk_clock.clk_minutes[3] ;
 wire \desk_clock.clk_minutes[4] ;
 wire \desk_clock.clk_minutes[5] ;
 wire \desk_clock.clk_seconds[0] ;
 wire \desk_clock.clk_seconds[1] ;
 wire \desk_clock.clk_seconds[2] ;
 wire \desk_clock.clk_seconds[3] ;
 wire \desk_clock.clk_seconds[4] ;
 wire \desk_clock.clk_seconds[5] ;
 wire \desk_clock.display_control_inst.display_update ;
 wire \desk_clock.display_control_inst.o_write_config ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[0] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[1] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[2] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[3] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[4] ;
 wire \desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[0] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[10] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[11] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[12] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[13] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[14] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[15] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[1] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[2] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[3] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[4] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[5] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[6] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[7] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[8] ;
 wire \desk_clock.display_inst.disp_driver.data_reg[9] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[0] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[1] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[2] ;
 wire \desk_clock.display_inst.disp_driver.i_addr[3] ;
 wire \desk_clock.display_inst.disp_driver.i_data[0] ;
 wire \desk_clock.display_inst.disp_driver.i_data[1] ;
 wire \desk_clock.display_inst.disp_driver.i_data[2] ;
 wire \desk_clock.display_inst.disp_driver.i_data[3] ;
 wire \desk_clock.display_inst.disp_driver.i_data[4] ;
 wire \desk_clock.display_inst.disp_driver.i_data[7] ;
 wire \desk_clock.display_inst.disp_driver.o_serial_clk ;
 wire \desk_clock.display_inst.disp_driver.o_serial_load ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[0] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[1] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[2] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[3] ;
 wire \desk_clock.display_inst.disp_driver.transfer_state[4] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[0] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[1] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[2] ;
 wire \desk_clock.display_inst.display_settings.transfer_state[3] ;
 wire \desk_clock.display_inst.display_settings.write_config ;
 wire \desk_clock.display_inst.state[0] ;
 wire \desk_clock.display_inst.state[1] ;
 wire \desk_clock.display_inst.state[2] ;
 wire \desk_clock.display_inst.state[3] ;
 wire \desk_clock.input_debounce.en_12h_mode_reg[0] ;
 wire \desk_clock.input_debounce.en_12h_mode_reg[1] ;
 wire \desk_clock.input_debounce.en_12h_mode_reg[2] ;
 wire \desk_clock.input_debounce.en_12h_mode_reg[3] ;
 wire \desk_clock.input_debounce.en_12h_mode_reg[4] ;
 wire \desk_clock.input_debounce.en_12h_mode_reg[5] ;
 wire \desk_clock.input_debounce.fast_set_reg[0] ;
 wire \desk_clock.input_debounce.fast_set_reg[1] ;
 wire \desk_clock.input_debounce.fast_set_reg[2] ;
 wire \desk_clock.input_debounce.fast_set_reg[3] ;
 wire \desk_clock.input_debounce.fast_set_reg[4] ;
 wire \desk_clock.input_debounce.fast_set_reg[5] ;
 wire \desk_clock.input_debounce.set_hours_reg[0] ;
 wire \desk_clock.input_debounce.set_hours_reg[1] ;
 wire \desk_clock.input_debounce.set_hours_reg[2] ;
 wire \desk_clock.input_debounce.set_hours_reg[3] ;
 wire \desk_clock.input_debounce.set_hours_reg[4] ;
 wire \desk_clock.input_debounce.set_hours_reg[5] ;
 wire \desk_clock.input_debounce.set_minutes_reg[0] ;
 wire \desk_clock.input_debounce.set_minutes_reg[1] ;
 wire \desk_clock.input_debounce.set_minutes_reg[2] ;
 wire \desk_clock.input_debounce.set_minutes_reg[3] ;
 wire \desk_clock.input_debounce.set_minutes_reg[4] ;
 wire \desk_clock.input_debounce.set_minutes_reg[5] ;
 wire \desk_clock.refclk_sync_inst.refclk_sync_reg[0] ;
 wire net148;
 wire net149;
 wire net7;
 wire clk_regs;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;

 sg13g2_inv_1 _0810_ (.Y(_0130_),
    .A(net312));
 sg13g2_inv_1 _0811_ (.Y(_0131_),
    .A(net304));
 sg13g2_inv_1 _0812_ (.Y(_0132_),
    .A(net326));
 sg13g2_inv_1 _0813_ (.Y(_0133_),
    .A(net358));
 sg13g2_inv_1 _0814_ (.Y(_0134_),
    .A(net228));
 sg13g2_inv_1 _0815_ (.Y(_0135_),
    .A(net201));
 sg13g2_inv_1 _0816_ (.Y(_0136_),
    .A(net243));
 sg13g2_inv_1 _0817_ (.Y(_0137_),
    .A(net5));
 sg13g2_inv_1 _0818_ (.Y(_0138_),
    .A(net321));
 sg13g2_inv_1 _0819_ (.Y(_0139_),
    .A(net281));
 sg13g2_inv_1 _0820_ (.Y(_0140_),
    .A(net270));
 sg13g2_inv_1 _0821_ (.Y(_0141_),
    .A(net265));
 sg13g2_inv_1 _0822_ (.Y(_0142_),
    .A(net223));
 sg13g2_inv_1 _0823_ (.Y(_0143_),
    .A(net4));
 sg13g2_inv_1 _0824_ (.Y(_0144_),
    .A(net329));
 sg13g2_inv_1 _0825_ (.Y(_0145_),
    .A(net309));
 sg13g2_inv_1 _0826_ (.Y(_0146_),
    .A(net293));
 sg13g2_inv_1 _0827_ (.Y(_0147_),
    .A(net256));
 sg13g2_inv_1 _0828_ (.Y(_0148_),
    .A(net267));
 sg13g2_inv_1 _0829_ (.Y(_0149_),
    .A(net3));
 sg13g2_inv_1 _0830_ (.Y(_0150_),
    .A(net253));
 sg13g2_inv_1 _0831_ (.Y(_0151_),
    .A(net294));
 sg13g2_inv_1 _0832_ (.Y(_0152_),
    .A(net289));
 sg13g2_inv_1 _0833_ (.Y(_0153_),
    .A(net307));
 sg13g2_inv_1 _0834_ (.Y(_0154_),
    .A(net213));
 sg13g2_inv_1 _0835_ (.Y(_0155_),
    .A(net2));
 sg13g2_inv_1 _0836_ (.Y(_0156_),
    .A(net320));
 sg13g2_inv_1 _0837_ (.Y(_0157_),
    .A(net298));
 sg13g2_inv_1 _0838_ (.Y(_0158_),
    .A(net209));
 sg13g2_inv_1 _0839_ (.Y(_0159_),
    .A(net316));
 sg13g2_inv_1 _0840_ (.Y(_0160_),
    .A(net403));
 sg13g2_inv_1 _0841_ (.Y(_0161_),
    .A(\desk_clock.clk_hours[2] ));
 sg13g2_inv_1 _0842_ (.Y(_0162_),
    .A(net346));
 sg13g2_inv_1 _0843_ (.Y(_0163_),
    .A(net376));
 sg13g2_inv_1 _0844_ (.Y(_0164_),
    .A(net287));
 sg13g2_inv_1 _0845_ (.Y(_0165_),
    .A(net179));
 sg13g2_inv_1 _0846_ (.Y(_0166_),
    .A(net291));
 sg13g2_inv_1 _0847_ (.Y(_0167_),
    .A(net302));
 sg13g2_inv_1 _0848_ (.Y(_0168_),
    .A(net279));
 sg13g2_inv_1 _0849_ (.Y(_0169_),
    .A(net277));
 sg13g2_inv_1 _0850_ (.Y(_0170_),
    .A(net273));
 sg13g2_inv_1 _0851_ (.Y(_0171_),
    .A(net260));
 sg13g2_inv_1 _0852_ (.Y(_0172_),
    .A(net232));
 sg13g2_inv_1 _0853_ (.Y(_0173_),
    .A(net258));
 sg13g2_inv_1 _0854_ (.Y(_0174_),
    .A(net268));
 sg13g2_inv_1 _0855_ (.Y(_0175_),
    .A(net241));
 sg13g2_inv_1 _0856_ (.Y(_0176_),
    .A(net271));
 sg13g2_inv_1 _0857_ (.Y(_0177_),
    .A(net198));
 sg13g2_or3_1 _0858_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[3] ),
    .B(\desk_clock.display_inst.disp_driver.transfer_state[2] ),
    .C(\desk_clock.display_inst.disp_driver.transfer_state[1] ),
    .X(_0178_));
 sg13g2_nor2_1 _0859_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[0] ),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_nor3_1 _0860_ (.A(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .B(\desk_clock.display_inst.disp_driver.transfer_state[0] ),
    .C(_0178_),
    .Y(_0180_));
 sg13g2_nand2b_1 _0861_ (.Y(_0181_),
    .B(_0179_),
    .A_N(\desk_clock.display_inst.disp_driver.transfer_state[4] ));
 sg13g2_xor2_1 _0862_ (.B(_0179_),
    .A(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .X(\desk_clock.display_inst.disp_driver.o_serial_load ));
 sg13g2_nor2_1 _0863_ (.A(clknet_1_0__leaf_clk),
    .B(\desk_clock.display_inst.disp_driver.o_serial_load ),
    .Y(\desk_clock.display_inst.disp_driver.o_serial_clk ));
 sg13g2_and2_1 _0864_ (.A(net199),
    .B(net1),
    .X(_0008_));
 sg13g2_and2_1 _0865_ (.A(net199),
    .B(net203),
    .X(_0009_));
 sg13g2_or2_2 _0866_ (.X(_0182_),
    .B(net183),
    .A(net181));
 sg13g2_nor3_2 _0867_ (.A(net179),
    .B(net180),
    .C(net182),
    .Y(_0183_));
 sg13g2_nand2_1 _0868_ (.Y(_0184_),
    .A(net179),
    .B(net181));
 sg13g2_and2_1 _0869_ (.A(net181),
    .B(net183),
    .X(_0185_));
 sg13g2_nand3_1 _0870_ (.B(net180),
    .C(net182),
    .A(net179),
    .Y(_0186_));
 sg13g2_nor2b_2 _0871_ (.A(_0183_),
    .B_N(_0186_),
    .Y(_0187_));
 sg13g2_nand2b_2 _0872_ (.Y(_0188_),
    .B(_0186_),
    .A_N(_0183_));
 sg13g2_a21oi_2 _0873_ (.B1(net179),
    .Y(_0189_),
    .A2(net183),
    .A1(net180));
 sg13g2_a21o_1 _0874_ (.A2(net182),
    .A1(net181),
    .B1(net179),
    .X(_0190_));
 sg13g2_o21ai_1 _0875_ (.B1(\desk_clock.display_inst.state[2] ),
    .Y(_0191_),
    .A1(net180),
    .A2(net183));
 sg13g2_and2_1 _0876_ (.A(_0190_),
    .B(net177),
    .X(_0192_));
 sg13g2_nand3_1 _0877_ (.B(_0190_),
    .C(net177),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ),
    .Y(_0193_));
 sg13g2_nor2_1 _0878_ (.A(_0185_),
    .B(_0191_),
    .Y(_0194_));
 sg13g2_or3_1 _0879_ (.A(_0169_),
    .B(_0185_),
    .C(_0191_),
    .X(_0195_));
 sg13g2_and2_1 _0880_ (.A(_0182_),
    .B(_0189_),
    .X(_0196_));
 sg13g2_nand3_1 _0881_ (.B(_0182_),
    .C(_0189_),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ),
    .Y(_0197_));
 sg13g2_nand4_1 _0882_ (.B(_0193_),
    .C(_0195_),
    .A(_0187_),
    .Y(_0198_),
    .D(_0197_));
 sg13g2_or3_1 _0883_ (.A(_0168_),
    .B(_0185_),
    .C(net177),
    .X(_0199_));
 sg13g2_nand3_1 _0884_ (.B(_0190_),
    .C(net177),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ),
    .Y(_0200_));
 sg13g2_and2_1 _0885_ (.A(_0199_),
    .B(_0200_),
    .X(_0201_));
 sg13g2_nand3_1 _0886_ (.B(_0182_),
    .C(_0189_),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ),
    .Y(_0202_));
 sg13g2_nand3_1 _0887_ (.B(_0200_),
    .C(_0202_),
    .A(_0199_),
    .Y(_0203_));
 sg13g2_nor2_1 _0888_ (.A(net163),
    .B(_0203_),
    .Y(_0204_));
 sg13g2_or2_1 _0889_ (.X(_0205_),
    .B(_0203_),
    .A(net163));
 sg13g2_or3_1 _0890_ (.A(_0170_),
    .B(_0185_),
    .C(net177),
    .X(_0206_));
 sg13g2_nand3_1 _0891_ (.B(_0190_),
    .C(net177),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ),
    .Y(_0207_));
 sg13g2_nand2_1 _0892_ (.Y(_0208_),
    .A(_0206_),
    .B(_0207_));
 sg13g2_nor3_1 _0893_ (.A(net163),
    .B(_0203_),
    .C(_0208_),
    .Y(_0209_));
 sg13g2_nand3_1 _0894_ (.B(_0190_),
    .C(net177),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ),
    .Y(_0210_));
 sg13g2_or3_1 _0895_ (.A(_0167_),
    .B(_0185_),
    .C(net177),
    .X(_0211_));
 sg13g2_nand3_1 _0896_ (.B(_0182_),
    .C(_0189_),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ),
    .Y(_0212_));
 sg13g2_and4_2 _0897_ (.A(_0187_),
    .B(_0210_),
    .C(_0211_),
    .D(_0212_),
    .X(_0213_));
 sg13g2_nand4_1 _0898_ (.B(_0210_),
    .C(_0211_),
    .A(_0187_),
    .Y(_0214_),
    .D(_0212_));
 sg13g2_nor2_1 _0899_ (.A(_0188_),
    .B(_0203_),
    .Y(_0215_));
 sg13g2_nand4_1 _0900_ (.B(_0199_),
    .C(_0200_),
    .A(_0187_),
    .Y(_0216_),
    .D(_0202_));
 sg13g2_and2_1 _0901_ (.A(net163),
    .B(_0216_),
    .X(_0217_));
 sg13g2_nand2_1 _0902_ (.Y(_0218_),
    .A(net163),
    .B(_0216_));
 sg13g2_a221oi_1 _0903_ (.B2(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ),
    .C1(_0188_),
    .B1(_0194_),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ),
    .Y(_0219_),
    .A2(_0192_));
 sg13g2_inv_1 _0904_ (.Y(_0220_),
    .A(_0219_));
 sg13g2_nor4_1 _0905_ (.A(_0209_),
    .B(_0213_),
    .C(_0217_),
    .D(_0219_),
    .Y(_0221_));
 sg13g2_nand3_1 _0906_ (.B(_0182_),
    .C(_0189_),
    .A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ),
    .Y(_0222_));
 sg13g2_and4_1 _0907_ (.A(_0187_),
    .B(_0206_),
    .C(_0207_),
    .D(_0222_),
    .X(_0223_));
 sg13g2_nand4_1 _0908_ (.B(_0206_),
    .C(_0207_),
    .A(_0187_),
    .Y(_0224_),
    .D(_0222_));
 sg13g2_nand4_1 _0909_ (.B(_0214_),
    .C(_0216_),
    .A(net163),
    .Y(_0225_),
    .D(_0224_));
 sg13g2_a21oi_2 _0910_ (.B1(_0219_),
    .Y(_0226_),
    .A2(_0213_),
    .A1(_0201_));
 sg13g2_inv_1 _0911_ (.Y(_0227_),
    .A(_0226_));
 sg13g2_a21oi_1 _0912_ (.A1(_0219_),
    .A2(_0225_),
    .Y(_0228_),
    .B1(_0226_));
 sg13g2_o21ai_1 _0913_ (.B1(_0219_),
    .Y(_0229_),
    .A1(_0204_),
    .A2(_0213_));
 sg13g2_a21oi_1 _0914_ (.A1(_0216_),
    .A2(_0224_),
    .Y(_0230_),
    .B1(_0214_));
 sg13g2_a221oi_1 _0915_ (.B2(_0230_),
    .C1(_0220_),
    .B1(_0218_),
    .A1(_0205_),
    .Y(_0231_),
    .A2(_0214_));
 sg13g2_nor2_1 _0916_ (.A(_0228_),
    .B(_0231_),
    .Y(_0232_));
 sg13g2_or3_1 _0917_ (.A(_0221_),
    .B(_0228_),
    .C(_0231_),
    .X(_0233_));
 sg13g2_nor2_1 _0918_ (.A(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .B(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .Y(_0234_));
 sg13g2_nor3_2 _0919_ (.A(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .B(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .C(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .Y(_0235_));
 sg13g2_and2_1 _0920_ (.A(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .B(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .X(_0236_));
 sg13g2_nand2_1 _0921_ (.Y(_0237_),
    .A(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .B(_0236_));
 sg13g2_a21oi_1 _0922_ (.A1(net391),
    .A2(_0236_),
    .Y(_0238_),
    .B1(\desk_clock.display_inst.display_settings.transfer_state[3] ));
 sg13g2_nor2b_1 _0923_ (.A(_0235_),
    .B_N(_0238_),
    .Y(_0239_));
 sg13g2_nor2b_1 _0924_ (.A(\desk_clock.display_inst.state[3] ),
    .B_N(_0183_),
    .Y(_0240_));
 sg13g2_nor2_1 _0925_ (.A(\desk_clock.display_inst.state[3] ),
    .B(_0186_),
    .Y(_0241_));
 sg13g2_nor3_2 _0926_ (.A(_0239_),
    .B(_0240_),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_nor2b_2 _0927_ (.A(net364),
    .B_N(_0242_),
    .Y(_0243_));
 sg13g2_nand2b_2 _0928_ (.Y(_0244_),
    .B(_0242_),
    .A_N(\desk_clock.display_control_inst.o_write_config ));
 sg13g2_nand3_1 _0929_ (.B(net153),
    .C(_0243_),
    .A(net183),
    .Y(_0245_));
 sg13g2_nand2b_1 _0930_ (.Y(_0246_),
    .B(_0235_),
    .A_N(\desk_clock.display_inst.display_settings.transfer_state[3] ));
 sg13g2_nand3b_1 _0931_ (.B(_0246_),
    .C(net363),
    .Y(_0247_),
    .A_N(_0242_));
 sg13g2_xor2_1 _0932_ (.B(_0235_),
    .A(\desk_clock.display_inst.display_settings.transfer_state[3] ),
    .X(_0248_));
 sg13g2_nor3_2 _0933_ (.A(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .B(net204),
    .C(_0248_),
    .Y(_0249_));
 sg13g2_xnor2_1 _0934_ (.Y(_0250_),
    .A(_0001_),
    .B(_0234_));
 sg13g2_nor2_1 _0935_ (.A(_0248_),
    .B(_0250_),
    .Y(_0251_));
 sg13g2_a21oi_1 _0936_ (.A1(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .A2(_0249_),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_nor2_1 _0937_ (.A(_0247_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_nand2_2 _0938_ (.Y(_0254_),
    .A(net324),
    .B(_0242_));
 sg13g2_o21ai_1 _0939_ (.B1(_0254_),
    .Y(_0255_),
    .A1(_0247_),
    .A2(_0252_));
 sg13g2_inv_1 _0940_ (.Y(_0256_),
    .A(net151));
 sg13g2_o21ai_1 _0941_ (.B1(net151),
    .Y(_0257_),
    .A1(_0247_),
    .A2(_0249_));
 sg13g2_nor2_1 _0942_ (.A(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .B(_0247_),
    .Y(_0258_));
 sg13g2_inv_1 _0943_ (.Y(_0259_),
    .A(_0258_));
 sg13g2_a21oi_1 _0944_ (.A1(net179),
    .A2(_0174_),
    .Y(_0260_),
    .B1(net180));
 sg13g2_a221oi_1 _0945_ (.B2(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ),
    .C1(_0260_),
    .B1(_0196_),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ),
    .Y(_0261_),
    .A2(_0194_));
 sg13g2_nor2_1 _0946_ (.A(net182),
    .B(_0244_),
    .Y(_0262_));
 sg13g2_nor3_1 _0947_ (.A(net182),
    .B(_0244_),
    .C(_0261_),
    .Y(_0263_));
 sg13g2_nor3_1 _0948_ (.A(_0257_),
    .B(_0258_),
    .C(_0263_),
    .Y(_0264_));
 sg13g2_o21ai_1 _0949_ (.B1(net191),
    .Y(_0265_),
    .A1(net359),
    .A2(net151));
 sg13g2_a21oi_1 _0950_ (.A1(_0245_),
    .A2(_0264_),
    .Y(_0010_),
    .B1(_0265_));
 sg13g2_a21oi_1 _0951_ (.A1(_0223_),
    .A2(net152),
    .Y(_0266_),
    .B1(net348));
 sg13g2_o21ai_1 _0952_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_0223_),
    .A2(net152));
 sg13g2_o21ai_1 _0953_ (.B1(_0226_),
    .Y(_0268_),
    .A1(_0209_),
    .A2(_0213_));
 sg13g2_nand3b_1 _0954_ (.B(_0229_),
    .C(_0268_),
    .Y(_0269_),
    .A_N(_0221_));
 sg13g2_a21oi_1 _0955_ (.A1(net182),
    .A2(_0269_),
    .Y(_0270_),
    .B1(_0244_));
 sg13g2_nand2_1 _0956_ (.Y(_0271_),
    .A(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .B(_0251_));
 sg13g2_a21oi_1 _0957_ (.A1(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .A2(_0251_),
    .Y(_0272_),
    .B1(_0249_));
 sg13g2_o21ai_1 _0958_ (.B1(_0257_),
    .Y(_0273_),
    .A1(_0256_),
    .A2(_0271_));
 sg13g2_o21ai_1 _0959_ (.B1(_0273_),
    .Y(_0274_),
    .A1(_0259_),
    .A2(_0271_));
 sg13g2_a21oi_1 _0960_ (.A1(_0267_),
    .A2(_0270_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_o21ai_1 _0961_ (.B1(net191),
    .Y(_0276_),
    .A1(net246),
    .A2(net151));
 sg13g2_nor2_1 _0962_ (.A(_0275_),
    .B(_0276_),
    .Y(_0011_));
 sg13g2_nand3_1 _0963_ (.B(net153),
    .C(_0269_),
    .A(net163),
    .Y(_0277_));
 sg13g2_a21oi_1 _0964_ (.A1(net153),
    .A2(_0269_),
    .Y(_0278_),
    .B1(_0198_));
 sg13g2_a21o_1 _0965_ (.A2(_0269_),
    .A1(net152),
    .B1(_0198_),
    .X(_0279_));
 sg13g2_a21oi_1 _0966_ (.A1(_0277_),
    .A2(_0279_),
    .Y(_0280_),
    .B1(_0224_));
 sg13g2_nand3_1 _0967_ (.B(_0277_),
    .C(_0279_),
    .A(_0224_),
    .Y(_0281_));
 sg13g2_nand2_1 _0968_ (.Y(_0282_),
    .A(net152),
    .B(_0281_));
 sg13g2_nand2b_1 _0969_ (.Y(_0283_),
    .B(_0269_),
    .A_N(net152));
 sg13g2_nor2b_1 _0970_ (.A(_0283_),
    .B_N(net163),
    .Y(_0284_));
 sg13g2_nor3_1 _0971_ (.A(_0198_),
    .B(net152),
    .C(_0269_),
    .Y(_0285_));
 sg13g2_nor3_1 _0972_ (.A(net348),
    .B(_0284_),
    .C(_0285_),
    .Y(_0286_));
 sg13g2_o21ai_1 _0973_ (.B1(_0286_),
    .Y(_0287_),
    .A1(_0280_),
    .A2(_0282_));
 sg13g2_a21oi_1 _0974_ (.A1(net182),
    .A2(_0227_),
    .Y(_0288_),
    .B1(_0244_));
 sg13g2_a21oi_1 _0975_ (.A1(_0287_),
    .A2(_0288_),
    .Y(_0289_),
    .B1(_0257_));
 sg13g2_o21ai_1 _0976_ (.B1(net191),
    .Y(_0290_),
    .A1(net351),
    .A2(net151));
 sg13g2_nor2_1 _0977_ (.A(_0289_),
    .B(_0290_),
    .Y(_0012_));
 sg13g2_o21ai_1 _0978_ (.B1(_0277_),
    .Y(_0291_),
    .A1(_0223_),
    .A2(_0278_));
 sg13g2_xnor2_1 _0979_ (.Y(_0292_),
    .A(_0216_),
    .B(_0232_));
 sg13g2_xnor2_1 _0980_ (.Y(_0293_),
    .A(_0291_),
    .B(_0292_));
 sg13g2_nor3_1 _0981_ (.A(_0215_),
    .B(_0226_),
    .C(_0283_),
    .Y(_0294_));
 sg13g2_nor2_1 _0982_ (.A(_0216_),
    .B(_0268_),
    .Y(_0295_));
 sg13g2_nor2_1 _0983_ (.A(_0204_),
    .B(_0217_),
    .Y(_0296_));
 sg13g2_xnor2_1 _0984_ (.Y(_0297_),
    .A(_0227_),
    .B(_0296_));
 sg13g2_nor3_1 _0985_ (.A(net152),
    .B(_0269_),
    .C(_0297_),
    .Y(_0298_));
 sg13g2_or4_1 _0986_ (.A(net183),
    .B(_0294_),
    .C(_0295_),
    .D(_0298_),
    .X(_0299_));
 sg13g2_a21oi_1 _0987_ (.A1(net152),
    .A2(_0293_),
    .Y(_0300_),
    .B1(_0299_));
 sg13g2_nand2b_1 _0988_ (.Y(_0301_),
    .B(_0262_),
    .A_N(_0300_));
 sg13g2_o21ai_1 _0989_ (.B1(net192),
    .Y(_0302_),
    .A1(net370),
    .A2(net151));
 sg13g2_a21oi_1 _0990_ (.A1(_0273_),
    .A2(_0301_),
    .Y(_0013_),
    .B1(_0302_));
 sg13g2_nor2_1 _0991_ (.A(_0150_),
    .B(_0151_),
    .Y(_0303_));
 sg13g2_nand4_1 _0992_ (.B(\desk_clock.input_debounce.set_hours_reg[1] ),
    .C(\desk_clock.input_debounce.set_hours_reg[0] ),
    .A(\desk_clock.input_debounce.set_hours_reg[2] ),
    .Y(_0304_),
    .D(_0303_));
 sg13g2_nand3_1 _0993_ (.B(\desk_clock.input_debounce.set_minutes_reg[1] ),
    .C(\desk_clock.input_debounce.set_minutes_reg[0] ),
    .A(\desk_clock.input_debounce.set_minutes_reg[2] ),
    .Y(_0305_));
 sg13g2_nor3_2 _0994_ (.A(_0144_),
    .B(_0145_),
    .C(_0305_),
    .Y(_0306_));
 sg13g2_inv_1 _0995_ (.Y(_0307_),
    .A(_0306_));
 sg13g2_nand2_2 _0996_ (.Y(_0308_),
    .A(_0304_),
    .B(_0307_));
 sg13g2_o21ai_1 _0997_ (.B1(net180),
    .Y(_0309_),
    .A1(\desk_clock.clk_seconds[0] ),
    .A2(_0308_));
 sg13g2_nand3_1 _0998_ (.B(_0304_),
    .C(_0307_),
    .A(\desk_clock.display_inst.state[2] ),
    .Y(_0310_));
 sg13g2_nor2_1 _0999_ (.A(_0138_),
    .B(_0139_),
    .Y(_0311_));
 sg13g2_nand4_1 _1000_ (.B(\desk_clock.input_debounce.en_12h_mode_reg[1] ),
    .C(\desk_clock.input_debounce.en_12h_mode_reg[0] ),
    .A(\desk_clock.input_debounce.en_12h_mode_reg[2] ),
    .Y(_0312_),
    .D(_0311_));
 sg13g2_a21oi_1 _1001_ (.A1(\desk_clock.clk_hours[3] ),
    .A2(\desk_clock.clk_hours[2] ),
    .Y(_0313_),
    .B1(\desk_clock.clk_hours[4] ));
 sg13g2_nor3_1 _1002_ (.A(net183),
    .B(_0312_),
    .C(_0313_),
    .Y(_0314_));
 sg13g2_o21ai_1 _1003_ (.B1(_0182_),
    .Y(_0315_),
    .A1(_0184_),
    .A2(_0314_));
 sg13g2_a21oi_1 _1004_ (.A1(_0309_),
    .A2(_0310_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_o21ai_1 _1005_ (.B1(_0243_),
    .Y(_0317_),
    .A1(_0188_),
    .A2(_0316_));
 sg13g2_o21ai_1 _1006_ (.B1(net190),
    .Y(_0318_),
    .A1(net356),
    .A2(net151));
 sg13g2_a21oi_1 _1007_ (.A1(_0273_),
    .A2(_0317_),
    .Y(_0014_),
    .B1(_0318_));
 sg13g2_nor3_1 _1008_ (.A(\desk_clock.display_inst.display_settings.transfer_state[3] ),
    .B(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .C(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .Y(_0319_));
 sg13g2_nor2_1 _1009_ (.A(\desk_clock.display_inst.display_settings.transfer_state[3] ),
    .B(_0237_),
    .Y(_0320_));
 sg13g2_nor2_2 _1010_ (.A(_0319_),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_and2_1 _1011_ (.A(\desk_clock.display_inst.disp_driver.o_serial_load ),
    .B(_0321_),
    .X(_0322_));
 sg13g2_nand2_1 _1012_ (.Y(_0323_),
    .A(\desk_clock.display_inst.disp_driver.o_serial_load ),
    .B(_0321_));
 sg13g2_nor2_2 _1013_ (.A(net164),
    .B(_0321_),
    .Y(_0324_));
 sg13g2_nand2_1 _1014_ (.Y(_0325_),
    .A(net167),
    .B(net154));
 sg13g2_a22oi_1 _1015_ (.Y(_0326_),
    .B1(_0324_),
    .B2(net221),
    .A2(net156),
    .A1(\desk_clock.display_inst.disp_driver.i_data[0] ));
 sg13g2_nor2_1 _1016_ (.A(net186),
    .B(net222),
    .Y(_0015_));
 sg13g2_nand2_1 _1017_ (.Y(_0327_),
    .A(net221),
    .B(net165));
 sg13g2_a21oi_1 _1018_ (.A1(\desk_clock.display_inst.disp_driver.data_reg[1] ),
    .A2(net166),
    .Y(_0328_),
    .B1(net156));
 sg13g2_o21ai_1 _1019_ (.B1(net191),
    .Y(_0329_),
    .A1(net246),
    .A2(net154));
 sg13g2_a21oi_1 _1020_ (.A1(_0327_),
    .A2(_0328_),
    .Y(_0016_),
    .B1(_0329_));
 sg13g2_and2_1 _1021_ (.A(\desk_clock.display_inst.disp_driver.data_reg[1] ),
    .B(net165),
    .X(_0330_));
 sg13g2_a21oi_1 _1022_ (.A1(net234),
    .A2(net166),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_o21ai_1 _1023_ (.B1(net191),
    .Y(_0332_),
    .A1(net351),
    .A2(net154));
 sg13g2_a21oi_1 _1024_ (.A1(net154),
    .A2(_0331_),
    .Y(_0017_),
    .B1(_0332_));
 sg13g2_nand2_1 _1025_ (.Y(_0333_),
    .A(net234),
    .B(net165));
 sg13g2_a21oi_1 _1026_ (.A1(\desk_clock.display_inst.disp_driver.data_reg[3] ),
    .A2(net167),
    .Y(_0334_),
    .B1(net156));
 sg13g2_o21ai_1 _1027_ (.B1(net191),
    .Y(_0335_),
    .A1(\desk_clock.display_inst.disp_driver.i_data[3] ),
    .A2(_0323_));
 sg13g2_a21oi_1 _1028_ (.A1(_0333_),
    .A2(_0334_),
    .Y(_0018_),
    .B1(_0335_));
 sg13g2_a21o_1 _1029_ (.A2(_0322_),
    .A1(\desk_clock.display_inst.disp_driver.i_data[4] ),
    .B1(_0324_),
    .X(_0336_));
 sg13g2_a21oi_1 _1030_ (.A1(net318),
    .A2(net154),
    .Y(_0337_),
    .B1(_0336_));
 sg13g2_o21ai_1 _1031_ (.B1(net190),
    .Y(_0338_),
    .A1(net299),
    .A2(_0325_));
 sg13g2_nor2_1 _1032_ (.A(net319),
    .B(_0338_),
    .Y(_0019_));
 sg13g2_a21oi_1 _1033_ (.A1(net299),
    .A2(net154),
    .Y(_0339_),
    .B1(_0336_));
 sg13g2_o21ai_1 _1034_ (.B1(net190),
    .Y(_0340_),
    .A1(\desk_clock.display_inst.disp_driver.data_reg[5] ),
    .A2(_0325_));
 sg13g2_nor2_1 _1035_ (.A(net300),
    .B(_0340_),
    .Y(_0020_));
 sg13g2_a21oi_1 _1036_ (.A1(net310),
    .A2(net154),
    .Y(_0341_),
    .B1(_0336_));
 sg13g2_o21ai_1 _1037_ (.B1(net190),
    .Y(_0342_),
    .A1(net285),
    .A2(_0325_));
 sg13g2_nor2_1 _1038_ (.A(net311),
    .B(_0342_),
    .Y(_0021_));
 sg13g2_nand2_1 _1039_ (.Y(_0343_),
    .A(net285),
    .B(net164));
 sg13g2_a21oi_1 _1040_ (.A1(net275),
    .A2(net166),
    .Y(_0344_),
    .B1(net156));
 sg13g2_o21ai_1 _1041_ (.B1(net190),
    .Y(_0345_),
    .A1(\desk_clock.display_inst.disp_driver.i_data[7] ),
    .A2(net155));
 sg13g2_a21oi_1 _1042_ (.A1(_0343_),
    .A2(_0344_),
    .Y(_0022_),
    .B1(_0345_));
 sg13g2_nand2_1 _1043_ (.Y(_0346_),
    .A(net275),
    .B(net164));
 sg13g2_a21oi_1 _1044_ (.A1(net238),
    .A2(net166),
    .Y(_0347_),
    .B1(net156));
 sg13g2_o21ai_1 _1045_ (.B1(net189),
    .Y(_0348_),
    .A1(\desk_clock.display_inst.disp_driver.i_addr[0] ),
    .A2(net155));
 sg13g2_a21oi_1 _1046_ (.A1(_0346_),
    .A2(_0347_),
    .Y(_0023_),
    .B1(_0348_));
 sg13g2_nand2_1 _1047_ (.Y(_0349_),
    .A(net238),
    .B(net164));
 sg13g2_a21oi_1 _1048_ (.A1(net211),
    .A2(net166),
    .Y(_0350_),
    .B1(net156));
 sg13g2_o21ai_1 _1049_ (.B1(net189),
    .Y(_0351_),
    .A1(\desk_clock.display_inst.disp_driver.i_addr[1] ),
    .A2(net155));
 sg13g2_a21oi_1 _1050_ (.A1(_0349_),
    .A2(_0350_),
    .Y(_0024_),
    .B1(_0351_));
 sg13g2_nand2_1 _1051_ (.Y(_0352_),
    .A(net211),
    .B(net164));
 sg13g2_a21oi_1 _1052_ (.A1(\desk_clock.display_inst.disp_driver.data_reg[10] ),
    .A2(net166),
    .Y(_0353_),
    .B1(net156));
 sg13g2_o21ai_1 _1053_ (.B1(net189),
    .Y(_0354_),
    .A1(\desk_clock.display_inst.disp_driver.i_addr[2] ),
    .A2(net155));
 sg13g2_a21oi_1 _1054_ (.A1(_0352_),
    .A2(_0353_),
    .Y(_0025_),
    .B1(_0354_));
 sg13g2_a22oi_1 _1055_ (.Y(_0355_),
    .B1(_0324_),
    .B2(\desk_clock.display_inst.disp_driver.data_reg[11] ),
    .A2(net156),
    .A1(\desk_clock.display_inst.disp_driver.i_addr[3] ));
 sg13g2_nand2_1 _1056_ (.Y(_0356_),
    .A(net191),
    .B(net154));
 sg13g2_nand4_1 _1057_ (.B(net189),
    .C(net164),
    .A(net230),
    .Y(_0357_),
    .D(net155));
 sg13g2_o21ai_1 _1058_ (.B1(_0357_),
    .Y(_0026_),
    .A1(net186),
    .A2(_0355_));
 sg13g2_nand2_1 _1059_ (.Y(_0358_),
    .A(net206),
    .B(net164));
 sg13g2_nor2b_1 _1060_ (.A(net206),
    .B_N(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .Y(_0359_));
 sg13g2_a21oi_1 _1061_ (.A1(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .A2(_0178_),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_nand2_1 _1062_ (.Y(_0361_),
    .A(net190),
    .B(_0360_));
 sg13g2_a21oi_1 _1063_ (.A1(net155),
    .A2(_0358_),
    .Y(_0027_),
    .B1(_0361_));
 sg13g2_nor2_1 _1064_ (.A(\desk_clock.display_inst.state[3] ),
    .B(_0188_),
    .Y(_0362_));
 sg13g2_nor2b_2 _1065_ (.A(_0362_),
    .B_N(\desk_clock.display_control_inst.display_update ),
    .Y(_0363_));
 sg13g2_o21ai_1 _1066_ (.B1(\desk_clock.display_control_inst.display_update ),
    .Y(_0364_),
    .A1(\desk_clock.display_inst.state[3] ),
    .A2(_0188_));
 sg13g2_o21ai_1 _1067_ (.B1(net188),
    .Y(_0365_),
    .A1(\desk_clock.clk_hours[0] ),
    .A2(net159));
 sg13g2_a21oi_1 _1068_ (.A1(_0176_),
    .A2(net159),
    .Y(_0028_),
    .B1(_0365_));
 sg13g2_o21ai_1 _1069_ (.B1(net188),
    .Y(_0366_),
    .A1(\desk_clock.clk_hours[1] ),
    .A2(net159));
 sg13g2_a21oi_1 _1070_ (.A1(_0175_),
    .A2(net162),
    .Y(_0029_),
    .B1(_0366_));
 sg13g2_o21ai_1 _1071_ (.B1(\desk_clock.clk_hours[2] ),
    .Y(_0367_),
    .A1(net178),
    .A2(_0160_));
 sg13g2_a21oi_1 _1072_ (.A1(_0160_),
    .A2(_0005_),
    .Y(_0368_),
    .B1(\desk_clock.clk_hours[2] ));
 sg13g2_nor3_1 _1073_ (.A(\desk_clock.clk_hours[1] ),
    .B(\desk_clock.clk_hours[0] ),
    .C(_0368_),
    .Y(_0369_));
 sg13g2_a21oi_1 _1074_ (.A1(_0367_),
    .A2(_0369_),
    .Y(_0370_),
    .B1(_0312_));
 sg13g2_a21oi_1 _1075_ (.A1(net178),
    .A2(\desk_clock.clk_hours[3] ),
    .Y(_0371_),
    .B1(_0313_));
 sg13g2_xor2_1 _1076_ (.B(_0371_),
    .A(_0006_),
    .X(_0372_));
 sg13g2_a221oi_1 _1077_ (.B2(_0372_),
    .C1(net159),
    .B1(_0370_),
    .A1(_0161_),
    .Y(_0373_),
    .A2(_0312_));
 sg13g2_a21oi_1 _1078_ (.A1(net339),
    .A2(net159),
    .Y(_0374_),
    .B1(_0373_));
 sg13g2_nor2_1 _1079_ (.A(net184),
    .B(net340),
    .Y(_0030_));
 sg13g2_nand3b_1 _1080_ (.B(\desk_clock.clk_hours[3] ),
    .C(_0161_),
    .Y(_0375_),
    .A_N(net178));
 sg13g2_nand3_1 _1081_ (.B(_0160_),
    .C(\desk_clock.clk_hours[2] ),
    .A(net178),
    .Y(_0376_));
 sg13g2_nand3_1 _1082_ (.B(_0375_),
    .C(_0376_),
    .A(_0370_),
    .Y(_0377_));
 sg13g2_a21oi_1 _1083_ (.A1(_0160_),
    .A2(_0312_),
    .Y(_0378_),
    .B1(net160));
 sg13g2_a22oi_1 _1084_ (.Y(_0379_),
    .B1(_0377_),
    .B2(_0378_),
    .A2(net160),
    .A1(net314));
 sg13g2_nor2_1 _1085_ (.A(net184),
    .B(net315),
    .Y(_0031_));
 sg13g2_a21oi_1 _1086_ (.A1(net178),
    .A2(_0312_),
    .Y(_0380_),
    .B1(net159));
 sg13g2_o21ai_1 _1087_ (.B1(net188),
    .Y(_0381_),
    .A1(net336),
    .A2(_0363_));
 sg13g2_nor2_1 _1088_ (.A(_0380_),
    .B(net337),
    .Y(_0032_));
 sg13g2_o21ai_1 _1089_ (.B1(net188),
    .Y(_0382_),
    .A1(\desk_clock.clk_minutes[0] ),
    .A2(net158));
 sg13g2_a21oi_1 _1090_ (.A1(_0174_),
    .A2(net158),
    .Y(_0033_),
    .B1(_0382_));
 sg13g2_o21ai_1 _1091_ (.B1(net187),
    .Y(_0383_),
    .A1(\desk_clock.clk_minutes[1] ),
    .A2(net158));
 sg13g2_a21oi_1 _1092_ (.A1(_0173_),
    .A2(net158),
    .Y(_0034_),
    .B1(_0383_));
 sg13g2_o21ai_1 _1093_ (.B1(net188),
    .Y(_0384_),
    .A1(net343),
    .A2(_0363_));
 sg13g2_a21oi_1 _1094_ (.A1(_0164_),
    .A2(_0363_),
    .Y(_0035_),
    .B1(net344));
 sg13g2_o21ai_1 _1095_ (.B1(net187),
    .Y(_0385_),
    .A1(net353),
    .A2(net157));
 sg13g2_a21oi_1 _1096_ (.A1(_0163_),
    .A2(net157),
    .Y(_0036_),
    .B1(_0385_));
 sg13g2_o21ai_1 _1097_ (.B1(net187),
    .Y(_0386_),
    .A1(\desk_clock.clk_minutes[4] ),
    .A2(net158));
 sg13g2_a21oi_1 _1098_ (.A1(_0172_),
    .A2(net158),
    .Y(_0037_),
    .B1(_0386_));
 sg13g2_o21ai_1 _1099_ (.B1(net187),
    .Y(_0387_),
    .A1(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ),
    .A2(net157));
 sg13g2_a21oi_1 _1100_ (.A1(_0162_),
    .A2(net157),
    .Y(_0038_),
    .B1(_0387_));
 sg13g2_o21ai_1 _1101_ (.B1(net193),
    .Y(_0388_),
    .A1(\desk_clock.clk_seconds[0] ),
    .A2(net161));
 sg13g2_a21oi_1 _1102_ (.A1(_0171_),
    .A2(net159),
    .Y(_0039_),
    .B1(_0388_));
 sg13g2_o21ai_1 _1103_ (.B1(net193),
    .Y(_0389_),
    .A1(\desk_clock.clk_seconds[1] ),
    .A2(net161));
 sg13g2_a21oi_1 _1104_ (.A1(_0170_),
    .A2(net159),
    .Y(_0040_),
    .B1(_0389_));
 sg13g2_o21ai_1 _1105_ (.B1(net193),
    .Y(_0390_),
    .A1(\desk_clock.clk_seconds[2] ),
    .A2(net160));
 sg13g2_a21oi_1 _1106_ (.A1(_0169_),
    .A2(net160),
    .Y(_0041_),
    .B1(_0390_));
 sg13g2_o21ai_1 _1107_ (.B1(net193),
    .Y(_0391_),
    .A1(\desk_clock.clk_seconds[3] ),
    .A2(net161));
 sg13g2_a21oi_1 _1108_ (.A1(_0168_),
    .A2(net160),
    .Y(_0042_),
    .B1(_0391_));
 sg13g2_o21ai_1 _1109_ (.B1(net193),
    .Y(_0392_),
    .A1(\desk_clock.clk_seconds[4] ),
    .A2(net161));
 sg13g2_a21oi_1 _1110_ (.A1(_0167_),
    .A2(net160),
    .Y(_0043_),
    .B1(_0392_));
 sg13g2_o21ai_1 _1111_ (.B1(net193),
    .Y(_0393_),
    .A1(\desk_clock.clk_seconds[5] ),
    .A2(net160));
 sg13g2_a21oi_1 _1112_ (.A1(_0166_),
    .A2(net160),
    .Y(_0044_),
    .B1(_0393_));
 sg13g2_nor3_2 _1113_ (.A(\desk_clock.display_inst.display_settings.transfer_state[3] ),
    .B(_0237_),
    .C(_0240_),
    .Y(_0394_));
 sg13g2_mux2_1 _1114_ (.A0(net182),
    .A1(_0003_),
    .S(_0394_),
    .X(_0395_));
 sg13g2_nor2_1 _1115_ (.A(net157),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_nand3b_1 _1116_ (.B(net187),
    .C(_0186_),
    .Y(_0397_),
    .A_N(net382));
 sg13g2_nor2_1 _1117_ (.A(net324),
    .B(net162),
    .Y(_0398_));
 sg13g2_nor3_1 _1118_ (.A(_0396_),
    .B(_0397_),
    .C(_0398_),
    .Y(_0045_));
 sg13g2_nor2_1 _1119_ (.A(net157),
    .B(_0394_),
    .Y(_0399_));
 sg13g2_nand3b_1 _1120_ (.B(net158),
    .C(_0394_),
    .Y(_0400_),
    .A_N(_0192_));
 sg13g2_a22oi_1 _1121_ (.Y(_0401_),
    .B1(_0399_),
    .B2(net180),
    .A2(net157),
    .A1(net364));
 sg13g2_a21oi_1 _1122_ (.A1(_0400_),
    .A2(_0401_),
    .Y(_0046_),
    .B1(_0397_));
 sg13g2_nand3b_1 _1123_ (.B(net158),
    .C(_0394_),
    .Y(_0402_),
    .A_N(_0196_));
 sg13g2_a22oi_1 _1124_ (.Y(_0403_),
    .B1(_0399_),
    .B2(net179),
    .A2(net157),
    .A1(net364));
 sg13g2_a21oi_1 _1125_ (.A1(_0402_),
    .A2(_0403_),
    .Y(_0047_),
    .B1(_0397_));
 sg13g2_nor2b_1 _1126_ (.A(_0178_),
    .B_N(_0359_),
    .Y(_0404_));
 sg13g2_o21ai_1 _1127_ (.B1(_0246_),
    .Y(_0405_),
    .A1(_0319_),
    .A2(_0404_));
 sg13g2_nand2b_2 _1128_ (.Y(_0406_),
    .B(_0405_),
    .A_N(_0242_));
 sg13g2_nor2_1 _1129_ (.A(net371),
    .B(_0242_),
    .Y(_0407_));
 sg13g2_o21ai_1 _1130_ (.B1(_0406_),
    .Y(_0408_),
    .A1(_0243_),
    .A2(_0407_));
 sg13g2_nand2_2 _1131_ (.Y(_0409_),
    .A(net187),
    .B(_0238_));
 sg13g2_o21ai_1 _1132_ (.B1(_0408_),
    .Y(_0410_),
    .A1(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .A2(_0406_));
 sg13g2_nor2_1 _1133_ (.A(_0409_),
    .B(net372),
    .Y(_0049_));
 sg13g2_nand2_1 _1134_ (.Y(_0411_),
    .A(_0236_),
    .B(_0406_));
 sg13g2_nand2b_1 _1135_ (.Y(_0412_),
    .B(_0411_),
    .A_N(_0234_));
 sg13g2_a21oi_1 _1136_ (.A1(_0254_),
    .A2(_0412_),
    .Y(_0413_),
    .B1(_0409_));
 sg13g2_o21ai_1 _1137_ (.B1(_0413_),
    .Y(_0414_),
    .A1(net390),
    .A2(_0406_));
 sg13g2_inv_1 _1138_ (.Y(_0050_),
    .A(_0414_));
 sg13g2_nor3_1 _1139_ (.A(\desk_clock.display_inst.display_settings.transfer_state[3] ),
    .B(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .C(_0236_),
    .Y(_0415_));
 sg13g2_nand3_1 _1140_ (.B(_0406_),
    .C(_0415_),
    .A(_0254_),
    .Y(_0416_));
 sg13g2_o21ai_1 _1141_ (.B1(_0416_),
    .Y(_0417_),
    .A1(net391),
    .A2(_0406_));
 sg13g2_nor2_1 _1142_ (.A(_0409_),
    .B(_0417_),
    .Y(_0051_));
 sg13g2_nor3_1 _1143_ (.A(net204),
    .B(_0409_),
    .C(_0411_),
    .Y(_0052_));
 sg13g2_nor3_1 _1144_ (.A(_0247_),
    .B(_0252_),
    .C(_0272_),
    .Y(_0418_));
 sg13g2_o21ai_1 _1145_ (.B1(net189),
    .Y(_0419_),
    .A1(net369),
    .A2(_0253_));
 sg13g2_nor3_1 _1146_ (.A(_0243_),
    .B(_0418_),
    .C(_0419_),
    .Y(_0053_));
 sg13g2_nor3_1 _1147_ (.A(\desk_clock.display_inst.display_settings.transfer_state[0] ),
    .B(_0243_),
    .C(_0272_),
    .Y(_0420_));
 sg13g2_o21ai_1 _1148_ (.B1(net150),
    .Y(_0421_),
    .A1(_0262_),
    .A2(_0420_));
 sg13g2_o21ai_1 _1149_ (.B1(net189),
    .Y(_0422_),
    .A1(net357),
    .A2(net150));
 sg13g2_nor2b_1 _1150_ (.A(_0422_),
    .B_N(_0421_),
    .Y(_0054_));
 sg13g2_nor3_1 _1151_ (.A(_0234_),
    .B(_0243_),
    .C(_0272_),
    .Y(_0423_));
 sg13g2_a21oi_1 _1152_ (.A1(net180),
    .A2(_0243_),
    .Y(_0424_),
    .B1(_0423_));
 sg13g2_o21ai_1 _1153_ (.B1(net189),
    .Y(_0425_),
    .A1(net349),
    .A2(net150));
 sg13g2_a21oi_1 _1154_ (.A1(net150),
    .A2(_0424_),
    .Y(_0055_),
    .B1(_0425_));
 sg13g2_o21ai_1 _1155_ (.B1(net150),
    .Y(_0426_),
    .A1(_0165_),
    .A2(_0244_));
 sg13g2_a21oi_1 _1156_ (.A1(_0244_),
    .A2(_0249_),
    .Y(_0427_),
    .B1(_0426_));
 sg13g2_o21ai_1 _1157_ (.B1(net189),
    .Y(_0428_),
    .A1(net342),
    .A2(net150));
 sg13g2_nor2_1 _1158_ (.A(_0427_),
    .B(_0428_),
    .Y(_0056_));
 sg13g2_nor2_1 _1159_ (.A(_0183_),
    .B(_0244_),
    .Y(_0429_));
 sg13g2_o21ai_1 _1160_ (.B1(net190),
    .Y(_0430_),
    .A1(net341),
    .A2(net150));
 sg13g2_a21oi_1 _1161_ (.A1(net150),
    .A2(_0429_),
    .Y(_0057_),
    .B1(_0430_));
 sg13g2_nor2_1 _1162_ (.A(_0156_),
    .B(_0157_),
    .Y(_0431_));
 sg13g2_nand4_1 _1163_ (.B(\desk_clock.input_debounce.fast_set_reg[1] ),
    .C(\desk_clock.input_debounce.fast_set_reg[0] ),
    .A(\desk_clock.input_debounce.fast_set_reg[2] ),
    .Y(_0432_),
    .D(_0431_));
 sg13g2_nor2b_1 _1164_ (.A(\desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold ),
    .B_N(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .Y(_0433_));
 sg13g2_o21ai_1 _1165_ (.B1(_0432_),
    .Y(_0434_),
    .A1(_0131_),
    .A2(\desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold ));
 sg13g2_o21ai_1 _1166_ (.B1(_0434_),
    .Y(_0435_),
    .A1(_0432_),
    .A2(_0433_));
 sg13g2_nor3_1 _1167_ (.A(\desk_clock.display_control_inst.o_write_config ),
    .B(\desk_clock.display_inst.state[3] ),
    .C(_0186_),
    .Y(_0436_));
 sg13g2_nor2_2 _1168_ (.A(_0130_),
    .B(\desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold ),
    .Y(_0437_));
 sg13g2_a22oi_1 _1169_ (.Y(_0438_),
    .B1(_0436_),
    .B2(net395),
    .A2(_0435_),
    .A1(_0308_));
 sg13g2_o21ai_1 _1170_ (.B1(net396),
    .Y(_0439_),
    .A1(_0308_),
    .A2(_0437_));
 sg13g2_nand2b_1 _1171_ (.Y(_0440_),
    .B(_0241_),
    .A_N(net324));
 sg13g2_nand3_1 _1172_ (.B(net397),
    .C(_0440_),
    .A(net188),
    .Y(_0058_));
 sg13g2_nand2b_2 _1173_ (.Y(_0441_),
    .B(net155),
    .A_N(_0361_));
 sg13g2_xnor2_1 _1174_ (.Y(_0442_),
    .A(net361),
    .B(\desk_clock.display_inst.disp_driver.transfer_state[0] ));
 sg13g2_nor2_1 _1175_ (.A(_0441_),
    .B(net362),
    .Y(_0059_));
 sg13g2_and3_1 _1176_ (.X(_0443_),
    .A(net262),
    .B(\desk_clock.display_inst.disp_driver.transfer_state[1] ),
    .C(\desk_clock.display_inst.disp_driver.transfer_state[0] ));
 sg13g2_a21oi_1 _1177_ (.A1(\desk_clock.display_inst.disp_driver.transfer_state[1] ),
    .A2(\desk_clock.display_inst.disp_driver.transfer_state[0] ),
    .Y(_0444_),
    .B1(net262));
 sg13g2_nor3_1 _1178_ (.A(_0441_),
    .B(_0443_),
    .C(net263),
    .Y(_0060_));
 sg13g2_nand2_1 _1179_ (.Y(_0445_),
    .A(net332),
    .B(_0443_));
 sg13g2_xnor2_1 _1180_ (.Y(_0446_),
    .A(net332),
    .B(_0443_));
 sg13g2_nor2_1 _1181_ (.A(_0441_),
    .B(net333),
    .Y(_0061_));
 sg13g2_xor2_1 _1182_ (.B(_0445_),
    .A(net387),
    .X(_0447_));
 sg13g2_nor2_1 _1183_ (.A(_0441_),
    .B(_0447_),
    .Y(_0062_));
 sg13g2_nand2_1 _1184_ (.Y(_0448_),
    .A(net255),
    .B(net164));
 sg13g2_nand2_1 _1185_ (.Y(_0449_),
    .A(net240),
    .B(net167));
 sg13g2_a21oi_1 _1186_ (.A1(_0448_),
    .A2(_0449_),
    .Y(_0063_),
    .B1(_0356_));
 sg13g2_nand2_1 _1187_ (.Y(_0450_),
    .A(net240),
    .B(net165));
 sg13g2_nand2_1 _1188_ (.Y(_0451_),
    .A(net236),
    .B(net167));
 sg13g2_a21oi_1 _1189_ (.A1(_0450_),
    .A2(_0451_),
    .Y(_0064_),
    .B1(_0356_));
 sg13g2_nand2_1 _1190_ (.Y(_0452_),
    .A(net236),
    .B(net165));
 sg13g2_nand2_1 _1191_ (.Y(_0453_),
    .A(\desk_clock.display_inst.disp_driver.data_reg[14] ),
    .B(net166));
 sg13g2_a21oi_1 _1192_ (.A1(_0452_),
    .A2(_0453_),
    .Y(_0065_),
    .B1(_0356_));
 sg13g2_nand2_1 _1193_ (.Y(_0454_),
    .A(\desk_clock.display_inst.disp_driver.data_reg[14] ),
    .B(net165));
 sg13g2_nand2_1 _1194_ (.Y(_0455_),
    .A(net248),
    .B(net166));
 sg13g2_a21oi_1 _1195_ (.A1(_0454_),
    .A2(_0455_),
    .Y(_0066_),
    .B1(_0356_));
 sg13g2_a21o_1 _1196_ (.A2(_0440_),
    .A1(net364),
    .B1(net186),
    .X(_0067_));
 sg13g2_nor2_1 _1197_ (.A(_0131_),
    .B(net185),
    .Y(_0068_));
 sg13g2_nand4_1 _1198_ (.B(\desk_clock.clk_seconds[4] ),
    .C(\desk_clock.clk_seconds[3] ),
    .A(\desk_clock.clk_seconds[5] ),
    .Y(_0456_),
    .D(\desk_clock.clk_seconds[2] ));
 sg13g2_and2_1 _1199_ (.A(net193),
    .B(_0456_),
    .X(_0457_));
 sg13g2_o21ai_1 _1200_ (.B1(_0457_),
    .Y(_0458_),
    .A1(_0304_),
    .A2(_0307_));
 sg13g2_xnor2_1 _1201_ (.Y(_0459_),
    .A(net385),
    .B(_0437_));
 sg13g2_nor2_1 _1202_ (.A(_0458_),
    .B(net386),
    .Y(_0069_));
 sg13g2_and3_1 _1203_ (.X(_0460_),
    .A(net295),
    .B(\desk_clock.clk_seconds[0] ),
    .C(_0437_));
 sg13g2_a21oi_1 _1204_ (.A1(\desk_clock.clk_seconds[0] ),
    .A2(_0437_),
    .Y(_0461_),
    .B1(net295));
 sg13g2_nor3_1 _1205_ (.A(_0458_),
    .B(_0460_),
    .C(net296),
    .Y(_0070_));
 sg13g2_nor2_1 _1206_ (.A(net377),
    .B(_0460_),
    .Y(_0462_));
 sg13g2_and2_1 _1207_ (.A(net377),
    .B(_0460_),
    .X(_0463_));
 sg13g2_and4_1 _1208_ (.A(net322),
    .B(net368),
    .C(net365),
    .D(_0437_),
    .X(_0464_));
 sg13g2_nor4_1 _1209_ (.A(_0458_),
    .B(net378),
    .C(_0463_),
    .D(_0464_),
    .Y(_0071_));
 sg13g2_a21oi_1 _1210_ (.A1(\desk_clock.clk_seconds[1] ),
    .A2(\desk_clock.clk_seconds[0] ),
    .Y(_0465_),
    .B1(\desk_clock.clk_seconds[2] ));
 sg13g2_nor2b_1 _1211_ (.A(_0465_),
    .B_N(_0464_),
    .Y(_0466_));
 sg13g2_or2_1 _1212_ (.X(_0467_),
    .B(_0466_),
    .A(_0458_));
 sg13g2_and2_1 _1213_ (.A(net365),
    .B(_0463_),
    .X(_0468_));
 sg13g2_nor2_1 _1214_ (.A(net365),
    .B(_0463_),
    .Y(_0469_));
 sg13g2_nor3_1 _1215_ (.A(_0467_),
    .B(_0468_),
    .C(net366),
    .Y(_0072_));
 sg13g2_nor2_1 _1216_ (.A(net368),
    .B(_0468_),
    .Y(_0470_));
 sg13g2_and2_1 _1217_ (.A(net368),
    .B(_0468_),
    .X(_0471_));
 sg13g2_nor3_1 _1218_ (.A(_0467_),
    .B(_0470_),
    .C(_0471_),
    .Y(_0073_));
 sg13g2_nor2_1 _1219_ (.A(net322),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_nor2_1 _1220_ (.A(_0467_),
    .B(net323),
    .Y(_0074_));
 sg13g2_nor2b_1 _1221_ (.A(_0308_),
    .B_N(_0466_),
    .Y(_0473_));
 sg13g2_inv_1 _1222_ (.Y(_0474_),
    .A(_0473_));
 sg13g2_nand2_1 _1223_ (.Y(_0475_),
    .A(_0304_),
    .B(_0306_));
 sg13g2_o21ai_1 _1224_ (.B1(_0474_),
    .Y(_0476_),
    .A1(_0435_),
    .A2(_0475_));
 sg13g2_nor2_1 _1225_ (.A(net367),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nand3_1 _1226_ (.B(\desk_clock.clk_minutes[4] ),
    .C(\desk_clock.clk_minutes[3] ),
    .A(\desk_clock.clk_minutes[5] ),
    .Y(_0478_));
 sg13g2_o21ai_1 _1227_ (.B1(net187),
    .Y(_0479_),
    .A1(_0164_),
    .A2(_0478_));
 sg13g2_and2_1 _1228_ (.A(net367),
    .B(_0476_),
    .X(_0480_));
 sg13g2_nor3_1 _1229_ (.A(_0477_),
    .B(_0479_),
    .C(_0480_),
    .Y(_0075_));
 sg13g2_xnor2_1 _1230_ (.Y(_0481_),
    .A(net374),
    .B(_0480_));
 sg13g2_nor2_1 _1231_ (.A(_0479_),
    .B(_0481_),
    .Y(_0076_));
 sg13g2_nand2b_1 _1232_ (.Y(_0482_),
    .B(_0475_),
    .A_N(_0466_));
 sg13g2_a21oi_1 _1233_ (.A1(\desk_clock.clk_minutes[1] ),
    .A2(\desk_clock.clk_minutes[0] ),
    .Y(_0483_),
    .B1(\desk_clock.clk_minutes[2] ));
 sg13g2_nor2_1 _1234_ (.A(_0478_),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_nand2_1 _1235_ (.Y(_0485_),
    .A(_0482_),
    .B(_0484_));
 sg13g2_nand3_1 _1236_ (.B(net374),
    .C(net367),
    .A(net287),
    .Y(_0486_));
 sg13g2_nand2_1 _1237_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_a21o_1 _1238_ (.A2(_0487_),
    .A1(_0476_),
    .B1(_0479_),
    .X(_0488_));
 sg13g2_a21oi_1 _1239_ (.A1(\desk_clock.clk_minutes[1] ),
    .A2(_0480_),
    .Y(_0489_),
    .B1(net287));
 sg13g2_nor2_1 _1240_ (.A(_0488_),
    .B(net288),
    .Y(_0077_));
 sg13g2_nand2_1 _1241_ (.Y(_0490_),
    .A(_0476_),
    .B(_0485_));
 sg13g2_or2_1 _1242_ (.X(_0491_),
    .B(_0490_),
    .A(_0486_));
 sg13g2_nand2_1 _1243_ (.Y(_0492_),
    .A(_0163_),
    .B(net187));
 sg13g2_a22oi_1 _1244_ (.Y(_0078_),
    .B1(_0492_),
    .B2(_0488_),
    .A2(_0491_),
    .A1(_0163_));
 sg13g2_nor2_1 _1245_ (.A(_0163_),
    .B(_0486_),
    .Y(_0493_));
 sg13g2_nand2_1 _1246_ (.Y(_0494_),
    .A(net305),
    .B(_0493_));
 sg13g2_nand2_1 _1247_ (.Y(_0495_),
    .A(_0485_),
    .B(_0494_));
 sg13g2_a21o_1 _1248_ (.A2(_0495_),
    .A1(_0476_),
    .B1(_0479_),
    .X(_0496_));
 sg13g2_a21oi_1 _1249_ (.A1(_0476_),
    .A2(_0493_),
    .Y(_0497_),
    .B1(net305));
 sg13g2_nor2_1 _1250_ (.A(_0496_),
    .B(net306),
    .Y(_0079_));
 sg13g2_o21ai_1 _1251_ (.B1(_0162_),
    .Y(_0498_),
    .A1(_0490_),
    .A2(_0494_));
 sg13g2_o21ai_1 _1252_ (.B1(_0496_),
    .Y(_0499_),
    .A1(net346),
    .A2(net186));
 sg13g2_and2_1 _1253_ (.A(_0498_),
    .B(_0499_),
    .X(_0080_));
 sg13g2_nor3_1 _1254_ (.A(_0304_),
    .B(_0306_),
    .C(_0435_),
    .Y(_0500_));
 sg13g2_a21o_2 _1255_ (.A2(_0484_),
    .A1(_0473_),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_nand2_1 _1256_ (.Y(_0502_),
    .A(\desk_clock.clk_hours[0] ),
    .B(_0501_));
 sg13g2_a21o_2 _1257_ (.A2(net403),
    .A1(net178),
    .B1(net184),
    .X(_0503_));
 sg13g2_xnor2_1 _1258_ (.Y(_0504_),
    .A(net383),
    .B(_0501_));
 sg13g2_nor2_1 _1259_ (.A(_0503_),
    .B(_0504_),
    .Y(_0081_));
 sg13g2_nand2_1 _1260_ (.Y(_0505_),
    .A(net379),
    .B(\desk_clock.clk_hours[0] ));
 sg13g2_xor2_1 _1261_ (.B(_0502_),
    .A(net379),
    .X(_0506_));
 sg13g2_nor2_1 _1262_ (.A(_0503_),
    .B(net380),
    .Y(_0082_));
 sg13g2_nor2_1 _1263_ (.A(_0161_),
    .B(_0505_),
    .Y(_0507_));
 sg13g2_o21ai_1 _1264_ (.B1(net178),
    .Y(_0508_),
    .A1(\desk_clock.clk_hours[3] ),
    .A2(_0507_));
 sg13g2_xor2_1 _1265_ (.B(_0505_),
    .A(net398),
    .X(_0509_));
 sg13g2_nand2_1 _1266_ (.Y(_0510_),
    .A(_0508_),
    .B(_0509_));
 sg13g2_mux2_1 _1267_ (.A0(_0161_),
    .A1(_0510_),
    .S(_0501_),
    .X(_0511_));
 sg13g2_nor2_1 _1268_ (.A(_0503_),
    .B(net399),
    .Y(_0083_));
 sg13g2_nand2_1 _1269_ (.Y(_0512_),
    .A(\desk_clock.clk_hours[3] ),
    .B(_0507_));
 sg13g2_nand2_1 _1270_ (.Y(_0513_),
    .A(_0508_),
    .B(_0512_));
 sg13g2_nand2_1 _1271_ (.Y(_0514_),
    .A(_0501_),
    .B(_0507_));
 sg13g2_a221oi_1 _1272_ (.B2(_0160_),
    .C1(_0503_),
    .B1(_0514_),
    .A1(_0501_),
    .Y(_0084_),
    .A2(_0513_));
 sg13g2_o21ai_1 _1273_ (.B1(_0508_),
    .Y(_0515_),
    .A1(_0005_),
    .A2(_0512_));
 sg13g2_a21oi_1 _1274_ (.A1(net401),
    .A2(_0512_),
    .Y(_0516_),
    .B1(_0515_));
 sg13g2_mux2_1 _1275_ (.A0(net178),
    .A1(_0516_),
    .S(_0501_),
    .X(_0517_));
 sg13g2_nor2b_1 _1276_ (.A(_0503_),
    .B_N(_0517_),
    .Y(_0085_));
 sg13g2_nor2b_1 _1277_ (.A(\desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold ),
    .B_N(\desk_clock.clk_gen_inst.refclk_div[3] ),
    .Y(_0518_));
 sg13g2_o21ai_1 _1278_ (.B1(net198),
    .Y(_0519_),
    .A1(\desk_clock.input_debounce.fast_set_reg[0] ),
    .A2(net175));
 sg13g2_a21oi_1 _1279_ (.A1(_0159_),
    .A2(net175),
    .Y(_0086_),
    .B1(_0519_));
 sg13g2_o21ai_1 _1280_ (.B1(net198),
    .Y(_0520_),
    .A1(\desk_clock.input_debounce.fast_set_reg[1] ),
    .A2(net172));
 sg13g2_a21oi_1 _1281_ (.A1(_0158_),
    .A2(net172),
    .Y(_0087_),
    .B1(_0520_));
 sg13g2_o21ai_1 _1282_ (.B1(net198),
    .Y(_0521_),
    .A1(net209),
    .A2(net172));
 sg13g2_a21oi_1 _1283_ (.A1(_0157_),
    .A2(net172),
    .Y(_0088_),
    .B1(_0521_));
 sg13g2_o21ai_1 _1284_ (.B1(net198),
    .Y(_0522_),
    .A1(net298),
    .A2(net172));
 sg13g2_a21oi_1 _1285_ (.A1(_0156_),
    .A2(net172),
    .Y(_0089_),
    .B1(_0522_));
 sg13g2_o21ai_1 _1286_ (.B1(net197),
    .Y(_0523_),
    .A1(\desk_clock.input_debounce.fast_set_reg[4] ),
    .A2(net174));
 sg13g2_a21oi_1 _1287_ (.A1(_0154_),
    .A2(net174),
    .Y(_0090_),
    .B1(_0523_));
 sg13g2_o21ai_1 _1288_ (.B1(net197),
    .Y(_0524_),
    .A1(net213),
    .A2(net174));
 sg13g2_a21oi_1 _1289_ (.A1(_0155_),
    .A2(net174),
    .Y(_0091_),
    .B1(_0524_));
 sg13g2_o21ai_1 _1290_ (.B1(net196),
    .Y(_0525_),
    .A1(\desk_clock.input_debounce.set_hours_reg[0] ),
    .A2(net170));
 sg13g2_a21oi_1 _1291_ (.A1(_0153_),
    .A2(net170),
    .Y(_0092_),
    .B1(_0525_));
 sg13g2_o21ai_1 _1292_ (.B1(net196),
    .Y(_0526_),
    .A1(\desk_clock.input_debounce.set_hours_reg[1] ),
    .A2(net170));
 sg13g2_a21oi_1 _1293_ (.A1(_0152_),
    .A2(net170),
    .Y(_0093_),
    .B1(_0526_));
 sg13g2_o21ai_1 _1294_ (.B1(net196),
    .Y(_0527_),
    .A1(net289),
    .A2(net171));
 sg13g2_a21oi_1 _1295_ (.A1(_0151_),
    .A2(net170),
    .Y(_0094_),
    .B1(_0527_));
 sg13g2_o21ai_1 _1296_ (.B1(net195),
    .Y(_0528_),
    .A1(\desk_clock.input_debounce.set_hours_reg[3] ),
    .A2(net170));
 sg13g2_a21oi_1 _1297_ (.A1(_0150_),
    .A2(net170),
    .Y(_0095_),
    .B1(_0528_));
 sg13g2_o21ai_1 _1298_ (.B1(net196),
    .Y(_0529_),
    .A1(net253),
    .A2(net171));
 sg13g2_a21oi_1 _1299_ (.A1(_0148_),
    .A2(net173),
    .Y(_0096_),
    .B1(_0529_));
 sg13g2_o21ai_1 _1300_ (.B1(net197),
    .Y(_0530_),
    .A1(net267),
    .A2(net173));
 sg13g2_a21oi_1 _1301_ (.A1(_0149_),
    .A2(net173),
    .Y(_0097_),
    .B1(_0530_));
 sg13g2_o21ai_1 _1302_ (.B1(net195),
    .Y(_0531_),
    .A1(\desk_clock.input_debounce.set_minutes_reg[0] ),
    .A2(net168));
 sg13g2_a21oi_1 _1303_ (.A1(_0147_),
    .A2(net168),
    .Y(_0098_),
    .B1(_0531_));
 sg13g2_o21ai_1 _1304_ (.B1(net195),
    .Y(_0532_),
    .A1(net256),
    .A2(net168));
 sg13g2_a21oi_1 _1305_ (.A1(_0146_),
    .A2(net168),
    .Y(_0099_),
    .B1(_0532_));
 sg13g2_o21ai_1 _1306_ (.B1(net195),
    .Y(_0533_),
    .A1(net293),
    .A2(net168));
 sg13g2_a21oi_1 _1307_ (.A1(_0145_),
    .A2(net168),
    .Y(_0100_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1308_ (.B1(net195),
    .Y(_0534_),
    .A1(net309),
    .A2(net168));
 sg13g2_a21oi_1 _1309_ (.A1(_0144_),
    .A2(net168),
    .Y(_0101_),
    .B1(_0534_));
 sg13g2_o21ai_1 _1310_ (.B1(net196),
    .Y(_0535_),
    .A1(\desk_clock.input_debounce.set_minutes_reg[4] ),
    .A2(net170));
 sg13g2_a21oi_1 _1311_ (.A1(_0142_),
    .A2(net171),
    .Y(_0102_),
    .B1(_0535_));
 sg13g2_o21ai_1 _1312_ (.B1(net196),
    .Y(_0536_),
    .A1(net223),
    .A2(net171));
 sg13g2_a21oi_1 _1313_ (.A1(_0143_),
    .A2(net173),
    .Y(_0103_),
    .B1(_0536_));
 sg13g2_o21ai_1 _1314_ (.B1(net195),
    .Y(_0537_),
    .A1(\desk_clock.input_debounce.en_12h_mode_reg[0] ),
    .A2(net169));
 sg13g2_a21oi_1 _1315_ (.A1(_0141_),
    .A2(net169),
    .Y(_0104_),
    .B1(_0537_));
 sg13g2_o21ai_1 _1316_ (.B1(net195),
    .Y(_0538_),
    .A1(net265),
    .A2(net169));
 sg13g2_a21oi_1 _1317_ (.A1(_0140_),
    .A2(net169),
    .Y(_0105_),
    .B1(_0538_));
 sg13g2_o21ai_1 _1318_ (.B1(net195),
    .Y(_0539_),
    .A1(net270),
    .A2(net169));
 sg13g2_a21oi_1 _1319_ (.A1(_0139_),
    .A2(net169),
    .Y(_0106_),
    .B1(_0539_));
 sg13g2_o21ai_1 _1320_ (.B1(net196),
    .Y(_0540_),
    .A1(net281),
    .A2(net172));
 sg13g2_a21oi_1 _1321_ (.A1(_0138_),
    .A2(net172),
    .Y(_0107_),
    .B1(_0540_));
 sg13g2_o21ai_1 _1322_ (.B1(net197),
    .Y(_0541_),
    .A1(\desk_clock.input_debounce.en_12h_mode_reg[4] ),
    .A2(net173));
 sg13g2_a21oi_1 _1323_ (.A1(_0136_),
    .A2(net173),
    .Y(_0108_),
    .B1(_0541_));
 sg13g2_o21ai_1 _1324_ (.B1(net197),
    .Y(_0542_),
    .A1(net243),
    .A2(net173));
 sg13g2_a21oi_1 _1325_ (.A1(_0137_),
    .A2(net173),
    .Y(_0109_),
    .B1(_0542_));
 sg13g2_nor2b_2 _1326_ (.A(\desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold ),
    .B_N(net208),
    .Y(_0543_));
 sg13g2_o21ai_1 _1327_ (.B1(net197),
    .Y(_0544_),
    .A1(\desk_clock.clk_gen_inst.refclk_div[0] ),
    .A2(_0543_));
 sg13g2_a21oi_1 _1328_ (.A1(_0135_),
    .A2(_0543_),
    .Y(_0110_),
    .B1(_0544_));
 sg13g2_a21oi_1 _1329_ (.A1(\desk_clock.clk_gen_inst.refclk_div[0] ),
    .A2(_0543_),
    .Y(_0545_),
    .B1(net250));
 sg13g2_nand3_1 _1330_ (.B(\desk_clock.clk_gen_inst.refclk_div[0] ),
    .C(_0543_),
    .A(net250),
    .Y(_0546_));
 sg13g2_nand2_1 _1331_ (.Y(_0547_),
    .A(net197),
    .B(_0546_));
 sg13g2_nor2_1 _1332_ (.A(net251),
    .B(_0547_),
    .Y(_0111_));
 sg13g2_nor2b_1 _1333_ (.A(net282),
    .B_N(_0546_),
    .Y(_0548_));
 sg13g2_and4_1 _1334_ (.A(net282),
    .B(net250),
    .C(net330),
    .D(_0543_),
    .X(_0549_));
 sg13g2_nor3_1 _1335_ (.A(net185),
    .B(net283),
    .C(_0549_),
    .Y(_0112_));
 sg13g2_nor2_1 _1336_ (.A(net245),
    .B(net331),
    .Y(_0550_));
 sg13g2_and2_1 _1337_ (.A(net245),
    .B(_0549_),
    .X(_0551_));
 sg13g2_nor3_1 _1338_ (.A(net184),
    .B(_0550_),
    .C(_0551_),
    .Y(_0113_));
 sg13g2_xnor2_1 _1339_ (.Y(_0552_),
    .A(net355),
    .B(_0551_));
 sg13g2_nor2_1 _1340_ (.A(net185),
    .B(_0552_),
    .Y(_0114_));
 sg13g2_a21oi_1 _1341_ (.A1(\desk_clock.clk_gen_inst.refclk_div[4] ),
    .A2(_0551_),
    .Y(_0553_),
    .B1(net225));
 sg13g2_nand3_1 _1342_ (.B(\desk_clock.clk_gen_inst.refclk_div[4] ),
    .C(_0551_),
    .A(net225),
    .Y(_0554_));
 sg13g2_nand2_1 _1343_ (.Y(_0555_),
    .A(net198),
    .B(_0554_));
 sg13g2_nor2_1 _1344_ (.A(net226),
    .B(_0555_),
    .Y(_0115_));
 sg13g2_or2_1 _1345_ (.X(_0556_),
    .B(_0554_),
    .A(_0134_));
 sg13g2_nand2_1 _1346_ (.Y(_0557_),
    .A(net194),
    .B(_0556_));
 sg13g2_a21oi_1 _1347_ (.A1(_0134_),
    .A2(_0554_),
    .Y(_0116_),
    .B1(_0557_));
 sg13g2_and2_1 _1348_ (.A(_0133_),
    .B(_0556_),
    .X(_0558_));
 sg13g2_nor2_2 _1349_ (.A(_0133_),
    .B(_0556_),
    .Y(_0559_));
 sg13g2_nor3_1 _1350_ (.A(net184),
    .B(_0558_),
    .C(_0559_),
    .Y(_0117_));
 sg13g2_xnor2_1 _1351_ (.Y(_0560_),
    .A(net334),
    .B(_0559_));
 sg13g2_nor2_1 _1352_ (.A(net184),
    .B(net335),
    .Y(_0118_));
 sg13g2_a21oi_1 _1353_ (.A1(\desk_clock.clk_gen_inst.refclk_div[8] ),
    .A2(_0559_),
    .Y(_0561_),
    .B1(net218));
 sg13g2_nand3_1 _1354_ (.B(net334),
    .C(_0559_),
    .A(net218),
    .Y(_0562_));
 sg13g2_nand2_1 _1355_ (.Y(_0563_),
    .A(net194),
    .B(_0562_));
 sg13g2_nor2_1 _1356_ (.A(net219),
    .B(_0563_),
    .Y(_0119_));
 sg13g2_and2_1 _1357_ (.A(_0132_),
    .B(_0562_),
    .X(_0564_));
 sg13g2_nor2_2 _1358_ (.A(_0132_),
    .B(_0562_),
    .Y(_0565_));
 sg13g2_nor3_1 _1359_ (.A(net184),
    .B(_0564_),
    .C(net327),
    .Y(_0120_));
 sg13g2_xnor2_1 _1360_ (.Y(_0566_),
    .A(net313),
    .B(net327));
 sg13g2_nor2_1 _1361_ (.A(net184),
    .B(_0566_),
    .Y(_0121_));
 sg13g2_a21oi_1 _1362_ (.A1(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .A2(_0565_),
    .Y(_0567_),
    .B1(net215));
 sg13g2_nand3_1 _1363_ (.B(net313),
    .C(_0565_),
    .A(net215),
    .Y(_0568_));
 sg13g2_nand2_1 _1364_ (.Y(_0569_),
    .A(net194),
    .B(_0568_));
 sg13g2_nor2_1 _1365_ (.A(net216),
    .B(_0569_),
    .Y(_0122_));
 sg13g2_or2_1 _1366_ (.X(_0570_),
    .B(_0568_),
    .A(_0131_));
 sg13g2_nand2_1 _1367_ (.Y(_0571_),
    .A(net193),
    .B(_0570_));
 sg13g2_a21oi_1 _1368_ (.A1(_0131_),
    .A2(net328),
    .Y(_0123_),
    .B1(_0571_));
 sg13g2_o21ai_1 _1369_ (.B1(net194),
    .Y(_0572_),
    .A1(_0130_),
    .A2(_0570_));
 sg13g2_a21oi_1 _1370_ (.A1(_0130_),
    .A2(_0570_),
    .Y(_0124_),
    .B1(_0572_));
 sg13g2_and2_1 _1371_ (.A(net313),
    .B(net194),
    .X(_0125_));
 sg13g2_and2_1 _1372_ (.A(net197),
    .B(net208),
    .X(_0126_));
 sg13g2_and2_1 _1373_ (.A(net245),
    .B(net198),
    .X(_0127_));
 sg13g2_nor2_1 _1374_ (.A(_0130_),
    .B(net185),
    .Y(_0128_));
 sg13g2_o21ai_1 _1375_ (.B1(_0244_),
    .Y(_0573_),
    .A1(net363),
    .A2(_0242_));
 sg13g2_inv_1 _1376_ (.Y(_0129_),
    .A(_0573_));
 sg13g2_dfrbp_1 _1377_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net129),
    .D(_0008_),
    .Q_N(_0687_),
    .Q(\desk_clock.refclk_sync_inst.refclk_sync_reg[0] ));
 sg13g2_dfrbp_1 _1378_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net53),
    .D(_0009_),
    .Q_N(_0686_),
    .Q(\desk_clock.clk_gen_inst.i_refclk ));
 sg13g2_dfrbp_1 _1379_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net52),
    .D(net360),
    .Q_N(_0685_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[0] ));
 sg13g2_dfrbp_1 _1380_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0011_),
    .Q_N(_0684_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[1] ));
 sg13g2_dfrbp_1 _1381_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0012_),
    .Q_N(_0683_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[2] ));
 sg13g2_dfrbp_1 _1382_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0013_),
    .Q_N(_0682_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[3] ));
 sg13g2_dfrbp_1 _1383_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0014_),
    .Q_N(_0681_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[7] ));
 sg13g2_dfrbp_1 _1384_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net42),
    .D(_0015_),
    .Q_N(_0680_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[0] ));
 sg13g2_dfrbp_1 _1385_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net40),
    .D(net247),
    .Q_N(_0679_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[1] ));
 sg13g2_dfrbp_1 _1386_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net38),
    .D(net352),
    .Q_N(_0678_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[2] ));
 sg13g2_dfrbp_1 _1387_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net36),
    .D(net235),
    .Q_N(_0677_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[3] ));
 sg13g2_dfrbp_1 _1388_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0019_),
    .Q_N(_0676_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[4] ));
 sg13g2_dfrbp_1 _1389_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net32),
    .D(net301),
    .Q_N(_0675_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[5] ));
 sg13g2_dfrbp_1 _1390_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net30),
    .D(_0021_),
    .Q_N(_0674_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[6] ));
 sg13g2_dfrbp_1 _1391_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net28),
    .D(net286),
    .Q_N(_0673_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[7] ));
 sg13g2_dfrbp_1 _1392_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net26),
    .D(net276),
    .Q_N(_0672_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[8] ));
 sg13g2_dfrbp_1 _1393_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net146),
    .D(net239),
    .Q_N(_0671_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[9] ));
 sg13g2_dfrbp_1 _1394_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net144),
    .D(net212),
    .Q_N(_0670_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[10] ));
 sg13g2_dfrbp_1 _1395_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net142),
    .D(net231),
    .Q_N(_0669_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[11] ));
 sg13g2_dfrbp_1 _1396_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net140),
    .D(net207),
    .Q_N(_0000_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[0] ));
 sg13g2_dfrbp_1 _1397_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net138),
    .D(net272),
    .Q_N(_0668_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ));
 sg13g2_dfrbp_1 _1398_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net136),
    .D(net242),
    .Q_N(_0667_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ));
 sg13g2_dfrbp_1 _1399_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net134),
    .D(_0030_),
    .Q_N(_0666_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ));
 sg13g2_dfrbp_1 _1400_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net132),
    .D(_0031_),
    .Q_N(_0665_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ));
 sg13g2_dfrbp_1 _1401_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net130),
    .D(net338),
    .Q_N(_0664_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ));
 sg13g2_dfrbp_1 _1402_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net128),
    .D(net269),
    .Q_N(_0663_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[0] ));
 sg13g2_dfrbp_1 _1403_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net126),
    .D(net259),
    .Q_N(_0662_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ));
 sg13g2_dfrbp_1 _1404_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net124),
    .D(net345),
    .Q_N(_0661_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ));
 sg13g2_dfrbp_1 _1405_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net122),
    .D(net354),
    .Q_N(_0660_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ));
 sg13g2_dfrbp_1 _1406_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net120),
    .D(net233),
    .Q_N(_0659_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ));
 sg13g2_dfrbp_1 _1407_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net118),
    .D(net347),
    .Q_N(_0658_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[5] ));
 sg13g2_dfrbp_1 _1408_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net116),
    .D(net261),
    .Q_N(_0657_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ));
 sg13g2_dfrbp_1 _1409_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net114),
    .D(net274),
    .Q_N(_0656_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[1] ));
 sg13g2_dfrbp_1 _1410_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net112),
    .D(net278),
    .Q_N(_0655_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[2] ));
 sg13g2_dfrbp_1 _1411_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net110),
    .D(net280),
    .Q_N(_0654_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[3] ));
 sg13g2_dfrbp_1 _1412_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net108),
    .D(net303),
    .Q_N(_0653_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[4] ));
 sg13g2_dfrbp_1 _1413_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net106),
    .D(net292),
    .Q_N(_0652_),
    .Q(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ));
 sg13g2_dfrbp_1 _1414_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net104),
    .D(net325),
    .Q_N(_0003_),
    .Q(\desk_clock.display_inst.state[0] ));
 sg13g2_dfrbp_1 _1415_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net102),
    .D(net394),
    .Q_N(_0651_),
    .Q(\desk_clock.display_inst.state[1] ));
 sg13g2_dfrbp_1 _1416_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net100),
    .D(net389),
    .Q_N(_0650_),
    .Q(\desk_clock.display_inst.state[2] ));
 sg13g2_dfrbp_1 _1417_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net98),
    .D(net24),
    .Q_N(_0649_),
    .Q(\desk_clock.display_inst.state[3] ));
 sg13g2_dfrbp_1 _1418_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net96),
    .D(net373),
    .Q_N(_0004_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[0] ));
 sg13g2_dfrbp_1 _1419_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net94),
    .D(_0050_),
    .Q_N(_0648_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[1] ));
 sg13g2_dfrbp_1 _1420_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net92),
    .D(net392),
    .Q_N(_0001_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[2] ));
 sg13g2_dfrbp_1 _1421_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net90),
    .D(net205),
    .Q_N(_0647_),
    .Q(\desk_clock.display_inst.display_settings.transfer_state[3] ));
 sg13g2_dfrbp_1 _1422_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net88),
    .D(_0053_),
    .Q_N(_0646_),
    .Q(\desk_clock.display_inst.disp_driver.i_data[4] ));
 sg13g2_dfrbp_1 _1423_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net86),
    .D(_0054_),
    .Q_N(_0645_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[0] ));
 sg13g2_dfrbp_1 _1424_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net84),
    .D(net350),
    .Q_N(_0644_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[1] ));
 sg13g2_dfrbp_1 _1425_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net82),
    .D(_0056_),
    .Q_N(_0643_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[2] ));
 sg13g2_dfrbp_1 _1426_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0057_),
    .Q_N(_0642_),
    .Q(\desk_clock.display_inst.disp_driver.i_addr[3] ));
 sg13g2_dfrbp_1 _1427_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0058_),
    .Q_N(_0641_),
    .Q(\desk_clock.display_control_inst.display_update ));
 sg13g2_dfrbp_1 _1428_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net77),
    .D(_0059_),
    .Q_N(_0640_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[1] ));
 sg13g2_dfrbp_1 _1429_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net75),
    .D(net264),
    .Q_N(_0639_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[2] ));
 sg13g2_dfrbp_1 _1430_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net73),
    .D(_0061_),
    .Q_N(_0638_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[3] ));
 sg13g2_dfrbp_1 _1431_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0062_),
    .Q_N(_0637_),
    .Q(\desk_clock.display_inst.disp_driver.transfer_state[4] ));
 sg13g2_dfrbp_1 _1432_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net69),
    .D(_0063_),
    .Q_N(_0636_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[12] ));
 sg13g2_dfrbp_1 _1433_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net67),
    .D(_0064_),
    .Q_N(_0635_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[13] ));
 sg13g2_dfrbp_1 _1434_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net65),
    .D(net237),
    .Q_N(_0634_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[14] ));
 sg13g2_dfrbp_1 _1435_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net63),
    .D(net249),
    .Q_N(_0633_),
    .Q(\desk_clock.display_inst.disp_driver.data_reg[15] ));
 sg13g2_dfrbp_1 _1436_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net61),
    .D(_0067_),
    .Q_N(_0002_),
    .Q(\desk_clock.display_control_inst.o_write_config ));
 sg13g2_dfrbp_1 _1437_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0068_),
    .Q_N(_0632_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_slow_clk.sig_hold ));
 sg13g2_dfrbp_1 _1438_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0069_),
    .Q_N(_0631_),
    .Q(\desk_clock.clk_seconds[0] ));
 sg13g2_dfrbp_1 _1439_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net56),
    .D(net297),
    .Q_N(_0630_),
    .Q(\desk_clock.clk_seconds[1] ));
 sg13g2_dfrbp_1 _1440_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net54),
    .D(_0071_),
    .Q_N(_0629_),
    .Q(\desk_clock.clk_seconds[2] ));
 sg13g2_dfrbp_1 _1441_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net49),
    .D(_0072_),
    .Q_N(_0628_),
    .Q(\desk_clock.clk_seconds[3] ));
 sg13g2_dfrbp_1 _1442_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net45),
    .D(_0073_),
    .Q_N(_0627_),
    .Q(\desk_clock.clk_seconds[4] ));
 sg13g2_dfrbp_1 _1443_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net41),
    .D(_0074_),
    .Q_N(_0626_),
    .Q(\desk_clock.clk_seconds[5] ));
 sg13g2_dfrbp_1 _1444_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0075_),
    .Q_N(_0625_),
    .Q(\desk_clock.clk_minutes[0] ));
 sg13g2_dfrbp_1 _1445_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net33),
    .D(net375),
    .Q_N(_0624_),
    .Q(\desk_clock.clk_minutes[1] ));
 sg13g2_dfrbp_1 _1446_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net29),
    .D(_0077_),
    .Q_N(_0623_),
    .Q(\desk_clock.clk_minutes[2] ));
 sg13g2_dfrbp_1 _1447_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net25),
    .D(_0078_),
    .Q_N(_0622_),
    .Q(\desk_clock.clk_minutes[3] ));
 sg13g2_dfrbp_1 _1448_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net143),
    .D(_0079_),
    .Q_N(_0621_),
    .Q(\desk_clock.clk_minutes[4] ));
 sg13g2_dfrbp_1 _1449_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net139),
    .D(_0080_),
    .Q_N(_0620_),
    .Q(\desk_clock.clk_minutes[5] ));
 sg13g2_dfrbp_1 _1450_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net135),
    .D(net384),
    .Q_N(_0619_),
    .Q(\desk_clock.clk_hours[0] ));
 sg13g2_dfrbp_1 _1451_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net131),
    .D(net381),
    .Q_N(_0618_),
    .Q(\desk_clock.clk_hours[1] ));
 sg13g2_dfrbp_1 _1452_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net127),
    .D(net400),
    .Q_N(_0006_),
    .Q(\desk_clock.clk_hours[2] ));
 sg13g2_dfrbp_1 _1453_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net123),
    .D(net404),
    .Q_N(_0617_),
    .Q(\desk_clock.clk_hours[3] ));
 sg13g2_dfrbp_1 _1454_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net119),
    .D(net402),
    .Q_N(_0005_),
    .Q(\desk_clock.clk_hours[4] ));
 sg13g2_dfrbp_1 _1455_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net115),
    .D(net317),
    .Q_N(_0616_),
    .Q(\desk_clock.input_debounce.fast_set_reg[0] ));
 sg13g2_dfrbp_1 _1456_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net111),
    .D(net210),
    .Q_N(_0615_),
    .Q(\desk_clock.input_debounce.fast_set_reg[1] ));
 sg13g2_dfrbp_1 _1457_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net107),
    .D(_0088_),
    .Q_N(_0614_),
    .Q(\desk_clock.input_debounce.fast_set_reg[2] ));
 sg13g2_dfrbp_1 _1458_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net103),
    .D(_0089_),
    .Q_N(_0613_),
    .Q(\desk_clock.input_debounce.fast_set_reg[3] ));
 sg13g2_dfrbp_1 _1459_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net99),
    .D(net214),
    .Q_N(_0612_),
    .Q(\desk_clock.input_debounce.fast_set_reg[4] ));
 sg13g2_dfrbp_1 _1460_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net95),
    .D(_0091_),
    .Q_N(_0611_),
    .Q(\desk_clock.input_debounce.fast_set_reg[5] ));
 sg13g2_dfrbp_1 _1461_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net91),
    .D(net308),
    .Q_N(_0610_),
    .Q(\desk_clock.input_debounce.set_hours_reg[0] ));
 sg13g2_dfrbp_1 _1462_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net87),
    .D(net290),
    .Q_N(_0609_),
    .Q(\desk_clock.input_debounce.set_hours_reg[1] ));
 sg13g2_dfrbp_1 _1463_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net83),
    .D(_0094_),
    .Q_N(_0608_),
    .Q(\desk_clock.input_debounce.set_hours_reg[2] ));
 sg13g2_dfrbp_1 _1464_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net79),
    .D(net254),
    .Q_N(_0607_),
    .Q(\desk_clock.input_debounce.set_hours_reg[3] ));
 sg13g2_dfrbp_1 _1465_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net74),
    .D(_0096_),
    .Q_N(_0606_),
    .Q(\desk_clock.input_debounce.set_hours_reg[4] ));
 sg13g2_dfrbp_1 _1466_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0097_),
    .Q_N(_0605_),
    .Q(\desk_clock.input_debounce.set_hours_reg[5] ));
 sg13g2_dfrbp_1 _1467_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net66),
    .D(net257),
    .Q_N(_0604_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[0] ));
 sg13g2_dfrbp_1 _1468_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net62),
    .D(_0099_),
    .Q_N(_0603_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[1] ));
 sg13g2_dfrbp_1 _1469_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net57),
    .D(_0100_),
    .Q_N(_0602_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[2] ));
 sg13g2_dfrbp_1 _1470_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net51),
    .D(_0101_),
    .Q_N(_0601_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[3] ));
 sg13g2_dfrbp_1 _1471_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net43),
    .D(net224),
    .Q_N(_0600_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[4] ));
 sg13g2_dfrbp_1 _1472_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net35),
    .D(_0103_),
    .Q_N(_0599_),
    .Q(\desk_clock.input_debounce.set_minutes_reg[5] ));
 sg13g2_dfrbp_1 _1473_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net27),
    .D(net266),
    .Q_N(_0598_),
    .Q(\desk_clock.input_debounce.en_12h_mode_reg[0] ));
 sg13g2_dfrbp_1 _1474_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net141),
    .D(_0105_),
    .Q_N(_0597_),
    .Q(\desk_clock.input_debounce.en_12h_mode_reg[1] ));
 sg13g2_dfrbp_1 _1475_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net133),
    .D(_0106_),
    .Q_N(_0596_),
    .Q(\desk_clock.input_debounce.en_12h_mode_reg[2] ));
 sg13g2_dfrbp_1 _1476_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net125),
    .D(_0107_),
    .Q_N(_0595_),
    .Q(\desk_clock.input_debounce.en_12h_mode_reg[3] ));
 sg13g2_dfrbp_1 _1477_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net117),
    .D(net244),
    .Q_N(_0594_),
    .Q(\desk_clock.input_debounce.en_12h_mode_reg[4] ));
 sg13g2_dfrbp_1 _1478_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net109),
    .D(_0109_),
    .Q_N(_0593_),
    .Q(\desk_clock.input_debounce.en_12h_mode_reg[5] ));
 sg13g2_dfrbp_1 _1479_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net101),
    .D(net202),
    .Q_N(_0007_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[0] ));
 sg13g2_dfrbp_1 _1480_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net93),
    .D(net252),
    .Q_N(_0592_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[1] ));
 sg13g2_dfrbp_1 _1481_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net85),
    .D(net284),
    .Q_N(_0591_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[2] ));
 sg13g2_dfrbp_1 _1482_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net76),
    .D(_0113_),
    .Q_N(_0590_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[3] ));
 sg13g2_dfrbp_1 _1483_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net68),
    .D(_0114_),
    .Q_N(_0589_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[4] ));
 sg13g2_dfrbp_1 _1484_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net60),
    .D(net227),
    .Q_N(_0588_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[5] ));
 sg13g2_dfrbp_1 _1485_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net47),
    .D(net229),
    .Q_N(_0587_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[6] ));
 sg13g2_dfrbp_1 _1486_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net31),
    .D(_0117_),
    .Q_N(_0586_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[7] ));
 sg13g2_dfrbp_1 _1487_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net137),
    .D(_0118_),
    .Q_N(_0585_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[8] ));
 sg13g2_dfrbp_1 _1488_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net121),
    .D(net220),
    .Q_N(_0584_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[9] ));
 sg13g2_dfrbp_1 _1489_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net105),
    .D(_0120_),
    .Q_N(_0583_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[10] ));
 sg13g2_dfrbp_1 _1490_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net89),
    .D(_0121_),
    .Q_N(_0582_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[11] ));
 sg13g2_dfrbp_1 _1491_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net72),
    .D(net217),
    .Q_N(_0581_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[12] ));
 sg13g2_dfrbp_1 _1492_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net55),
    .D(_0123_),
    .Q_N(_0580_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[13] ));
 sg13g2_dfrbp_1 _1493_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net145),
    .D(_0124_),
    .Q_N(_0579_),
    .Q(\desk_clock.clk_gen_inst.refclk_div[14] ));
 sg13g2_dfrbp_1 _1494_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net113),
    .D(_0125_),
    .Q_N(_0578_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_fast_clk.sig_hold ));
 sg13g2_dfrbp_1 _1495_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0126_),
    .Q_N(_0577_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_refclk.sig_hold ));
 sg13g2_dfrbp_1 _1496_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net81),
    .D(_0127_),
    .Q_N(_0576_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_debounce_clk.sig_hold ));
 sg13g2_dfrbp_1 _1497_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0128_),
    .Q_N(_0575_),
    .Q(\desk_clock.clk_gen_inst.stb_gen_1hz.sig_hold ));
 sg13g2_dfrbp_1 _1498_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0129_),
    .Q_N(_0574_),
    .Q(\desk_clock.display_inst.display_settings.write_config ));
 sg13g2_tiehi _1392__26 (.L_HI(net26));
 sg13g2_tiehi _1473__27 (.L_HI(net27));
 sg13g2_tiehi _1391__28 (.L_HI(net28));
 sg13g2_tiehi _1446__29 (.L_HI(net29));
 sg13g2_tiehi _1390__30 (.L_HI(net30));
 sg13g2_tiehi _1486__31 (.L_HI(net31));
 sg13g2_tiehi _1389__32 (.L_HI(net32));
 sg13g2_tiehi _1445__33 (.L_HI(net33));
 sg13g2_tiehi _1388__34 (.L_HI(net34));
 sg13g2_tiehi _1472__35 (.L_HI(net35));
 sg13g2_tiehi _1387__36 (.L_HI(net36));
 sg13g2_tiehi _1444__37 (.L_HI(net37));
 sg13g2_tiehi _1386__38 (.L_HI(net38));
 sg13g2_tiehi _1498__39 (.L_HI(net39));
 sg13g2_tiehi _1385__40 (.L_HI(net40));
 sg13g2_tiehi _1443__41 (.L_HI(net41));
 sg13g2_tiehi _1384__42 (.L_HI(net42));
 sg13g2_tiehi _1471__43 (.L_HI(net43));
 sg13g2_tiehi _1383__44 (.L_HI(net44));
 sg13g2_tiehi _1442__45 (.L_HI(net45));
 sg13g2_tiehi _1382__46 (.L_HI(net46));
 sg13g2_tiehi _1485__47 (.L_HI(net47));
 sg13g2_tiehi _1381__48 (.L_HI(net48));
 sg13g2_tiehi _1441__49 (.L_HI(net49));
 sg13g2_tiehi _1380__50 (.L_HI(net50));
 sg13g2_tiehi _1470__51 (.L_HI(net51));
 sg13g2_tiehi _1379__52 (.L_HI(net52));
 sg13g2_tiehi _1378__53 (.L_HI(net53));
 sg13g2_tiehi _1440__54 (.L_HI(net54));
 sg13g2_tiehi _1492__55 (.L_HI(net55));
 sg13g2_tiehi _1439__56 (.L_HI(net56));
 sg13g2_tiehi _1469__57 (.L_HI(net57));
 sg13g2_tiehi _1438__58 (.L_HI(net58));
 sg13g2_tiehi _1437__59 (.L_HI(net59));
 sg13g2_tiehi _1484__60 (.L_HI(net60));
 sg13g2_tiehi _1436__61 (.L_HI(net61));
 sg13g2_tiehi _1468__62 (.L_HI(net62));
 sg13g2_tiehi _1435__63 (.L_HI(net63));
 sg13g2_tiehi _1497__64 (.L_HI(net64));
 sg13g2_tiehi _1434__65 (.L_HI(net65));
 sg13g2_tiehi _1467__66 (.L_HI(net66));
 sg13g2_tiehi _1433__67 (.L_HI(net67));
 sg13g2_tiehi _1483__68 (.L_HI(net68));
 sg13g2_tiehi _1432__69 (.L_HI(net69));
 sg13g2_tiehi _1466__70 (.L_HI(net70));
 sg13g2_tiehi _1431__71 (.L_HI(net71));
 sg13g2_tiehi _1491__72 (.L_HI(net72));
 sg13g2_tiehi _1430__73 (.L_HI(net73));
 sg13g2_tiehi _1465__74 (.L_HI(net74));
 sg13g2_tiehi _1429__75 (.L_HI(net75));
 sg13g2_tiehi _1482__76 (.L_HI(net76));
 sg13g2_tiehi _1428__77 (.L_HI(net77));
 sg13g2_tiehi _1427__78 (.L_HI(net78));
 sg13g2_tiehi _1464__79 (.L_HI(net79));
 sg13g2_tiehi _1426__80 (.L_HI(net80));
 sg13g2_tiehi _1496__81 (.L_HI(net81));
 sg13g2_tiehi _1425__82 (.L_HI(net82));
 sg13g2_tiehi _1463__83 (.L_HI(net83));
 sg13g2_tiehi _1424__84 (.L_HI(net84));
 sg13g2_tiehi _1481__85 (.L_HI(net85));
 sg13g2_tiehi _1423__86 (.L_HI(net86));
 sg13g2_tiehi _1462__87 (.L_HI(net87));
 sg13g2_tiehi _1422__88 (.L_HI(net88));
 sg13g2_tiehi _1490__89 (.L_HI(net89));
 sg13g2_tiehi _1421__90 (.L_HI(net90));
 sg13g2_tiehi _1461__91 (.L_HI(net91));
 sg13g2_tiehi _1420__92 (.L_HI(net92));
 sg13g2_tiehi _1480__93 (.L_HI(net93));
 sg13g2_tiehi _1419__94 (.L_HI(net94));
 sg13g2_tiehi _1460__95 (.L_HI(net95));
 sg13g2_tiehi _1418__96 (.L_HI(net96));
 sg13g2_tiehi _1495__97 (.L_HI(net97));
 sg13g2_tiehi _1417__98 (.L_HI(net98));
 sg13g2_tiehi _1459__99 (.L_HI(net99));
 sg13g2_tiehi _1416__100 (.L_HI(net100));
 sg13g2_tiehi _1479__101 (.L_HI(net101));
 sg13g2_tiehi _1415__102 (.L_HI(net102));
 sg13g2_tiehi _1458__103 (.L_HI(net103));
 sg13g2_tiehi _1414__104 (.L_HI(net104));
 sg13g2_tiehi _1489__105 (.L_HI(net105));
 sg13g2_tiehi _1413__106 (.L_HI(net106));
 sg13g2_tiehi _1457__107 (.L_HI(net107));
 sg13g2_tiehi _1412__108 (.L_HI(net108));
 sg13g2_tiehi _1478__109 (.L_HI(net109));
 sg13g2_tiehi _1411__110 (.L_HI(net110));
 sg13g2_tiehi _1456__111 (.L_HI(net111));
 sg13g2_tiehi _1410__112 (.L_HI(net112));
 sg13g2_tiehi _1494__113 (.L_HI(net113));
 sg13g2_tiehi _1409__114 (.L_HI(net114));
 sg13g2_tiehi _1455__115 (.L_HI(net115));
 sg13g2_tiehi _1408__116 (.L_HI(net116));
 sg13g2_tiehi _1477__117 (.L_HI(net117));
 sg13g2_tiehi _1407__118 (.L_HI(net118));
 sg13g2_tiehi _1454__119 (.L_HI(net119));
 sg13g2_tiehi _1406__120 (.L_HI(net120));
 sg13g2_tiehi _1488__121 (.L_HI(net121));
 sg13g2_tiehi _1405__122 (.L_HI(net122));
 sg13g2_tiehi _1453__123 (.L_HI(net123));
 sg13g2_tiehi _1404__124 (.L_HI(net124));
 sg13g2_tiehi _1476__125 (.L_HI(net125));
 sg13g2_tiehi _1403__126 (.L_HI(net126));
 sg13g2_tiehi _1452__127 (.L_HI(net127));
 sg13g2_tiehi _1402__128 (.L_HI(net128));
 sg13g2_tiehi _1377__129 (.L_HI(net129));
 sg13g2_tiehi _1401__130 (.L_HI(net130));
 sg13g2_tiehi _1451__131 (.L_HI(net131));
 sg13g2_tiehi _1400__132 (.L_HI(net132));
 sg13g2_tiehi _1475__133 (.L_HI(net133));
 sg13g2_tiehi _1399__134 (.L_HI(net134));
 sg13g2_tiehi _1450__135 (.L_HI(net135));
 sg13g2_tiehi _1398__136 (.L_HI(net136));
 sg13g2_tiehi _1487__137 (.L_HI(net137));
 sg13g2_tiehi _1397__138 (.L_HI(net138));
 sg13g2_tiehi _1449__139 (.L_HI(net139));
 sg13g2_tiehi _1396__140 (.L_HI(net140));
 sg13g2_tiehi _1474__141 (.L_HI(net141));
 sg13g2_tiehi _1395__142 (.L_HI(net142));
 sg13g2_tiehi _1448__143 (.L_HI(net143));
 sg13g2_tiehi _1394__144 (.L_HI(net144));
 sg13g2_tiehi _1493__145 (.L_HI(net145));
 sg13g2_tiehi _1393__146 (.L_HI(net146));
 sg13g2_tiehi tt_um_digital_clock_example_147 (.L_HI(net147));
 sg13g2_tiehi tt_um_digital_clock_example_148 (.L_HI(net148));
 sg13g2_tiehi tt_um_digital_clock_example_149 (.L_HI(net149));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_tielo tt_um_digital_clock_example_7 (.L_LO(net7));
 sg13g2_tielo tt_um_digital_clock_example_8 (.L_LO(net8));
 sg13g2_tielo tt_um_digital_clock_example_9 (.L_LO(net9));
 sg13g2_tielo tt_um_digital_clock_example_10 (.L_LO(net10));
 sg13g2_tielo tt_um_digital_clock_example_11 (.L_LO(net11));
 sg13g2_tielo tt_um_digital_clock_example_12 (.L_LO(net12));
 sg13g2_tielo tt_um_digital_clock_example_13 (.L_LO(net13));
 sg13g2_tielo tt_um_digital_clock_example_14 (.L_LO(net14));
 sg13g2_tielo tt_um_digital_clock_example_15 (.L_LO(net15));
 sg13g2_tielo tt_um_digital_clock_example_16 (.L_LO(net16));
 sg13g2_tielo tt_um_digital_clock_example_17 (.L_LO(net17));
 sg13g2_tielo tt_um_digital_clock_example_18 (.L_LO(net18));
 sg13g2_tielo tt_um_digital_clock_example_19 (.L_LO(net19));
 sg13g2_tielo tt_um_digital_clock_example_20 (.L_LO(net20));
 sg13g2_tielo tt_um_digital_clock_example_21 (.L_LO(net21));
 sg13g2_tielo tt_um_digital_clock_example_22 (.L_LO(net22));
 sg13g2_tielo tt_um_digital_clock_example_23 (.L_LO(net23));
 sg13g2_tielo _1417__24 (.L_LO(net24));
 sg13g2_tiehi _1447__25 (.L_HI(net25));
 sg13g2_buf_1 _1643_ (.A(\desk_clock.display_inst.disp_driver.o_serial_load ),
    .X(uio_out[0]));
 sg13g2_buf_1 _1644_ (.A(\desk_clock.display_inst.disp_driver.data_reg[15] ),
    .X(uio_out[1]));
 sg13g2_buf_1 _1645_ (.A(\desk_clock.display_inst.disp_driver.o_serial_clk ),
    .X(uio_out[3]));
 sg13g2_buf_2 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0255_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(_0233_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0323_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0322_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_0363_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(net162),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(net161),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0364_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0198_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0181_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_0181_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_0180_),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(_0180_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(net176),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(net176),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net176),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(net175),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net175),
    .X(net173));
 sg13g2_buf_1 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(_0518_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_0191_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(\desk_clock.clk_hours[4] ),
    .X(net178));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(net388));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net393));
 sg13g2_buf_1 fanout181 (.A(\desk_clock.display_inst.state[1] ),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net348),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net186));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(_0177_));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(net192));
 sg13g2_buf_2 fanout188 (.A(net192),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net200),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net200),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net200),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net199),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net199),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net200),
    .X(net199));
 sg13g2_buf_1 fanout200 (.A(rst_n),
    .X(net200));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_tielo tt_um_digital_clock_example_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0007_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0110_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold3 (.A(\desk_clock.refclk_sync_inst.refclk_sync_reg[0] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0001_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0052_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0027_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold8 (.A(\desk_clock.clk_gen_inst.i_refclk ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold9 (.A(\desk_clock.input_debounce.fast_set_reg[2] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0087_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold11 (.A(\desk_clock.display_inst.disp_driver.data_reg[9] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0025_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold13 (.A(\desk_clock.input_debounce.fast_set_reg[5] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0090_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold15 (.A(\desk_clock.clk_gen_inst.refclk_div[12] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0567_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0122_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold18 (.A(\desk_clock.clk_gen_inst.refclk_div[9] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0561_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0119_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold21 (.A(\desk_clock.display_inst.disp_driver.data_reg[0] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0326_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold23 (.A(\desk_clock.input_debounce.set_minutes_reg[5] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0102_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold25 (.A(\desk_clock.clk_gen_inst.refclk_div[5] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0553_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0115_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold28 (.A(\desk_clock.clk_gen_inst.refclk_div[6] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0116_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold30 (.A(\desk_clock.display_inst.disp_driver.data_reg[10] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0026_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold32 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0037_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold34 (.A(\desk_clock.display_inst.disp_driver.data_reg[2] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0018_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold36 (.A(\desk_clock.display_inst.disp_driver.data_reg[13] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0065_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold38 (.A(\desk_clock.display_inst.disp_driver.data_reg[8] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0024_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold40 (.A(\desk_clock.display_inst.disp_driver.data_reg[12] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold41 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[1] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0029_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold43 (.A(\desk_clock.input_debounce.en_12h_mode_reg[5] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0108_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold45 (.A(\desk_clock.clk_gen_inst.refclk_div[3] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold46 (.A(\desk_clock.display_inst.disp_driver.i_data[1] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0016_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold48 (.A(\desk_clock.display_inst.disp_driver.data_reg[15] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0066_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold50 (.A(\desk_clock.clk_gen_inst.refclk_div[1] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0545_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0111_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold53 (.A(\desk_clock.input_debounce.set_hours_reg[4] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0095_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold55 (.A(\desk_clock.display_inst.disp_driver.data_reg[11] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold56 (.A(\desk_clock.input_debounce.set_minutes_reg[1] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0098_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold58 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[1] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0034_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold60 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[0] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0039_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold62 (.A(\desk_clock.display_inst.disp_driver.transfer_state[2] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0444_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0060_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold65 (.A(\desk_clock.input_debounce.en_12h_mode_reg[1] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0104_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold67 (.A(\desk_clock.input_debounce.set_hours_reg[5] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold68 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[0] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0033_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold70 (.A(\desk_clock.input_debounce.en_12h_mode_reg[2] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold71 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[0] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0028_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold73 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[1] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0040_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold75 (.A(\desk_clock.display_inst.disp_driver.data_reg[7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0023_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold77 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[2] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0041_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold79 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[3] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0042_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold81 (.A(\desk_clock.input_debounce.en_12h_mode_reg[3] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold82 (.A(\desk_clock.clk_gen_inst.refclk_div[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0548_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0112_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold85 (.A(\desk_clock.display_inst.disp_driver.data_reg[6] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0022_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold87 (.A(\desk_clock.clk_minutes[2] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0489_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold89 (.A(\desk_clock.input_debounce.set_hours_reg[2] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0093_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold91 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[5] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0044_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold93 (.A(\desk_clock.input_debounce.set_minutes_reg[2] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold94 (.A(\desk_clock.input_debounce.set_hours_reg[3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold95 (.A(\desk_clock.clk_seconds[1] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0461_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0070_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold98 (.A(\desk_clock.input_debounce.fast_set_reg[3] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold99 (.A(\desk_clock.display_inst.disp_driver.data_reg[4] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0339_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0020_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold102 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_seconds[4] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0043_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold104 (.A(\desk_clock.clk_gen_inst.refclk_div[13] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold105 (.A(\desk_clock.clk_minutes[4] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0497_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold107 (.A(\desk_clock.input_debounce.set_hours_reg[1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0092_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold109 (.A(\desk_clock.input_debounce.set_minutes_reg[3] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold110 (.A(\desk_clock.display_inst.disp_driver.data_reg[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0341_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold112 (.A(\desk_clock.clk_gen_inst.refclk_div[14] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold113 (.A(\desk_clock.clk_gen_inst.refclk_div[11] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold114 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[3] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0379_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold116 (.A(\desk_clock.input_debounce.fast_set_reg[1] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0086_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold118 (.A(\desk_clock.display_inst.disp_driver.data_reg[3] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0337_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold120 (.A(\desk_clock.input_debounce.fast_set_reg[4] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold121 (.A(\desk_clock.input_debounce.en_12h_mode_reg[4] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold122 (.A(\desk_clock.clk_seconds[5] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0472_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0002_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0045_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold126 (.A(\desk_clock.clk_gen_inst.refclk_div[10] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0565_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0568_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold129 (.A(\desk_clock.input_debounce.set_minutes_reg[4] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold130 (.A(\desk_clock.clk_gen_inst.refclk_div[0] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0549_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold132 (.A(\desk_clock.display_inst.disp_driver.transfer_state[3] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0446_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold134 (.A(\desk_clock.clk_gen_inst.refclk_div[8] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0560_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold136 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[4] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0381_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0032_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold139 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.hours_int[2] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0374_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold141 (.A(\desk_clock.display_inst.disp_driver.i_addr[3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold142 (.A(\desk_clock.display_inst.disp_driver.i_addr[2] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold143 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[2] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0384_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0035_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold146 (.A(\desk_clock.clk_minutes[5] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0038_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold148 (.A(\desk_clock.display_inst.state[0] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold149 (.A(\desk_clock.display_inst.disp_driver.i_addr[1] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0055_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold151 (.A(\desk_clock.display_inst.disp_driver.i_data[2] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0017_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold153 (.A(\desk_clock.display_inst.clock_to_bcd_conv_inst.i_minutes[3] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0036_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold155 (.A(\desk_clock.clk_gen_inst.refclk_div[4] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold156 (.A(\desk_clock.display_inst.disp_driver.i_data[7] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold157 (.A(\desk_clock.display_inst.disp_driver.i_addr[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold158 (.A(\desk_clock.clk_gen_inst.refclk_div[7] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold159 (.A(\desk_clock.display_inst.disp_driver.i_data[0] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0010_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold161 (.A(\desk_clock.display_inst.disp_driver.transfer_state[1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0442_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold163 (.A(\desk_clock.display_inst.display_settings.write_config ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold164 (.A(\desk_clock.display_control_inst.o_write_config ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold165 (.A(\desk_clock.clk_seconds[3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0469_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold167 (.A(\desk_clock.clk_minutes[0] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold168 (.A(\desk_clock.clk_seconds[4] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold169 (.A(\desk_clock.display_inst.disp_driver.i_data[4] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold170 (.A(\desk_clock.display_inst.disp_driver.i_data[3] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0004_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0410_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0049_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold174 (.A(\desk_clock.clk_minutes[1] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0076_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold176 (.A(\desk_clock.clk_minutes[3] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold177 (.A(\desk_clock.clk_seconds[2] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0462_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold179 (.A(\desk_clock.clk_hours[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0506_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0082_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold182 (.A(\desk_clock.display_inst.state[3] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold183 (.A(\desk_clock.clk_hours[0] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0081_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold185 (.A(\desk_clock.clk_seconds[0] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0459_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold187 (.A(\desk_clock.display_inst.disp_driver.transfer_state[4] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold188 (.A(\desk_clock.display_inst.state[2] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0047_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold190 (.A(\desk_clock.display_inst.display_settings.transfer_state[1] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold191 (.A(\desk_clock.display_inst.display_settings.transfer_state[2] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0051_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold193 (.A(\desk_clock.display_inst.state[1] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0046_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold195 (.A(\desk_clock.display_control_inst.display_update ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0438_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0439_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0006_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0511_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0083_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0005_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0085_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold203 (.A(\desk_clock.clk_hours[3] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0084_),
    .X(net404));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_4 FILLER_8_119 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_decap_4 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_138 ();
 sg13g2_decap_8 FILLER_8_145 ();
 sg13g2_decap_8 FILLER_8_152 ();
 sg13g2_decap_8 FILLER_8_159 ();
 sg13g2_decap_8 FILLER_8_166 ();
 sg13g2_decap_8 FILLER_8_173 ();
 sg13g2_decap_8 FILLER_8_180 ();
 sg13g2_decap_8 FILLER_8_187 ();
 sg13g2_decap_8 FILLER_8_194 ();
 sg13g2_decap_8 FILLER_8_201 ();
 sg13g2_decap_8 FILLER_8_208 ();
 sg13g2_decap_8 FILLER_8_215 ();
 sg13g2_decap_8 FILLER_8_222 ();
 sg13g2_fill_2 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_4 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_4 FILLER_9_84 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_fill_2 FILLER_9_120 ();
 sg13g2_fill_1 FILLER_9_122 ();
 sg13g2_decap_8 FILLER_9_149 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_185 ();
 sg13g2_decap_8 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_fill_2 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_fill_2 FILLER_10_63 ();
 sg13g2_fill_1 FILLER_10_65 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_4 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_81 ();
 sg13g2_decap_4 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_96 ();
 sg13g2_fill_2 FILLER_10_157 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_192 ();
 sg13g2_decap_4 FILLER_10_196 ();
 sg13g2_fill_2 FILLER_10_226 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_285 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_4 FILLER_10_313 ();
 sg13g2_fill_2 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_fill_2 FILLER_11_93 ();
 sg13g2_fill_1 FILLER_11_95 ();
 sg13g2_decap_4 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_158 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_4 FILLER_11_223 ();
 sg13g2_fill_2 FILLER_11_227 ();
 sg13g2_fill_2 FILLER_11_237 ();
 sg13g2_fill_1 FILLER_11_239 ();
 sg13g2_fill_1 FILLER_11_284 ();
 sg13g2_fill_2 FILLER_11_290 ();
 sg13g2_fill_1 FILLER_11_296 ();
 sg13g2_fill_2 FILLER_11_305 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_58 ();
 sg13g2_decap_4 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_67 ();
 sg13g2_decap_4 FILLER_12_114 ();
 sg13g2_fill_1 FILLER_12_118 ();
 sg13g2_decap_8 FILLER_12_127 ();
 sg13g2_decap_8 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_decap_4 FILLER_12_153 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_decap_4 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_194 ();
 sg13g2_decap_4 FILLER_12_269 ();
 sg13g2_fill_2 FILLER_12_283 ();
 sg13g2_fill_1 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_fill_2 FILLER_13_92 ();
 sg13g2_fill_1 FILLER_13_94 ();
 sg13g2_fill_2 FILLER_13_136 ();
 sg13g2_decap_8 FILLER_13_198 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_decap_4 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_2 FILLER_13_282 ();
 sg13g2_decap_8 FILLER_13_344 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_fill_2 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_4 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_51 ();
 sg13g2_fill_2 FILLER_14_83 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_fill_2 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_108 ();
 sg13g2_decap_4 FILLER_14_117 ();
 sg13g2_fill_2 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_184 ();
 sg13g2_fill_1 FILLER_14_195 ();
 sg13g2_decap_4 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_decap_4 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_fill_1 FILLER_14_275 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_fill_2 FILLER_14_368 ();
 sg13g2_fill_1 FILLER_14_396 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_fill_2 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_decap_4 FILLER_15_124 ();
 sg13g2_fill_2 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_159 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_4 FILLER_15_232 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_4 FILLER_15_341 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_2 FILLER_15_363 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_fill_2 FILLER_15_386 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_fill_2 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_8 FILLER_16_135 ();
 sg13g2_decap_4 FILLER_16_142 ();
 sg13g2_decap_4 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_fill_2 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_43 ();
 sg13g2_fill_1 FILLER_17_50 ();
 sg13g2_decap_4 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_decap_8 FILLER_17_66 ();
 sg13g2_decap_8 FILLER_17_73 ();
 sg13g2_decap_4 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_4 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_4 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_275 ();
 sg13g2_fill_2 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_decap_4 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_157 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_2 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_201 ();
 sg13g2_decap_4 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_212 ();
 sg13g2_decap_4 FILLER_18_228 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_decap_4 FILLER_19_74 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_1 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_fill_1 FILLER_19_130 ();
 sg13g2_fill_2 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_159 ();
 sg13g2_decap_4 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_194 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_4 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_270 ();
 sg13g2_decap_4 FILLER_19_283 ();
 sg13g2_decap_4 FILLER_19_296 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_decap_4 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_375 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_31 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_fill_1 FILLER_20_48 ();
 sg13g2_decap_4 FILLER_20_72 ();
 sg13g2_decap_4 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_95 ();
 sg13g2_fill_1 FILLER_20_97 ();
 sg13g2_fill_2 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_106 ();
 sg13g2_decap_4 FILLER_20_123 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_decap_4 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_157 ();
 sg13g2_fill_1 FILLER_20_159 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_185 ();
 sg13g2_decap_4 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_196 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_298 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_20 ();
 sg13g2_fill_1 FILLER_21_27 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_44 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_decap_8 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_82 ();
 sg13g2_fill_1 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_decap_8 FILLER_21_121 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_fill_2 FILLER_21_163 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_fill_2 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_decap_4 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_4 FILLER_21_388 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_110 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_4 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_decap_4 FILLER_22_278 ();
 sg13g2_fill_1 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_fill_2 FILLER_22_372 ();
 sg13g2_fill_2 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_20 ();
 sg13g2_fill_1 FILLER_23_24 ();
 sg13g2_fill_2 FILLER_23_44 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_100 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_121 ();
 sg13g2_fill_1 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_decap_4 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_decap_4 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_decap_4 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_332 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_58 ();
 sg13g2_decap_4 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_88 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_2 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_142 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_2 FILLER_24_360 ();
 sg13g2_decap_4 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_371 ();
 sg13g2_decap_4 FILLER_24_398 ();
 sg13g2_fill_2 FILLER_24_402 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_33 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_decap_8 FILLER_25_72 ();
 sg13g2_decap_4 FILLER_25_79 ();
 sg13g2_decap_8 FILLER_25_110 ();
 sg13g2_decap_8 FILLER_25_117 ();
 sg13g2_decap_4 FILLER_25_124 ();
 sg13g2_fill_1 FILLER_25_128 ();
 sg13g2_decap_8 FILLER_25_134 ();
 sg13g2_fill_2 FILLER_25_141 ();
 sg13g2_fill_1 FILLER_25_143 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_decap_4 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_decap_4 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_decap_4 FILLER_26_113 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_2 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_decap_4 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_262 ();
 sg13g2_decap_4 FILLER_26_269 ();
 sg13g2_decap_4 FILLER_26_282 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_fill_2 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_320 ();
 sg13g2_decap_4 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_4 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_decap_8 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_decap_4 FILLER_27_104 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_181 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_decap_4 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_4 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_368 ();
 sg13g2_decap_4 FILLER_27_375 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_70 ();
 sg13g2_decap_4 FILLER_28_85 ();
 sg13g2_fill_2 FILLER_28_124 ();
 sg13g2_decap_8 FILLER_28_152 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_decap_8 FILLER_28_166 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_decap_8 FILLER_28_183 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_4 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_274 ();
 sg13g2_decap_4 FILLER_28_281 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_4 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_43 ();
 sg13g2_fill_2 FILLER_29_47 ();
 sg13g2_decap_4 FILLER_29_58 ();
 sg13g2_decap_8 FILLER_29_86 ();
 sg13g2_decap_4 FILLER_29_107 ();
 sg13g2_decap_4 FILLER_29_117 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_fill_2 FILLER_29_279 ();
 sg13g2_decap_4 FILLER_29_290 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_2 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_decap_8 FILLER_30_124 ();
 sg13g2_decap_8 FILLER_30_131 ();
 sg13g2_decap_4 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_1 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_decap_4 FILLER_30_270 ();
 sg13g2_decap_4 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_2 FILLER_30_391 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_55 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_301 ();
 sg13g2_decap_4 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_54 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_fill_2 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_2 FILLER_32_120 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_decap_4 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_decap_4 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_fill_1 FILLER_33_89 ();
 sg13g2_fill_2 FILLER_33_103 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_184 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_decap_8 FILLER_33_209 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_decap_4 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_323 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_decap_4 FILLER_33_342 ();
 sg13g2_decap_4 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_64 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_183 ();
 sg13g2_fill_1 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_58 ();
 sg13g2_fill_1 FILLER_35_82 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_134 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_decap_4 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_decap_8 FILLER_35_297 ();
 sg13g2_decap_4 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_51 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_105 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_decap_8 FILLER_36_211 ();
 sg13g2_decap_4 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_decap_4 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_decap_4 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_fill_1 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_104 ();
 sg13g2_decap_4 FILLER_37_111 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_fill_2 FILLER_37_248 ();
 sg13g2_decap_4 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_394 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_4 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_39 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_223 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_decap_4 FILLER_38_332 ();
 sg13g2_fill_1 FILLER_38_356 ();
 sg13g2_fill_1 FILLER_38_366 ();
 sg13g2_fill_2 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_383 ();
 assign uio_oe[0] = net147;
 assign uio_oe[1] = net148;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net149;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[2] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
 assign uio_out[7] = net15;
 assign uo_out[0] = net16;
 assign uo_out[1] = net17;
 assign uo_out[2] = net18;
 assign uo_out[3] = net19;
 assign uo_out[4] = net20;
 assign uo_out[5] = net21;
 assign uo_out[6] = net22;
 assign uo_out[7] = net23;
endmodule
