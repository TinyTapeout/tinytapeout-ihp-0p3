module tt_um_strau0106_simple_viii (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire clknet_leaf_0_clk;
 wire \cpu_instance.addr_reg_op[0] ;
 wire \cpu_instance.addr_reg_op[1] ;
 wire \cpu_instance.addr_reg_op[2] ;
 wire \cpu_instance.addr_sel ;
 wire \cpu_instance.alu_instance.op[0] ;
 wire \cpu_instance.alu_instance.op[1] ;
 wire \cpu_instance.alu_instance.op[2] ;
 wire \cpu_instance.alu_instance.op[3] ;
 wire \cpu_instance.ctrl_instance.flag_carry ;
 wire \cpu_instance.ctrl_instance.flag_zero ;
 wire \cpu_instance.ctrl_instance.jmp_op_addr_sel ;
 wire \cpu_instance.ctrl_instance.mem_op_done ;
 wire \cpu_instance.ctrl_instance.scan_in ;
 wire \cpu_instance.ctrl_instance.scan_out ;
 wire \cpu_instance.ctrl_instance.state[0] ;
 wire \cpu_instance.ctrl_instance.state[1] ;
 wire \cpu_instance.ctrl_instance.state[2] ;
 wire \cpu_instance.ctrl_instance.state[3] ;
 wire \cpu_instance.ctrl_instance.use_register_bank_in ;
 wire \cpu_instance.ctrl_instance.use_register_bank_out_1 ;
 wire \cpu_instance.mem_ctrl_op[0] ;
 wire \cpu_instance.mem_ctrl_op[1] ;
 wire \cpu_instance.mem_instance.addr[24] ;
 wire \cpu_instance.mem_instance.bus_data_out[0] ;
 wire \cpu_instance.mem_instance.bus_data_out[1] ;
 wire \cpu_instance.mem_instance.bus_data_out[2] ;
 wire \cpu_instance.mem_instance.bus_data_out[3] ;
 wire \cpu_instance.mem_instance.bus_data_out[4] ;
 wire \cpu_instance.mem_instance.bus_data_out[5] ;
 wire \cpu_instance.mem_instance.bus_data_out[6] ;
 wire \cpu_instance.mem_instance.bus_data_out[7] ;
 wire \cpu_instance.mem_instance.data_qi_mo[1] ;
 wire \cpu_instance.mem_instance.data_qi_mo[2] ;
 wire \cpu_instance.mem_instance.data_qi_mo[3] ;
 wire \cpu_instance.mem_instance.data_qi_mo[4] ;
 wire \cpu_instance.mem_instance.data_qi_mo[5] ;
 wire \cpu_instance.mem_instance.data_qi_mo[6] ;
 wire \cpu_instance.mem_instance.data_qi_mo[7] ;
 wire \cpu_instance.mem_instance.data_qo_mi[0] ;
 wire \cpu_instance.mem_instance.data_qo_mi[1] ;
 wire \cpu_instance.mem_instance.data_qo_mi[2] ;
 wire \cpu_instance.mem_instance.data_qo_mi[3] ;
 wire \cpu_instance.mem_instance.data_qo_mi[4] ;
 wire \cpu_instance.mem_instance.data_qo_mi[5] ;
 wire \cpu_instance.mem_instance.data_qo_mi[6] ;
 wire \cpu_instance.mem_instance.data_qo_mi[7] ;
 wire \cpu_instance.mem_instance.data_ready ;
 wire \cpu_instance.mem_instance.data_req ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][10] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][4] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][6] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][7] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][8] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.start_read ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.start_write ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.state[0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.state[1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.stop_txn ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[10] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[11] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[13] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[14] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[15] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[16] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[17] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[18] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[19] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[3] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[4] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[5] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[6] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[7] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[8] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[9] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.is_writing ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.last_ram_a_sel ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[3] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.stop_txn_reg ;
 wire \cpu_instance.mux_instance.sel[0] ;
 wire \cpu_instance.mux_instance.sel[1] ;
 wire \cpu_instance.reg_1_out_sel[0] ;
 wire \cpu_instance.reg_1_out_sel[1] ;
 wire \cpu_instance.reg_2_out_sel[0] ;
 wire \cpu_instance.reg_2_out_sel[1] ;
 wire \cpu_instance.reg_in_sel[0] ;
 wire \cpu_instance.reg_in_sel[1] ;
 wire \cpu_instance.reg_op ;
 wire \cpu_instance.registers_instance.register_bank[10][0] ;
 wire \cpu_instance.registers_instance.register_bank[10][1] ;
 wire \cpu_instance.registers_instance.register_bank[10][2] ;
 wire \cpu_instance.registers_instance.register_bank[10][3] ;
 wire \cpu_instance.registers_instance.register_bank[10][4] ;
 wire \cpu_instance.registers_instance.register_bank[10][5] ;
 wire \cpu_instance.registers_instance.register_bank[10][6] ;
 wire \cpu_instance.registers_instance.register_bank[10][7] ;
 wire \cpu_instance.registers_instance.register_bank[11][0] ;
 wire \cpu_instance.registers_instance.register_bank[11][1] ;
 wire \cpu_instance.registers_instance.register_bank[11][2] ;
 wire \cpu_instance.registers_instance.register_bank[11][3] ;
 wire \cpu_instance.registers_instance.register_bank[11][4] ;
 wire \cpu_instance.registers_instance.register_bank[11][5] ;
 wire \cpu_instance.registers_instance.register_bank[11][6] ;
 wire \cpu_instance.registers_instance.register_bank[11][7] ;
 wire \cpu_instance.registers_instance.register_bank[12][0] ;
 wire \cpu_instance.registers_instance.register_bank[12][1] ;
 wire \cpu_instance.registers_instance.register_bank[12][2] ;
 wire \cpu_instance.registers_instance.register_bank[12][3] ;
 wire \cpu_instance.registers_instance.register_bank[12][4] ;
 wire \cpu_instance.registers_instance.register_bank[12][5] ;
 wire \cpu_instance.registers_instance.register_bank[12][6] ;
 wire \cpu_instance.registers_instance.register_bank[12][7] ;
 wire \cpu_instance.registers_instance.register_bank[13][0] ;
 wire \cpu_instance.registers_instance.register_bank[13][1] ;
 wire \cpu_instance.registers_instance.register_bank[13][2] ;
 wire \cpu_instance.registers_instance.register_bank[13][3] ;
 wire \cpu_instance.registers_instance.register_bank[13][4] ;
 wire \cpu_instance.registers_instance.register_bank[13][5] ;
 wire \cpu_instance.registers_instance.register_bank[13][6] ;
 wire \cpu_instance.registers_instance.register_bank[13][7] ;
 wire \cpu_instance.registers_instance.register_bank[14][0] ;
 wire \cpu_instance.registers_instance.register_bank[14][1] ;
 wire \cpu_instance.registers_instance.register_bank[14][2] ;
 wire \cpu_instance.registers_instance.register_bank[14][3] ;
 wire \cpu_instance.registers_instance.register_bank[14][4] ;
 wire \cpu_instance.registers_instance.register_bank[14][5] ;
 wire \cpu_instance.registers_instance.register_bank[14][6] ;
 wire \cpu_instance.registers_instance.register_bank[14][7] ;
 wire \cpu_instance.registers_instance.register_bank[15][0] ;
 wire \cpu_instance.registers_instance.register_bank[15][1] ;
 wire \cpu_instance.registers_instance.register_bank[15][2] ;
 wire \cpu_instance.registers_instance.register_bank[15][3] ;
 wire \cpu_instance.registers_instance.register_bank[15][4] ;
 wire \cpu_instance.registers_instance.register_bank[15][5] ;
 wire \cpu_instance.registers_instance.register_bank[15][6] ;
 wire \cpu_instance.registers_instance.register_bank[15][7] ;
 wire \cpu_instance.registers_instance.register_bank[8][0] ;
 wire \cpu_instance.registers_instance.register_bank[8][1] ;
 wire \cpu_instance.registers_instance.register_bank[8][2] ;
 wire \cpu_instance.registers_instance.register_bank[8][3] ;
 wire \cpu_instance.registers_instance.register_bank[8][4] ;
 wire \cpu_instance.registers_instance.register_bank[8][5] ;
 wire \cpu_instance.registers_instance.register_bank[8][6] ;
 wire \cpu_instance.registers_instance.register_bank[8][7] ;
 wire \cpu_instance.registers_instance.register_bank[9][0] ;
 wire \cpu_instance.registers_instance.register_bank[9][1] ;
 wire \cpu_instance.registers_instance.register_bank[9][2] ;
 wire \cpu_instance.registers_instance.register_bank[9][3] ;
 wire \cpu_instance.registers_instance.register_bank[9][4] ;
 wire \cpu_instance.registers_instance.register_bank[9][5] ;
 wire \cpu_instance.registers_instance.register_bank[9][6] ;
 wire \cpu_instance.registers_instance.register_bank[9][7] ;
 wire \cpu_instance.registers_instance.registers[0][0] ;
 wire \cpu_instance.registers_instance.registers[0][1] ;
 wire \cpu_instance.registers_instance.registers[0][2] ;
 wire \cpu_instance.registers_instance.registers[0][3] ;
 wire \cpu_instance.registers_instance.registers[0][4] ;
 wire \cpu_instance.registers_instance.registers[0][5] ;
 wire \cpu_instance.registers_instance.registers[0][6] ;
 wire \cpu_instance.registers_instance.registers[0][7] ;
 wire \cpu_instance.registers_instance.registers[1][0] ;
 wire \cpu_instance.registers_instance.registers[1][1] ;
 wire \cpu_instance.registers_instance.registers[1][2] ;
 wire \cpu_instance.registers_instance.registers[1][3] ;
 wire \cpu_instance.registers_instance.registers[1][4] ;
 wire \cpu_instance.registers_instance.registers[1][5] ;
 wire \cpu_instance.registers_instance.registers[1][6] ;
 wire \cpu_instance.registers_instance.registers[1][7] ;
 wire \cpu_instance.registers_instance.registers[2][0] ;
 wire \cpu_instance.registers_instance.registers[2][1] ;
 wire \cpu_instance.registers_instance.registers[2][2] ;
 wire \cpu_instance.registers_instance.registers[2][3] ;
 wire \cpu_instance.registers_instance.registers[2][4] ;
 wire \cpu_instance.registers_instance.registers[2][5] ;
 wire \cpu_instance.registers_instance.registers[2][6] ;
 wire \cpu_instance.registers_instance.registers[2][7] ;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net904;
 wire net905;
 wire net906;

 sg13g2_inv_1 _2479_ (.Y(_1570_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ));
 sg13g2_inv_1 _2480_ (.Y(_1571_),
    .A(net609));
 sg13g2_inv_1 _2481_ (.Y(_1572_),
    .A(net617));
 sg13g2_inv_1 _2482_ (.Y(_1573_),
    .A(\cpu_instance.registers_instance.registers[2][2] ));
 sg13g2_inv_1 _2483_ (.Y(_1574_),
    .A(net579));
 sg13g2_inv_1 _2484_ (.Y(_1575_),
    .A(\cpu_instance.registers_instance.registers[2][0] ));
 sg13g2_inv_1 _2485_ (.Y(_1576_),
    .A(net587));
 sg13g2_inv_1 _2486_ (.Y(_1577_),
    .A(\cpu_instance.registers_instance.registers[1][2] ));
 sg13g2_inv_1 _2487_ (.Y(_1578_),
    .A(net602));
 sg13g2_inv_1 _2488_ (.Y(_1579_),
    .A(net318));
 sg13g2_inv_1 _2489_ (.Y(_1580_),
    .A(net374));
 sg13g2_inv_1 _2490_ (.Y(_1581_),
    .A(net552));
 sg13g2_inv_1 _2491_ (.Y(_1582_),
    .A(net344));
 sg13g2_inv_1 _2492_ (.Y(_1583_),
    .A(net340));
 sg13g2_inv_4 _2493_ (.A(\cpu_instance.mem_instance.addr[24] ),
    .Y(_1584_));
 sg13g2_inv_1 _2494_ (.Y(_1585_),
    .A(net815));
 sg13g2_inv_1 _2495_ (.Y(_1586_),
    .A(net804));
 sg13g2_inv_1 _2496_ (.Y(_1587_),
    .A(net384));
 sg13g2_inv_1 _2497_ (.Y(_1588_),
    .A(net366));
 sg13g2_inv_1 _2498_ (.Y(_1589_),
    .A(net422));
 sg13g2_inv_2 _2499_ (.Y(_1590_),
    .A(net397));
 sg13g2_inv_1 _2500_ (.Y(_1591_),
    .A(net407));
 sg13g2_inv_1 _2501_ (.Y(_1592_),
    .A(\cpu_instance.reg_1_out_sel[1] ));
 sg13g2_inv_1 _2502_ (.Y(_1593_),
    .A(net818));
 sg13g2_inv_1 _2503_ (.Y(_1594_),
    .A(net820));
 sg13g2_inv_2 _2504_ (.Y(_1595_),
    .A(net821));
 sg13g2_inv_1 _2505_ (.Y(_1596_),
    .A(\cpu_instance.ctrl_instance.use_register_bank_out_1 ));
 sg13g2_inv_1 _2506_ (.Y(_1597_),
    .A(net660));
 sg13g2_inv_1 _2507_ (.Y(_1598_),
    .A(net589));
 sg13g2_inv_1 _2508_ (.Y(_1599_),
    .A(\cpu_instance.reg_op ));
 sg13g2_inv_1 _2509_ (.Y(_1600_),
    .A(_0018_));
 sg13g2_inv_1 _2510_ (.Y(_1601_),
    .A(_0021_));
 sg13g2_inv_1 _2511_ (.Y(_1602_),
    .A(_0020_));
 sg13g2_inv_2 _2512_ (.Y(_1603_),
    .A(net841));
 sg13g2_inv_1 _2513_ (.Y(_1604_),
    .A(net321));
 sg13g2_inv_1 _2514_ (.Y(_1605_),
    .A(net874));
 sg13g2_inv_1 _2515_ (.Y(_1606_),
    .A(net324));
 sg13g2_inv_1 _2516_ (.Y(_1607_),
    .A(net356));
 sg13g2_inv_1 _2517_ (.Y(_1608_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.last_ram_a_sel ));
 sg13g2_inv_1 _2518_ (.Y(_1609_),
    .A(net567));
 sg13g2_inv_1 _2519_ (.Y(_1610_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ));
 sg13g2_inv_1 _2520_ (.Y(_1611_),
    .A(\cpu_instance.addr_reg_op[2] ));
 sg13g2_inv_2 _2521_ (.Y(_1612_),
    .A(net904));
 sg13g2_inv_1 _2522_ (.Y(_1613_),
    .A(_0026_));
 sg13g2_inv_1 _2523_ (.Y(_1614_),
    .A(\cpu_instance.mem_instance.data_ready ));
 sg13g2_inv_2 _2524_ (.Y(_1615_),
    .A(\cpu_instance.ctrl_instance.mem_op_done ));
 sg13g2_inv_1 _2525_ (.Y(_1616_),
    .A(_0001_));
 sg13g2_inv_1 _2526_ (.Y(_1617_),
    .A(_0002_));
 sg13g2_inv_1 _2527_ (.Y(_1618_),
    .A(\cpu_instance.reg_2_out_sel[1] ));
 sg13g2_inv_1 _2528_ (.Y(_1619_),
    .A(_0010_));
 sg13g2_inv_1 _2529_ (.Y(_1620_),
    .A(net335));
 sg13g2_inv_1 _2530_ (.Y(_1621_),
    .A(net332));
 sg13g2_inv_1 _2531_ (.Y(_1622_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[8] ));
 sg13g2_inv_1 _2532_ (.Y(_1623_),
    .A(net358));
 sg13g2_inv_1 _2533_ (.Y(_1624_),
    .A(net339));
 sg13g2_inv_1 _2534_ (.Y(_1625_),
    .A(net348));
 sg13g2_inv_1 _2535_ (.Y(_1626_),
    .A(net548));
 sg13g2_and2_2 _2536_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ),
    .B(net896),
    .X(uio_oe[5]));
 sg13g2_and2_1 _2537_ (.A(net806),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ),
    .X(_1627_));
 sg13g2_nand2_2 _2538_ (.Y(_1628_),
    .A(net806),
    .B(net808));
 sg13g2_nor2_2 _2539_ (.A(net807),
    .B(_1628_),
    .Y(_1629_));
 sg13g2_nand2b_2 _2540_ (.Y(_1630_),
    .B(net796),
    .A_N(net807));
 sg13g2_nor2b_1 _2541_ (.A(net807),
    .B_N(net808),
    .Y(_1631_));
 sg13g2_nand2_1 _2542_ (.Y(_1632_),
    .A(net805),
    .B(_1631_));
 sg13g2_nor2b_2 _2543_ (.A(net808),
    .B_N(net807),
    .Y(_1633_));
 sg13g2_nand2b_1 _2544_ (.Y(_1634_),
    .B(_1633_),
    .A_N(net806));
 sg13g2_nand3_1 _2545_ (.B(_1632_),
    .C(_1634_),
    .A(_1630_),
    .Y(_1635_));
 sg13g2_inv_1 _2546_ (.Y(_1636_),
    .A(_1635_));
 sg13g2_nor2_1 _2547_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ),
    .B(_1632_),
    .Y(_1637_));
 sg13g2_nand2_1 _2548_ (.Y(_1638_),
    .A(net801),
    .B(_1637_));
 sg13g2_nand2_1 _2549_ (.Y(_1639_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ),
    .B(net805));
 sg13g2_nor2_2 _2550_ (.A(net808),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_nand2_1 _2551_ (.Y(_1641_),
    .A(_0023_),
    .B(_1633_));
 sg13g2_a22oi_1 _2552_ (.Y(_1642_),
    .B1(_1640_),
    .B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ),
    .A2(_1629_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[4] ));
 sg13g2_a21oi_2 _2553_ (.B1(_1636_),
    .Y(uio_out[1]),
    .A2(_1642_),
    .A1(_1638_));
 sg13g2_a221oi_1 _2554_ (.B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ),
    .C1(_1637_),
    .B1(_1640_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[5] ),
    .Y(_1643_),
    .A2(_1629_));
 sg13g2_nand2_2 _2555_ (.Y(uio_out[2]),
    .A(_1635_),
    .B(_1643_));
 sg13g2_nand3_1 _2556_ (.B(_1635_),
    .C(_1640_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ),
    .Y(_1644_));
 sg13g2_o21ai_1 _2557_ (.B1(_1644_),
    .Y(uio_out[4]),
    .A1(_1626_),
    .A2(_1630_));
 sg13g2_a22oi_1 _2558_ (.Y(_1645_),
    .B1(_1640_),
    .B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ),
    .A2(_1629_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[7] ));
 sg13g2_nand3_1 _2559_ (.B(_1638_),
    .C(_1645_),
    .A(_1635_),
    .Y(uio_out[5]));
 sg13g2_nor2_1 _2560_ (.A(net798),
    .B(net833),
    .Y(\cpu_instance.ctrl_instance.scan_out ));
 sg13g2_nor2_1 _2561_ (.A(_0024_),
    .B(_1641_),
    .Y(_1646_));
 sg13g2_nand2b_2 _2562_ (.Y(_1647_),
    .B(_1640_),
    .A_N(_0024_));
 sg13g2_nor2_1 _2563_ (.A(net807),
    .B(net808),
    .Y(_1648_));
 sg13g2_and2_1 _2564_ (.A(net805),
    .B(_1648_),
    .X(_1649_));
 sg13g2_nand2_2 _2565_ (.Y(_1650_),
    .A(net805),
    .B(_1648_));
 sg13g2_nor2_2 _2566_ (.A(net324),
    .B(net356),
    .Y(_1651_));
 sg13g2_nor2_1 _2567_ (.A(_1650_),
    .B(_1651_),
    .Y(_1652_));
 sg13g2_nand2b_2 _2568_ (.Y(_1653_),
    .B(net790),
    .A_N(_1651_));
 sg13g2_nor2_2 _2569_ (.A(net771),
    .B(net770),
    .Y(_1654_));
 sg13g2_nand2_2 _2570_ (.Y(_1655_),
    .A(_1647_),
    .B(_1653_));
 sg13g2_a22oi_1 _2571_ (.Y(_1656_),
    .B1(_1654_),
    .B2(net316),
    .A2(net771),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ));
 sg13g2_inv_1 _2572_ (.Y(_0027_),
    .A(net317));
 sg13g2_a22oi_1 _2573_ (.Y(_1657_),
    .B1(_1654_),
    .B2(net314),
    .A2(net771),
    .A1(net323));
 sg13g2_inv_1 _2574_ (.Y(_0028_),
    .A(_1657_));
 sg13g2_a22oi_1 _2575_ (.Y(_1658_),
    .B1(_1654_),
    .B2(net310),
    .A2(net772),
    .A1(net320));
 sg13g2_inv_1 _2576_ (.Y(_0029_),
    .A(_1658_));
 sg13g2_a22oi_1 _2577_ (.Y(_1659_),
    .B1(net760),
    .B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[19] ),
    .A2(net771),
    .A1(net312));
 sg13g2_inv_1 _2578_ (.Y(_0030_),
    .A(net313));
 sg13g2_a22oi_1 _2579_ (.Y(_1660_),
    .B1(net760),
    .B2(net336),
    .A2(net771),
    .A1(net316));
 sg13g2_inv_1 _2580_ (.Y(_0031_),
    .A(_1660_));
 sg13g2_a22oi_1 _2581_ (.Y(_1661_),
    .B1(net760),
    .B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ),
    .A2(net771),
    .A1(net314));
 sg13g2_inv_1 _2582_ (.Y(_0032_),
    .A(net315));
 sg13g2_a22oi_1 _2583_ (.Y(_1662_),
    .B1(net760),
    .B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ),
    .A2(net771),
    .A1(net310));
 sg13g2_inv_1 _2584_ (.Y(_0033_),
    .A(net311));
 sg13g2_nor3_2 _2585_ (.A(\cpu_instance.addr_reg_op[1] ),
    .B(_1612_),
    .C(_1613_),
    .Y(_1663_));
 sg13g2_and2_2 _2586_ (.A(\cpu_instance.addr_reg_op[1] ),
    .B(_0026_),
    .X(_1664_));
 sg13g2_nand2_2 _2587_ (.Y(_1665_),
    .A(\cpu_instance.addr_reg_op[1] ),
    .B(_0026_));
 sg13g2_nor3_2 _2588_ (.A(_1611_),
    .B(\cpu_instance.addr_reg_op[1] ),
    .C(\cpu_instance.addr_reg_op[0] ),
    .Y(_1666_));
 sg13g2_nand3b_1 _2589_ (.B(_1612_),
    .C(\cpu_instance.addr_reg_op[2] ),
    .Y(_1667_),
    .A_N(\cpu_instance.addr_reg_op[1] ));
 sg13g2_nand2_2 _2590_ (.Y(_1668_),
    .A(_1665_),
    .B(_1667_));
 sg13g2_nor2_2 _2591_ (.A(_1663_),
    .B(_1668_),
    .Y(_1669_));
 sg13g2_nand2_1 _2592_ (.Y(_1670_),
    .A(net814),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ));
 sg13g2_nand2_2 _2593_ (.Y(_1671_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ),
    .B(net802));
 sg13g2_and2_2 _2594_ (.A(_1670_),
    .B(_1671_),
    .X(_1672_));
 sg13g2_nand2_1 _2595_ (.Y(_1673_),
    .A(_1670_),
    .B(_1671_));
 sg13g2_nor2_2 _2596_ (.A(\cpu_instance.mux_instance.sel[0] ),
    .B(\cpu_instance.mux_instance.sel[1] ),
    .Y(_1674_));
 sg13g2_inv_1 _2597_ (.Y(_1675_),
    .A(_1674_));
 sg13g2_nand2b_2 _2598_ (.Y(_1676_),
    .B(\cpu_instance.alu_instance.op[3] ),
    .A_N(\cpu_instance.alu_instance.op[2] ));
 sg13g2_nor2_1 _2599_ (.A(\cpu_instance.alu_instance.op[1] ),
    .B(\cpu_instance.alu_instance.op[0] ),
    .Y(_1677_));
 sg13g2_nor2b_2 _2600_ (.A(_1676_),
    .B_N(_1677_),
    .Y(_1678_));
 sg13g2_inv_1 _2601_ (.Y(_1679_),
    .A(_1678_));
 sg13g2_nor2_1 _2602_ (.A(net800),
    .B(net818),
    .Y(_1680_));
 sg13g2_nand2_1 _2603_ (.Y(_1681_),
    .A(net816),
    .B(net818));
 sg13g2_nor2_1 _2604_ (.A(net816),
    .B(_1593_),
    .Y(_1682_));
 sg13g2_nor2_2 _2605_ (.A(net816),
    .B(net818),
    .Y(_1683_));
 sg13g2_mux4_1 _2606_ (.S0(net800),
    .A0(_1575_),
    .A1(_0018_),
    .A2(_0001_),
    .A3(_1579_),
    .S1(net817),
    .X(_1684_));
 sg13g2_and2_1 _2607_ (.A(net798),
    .B(net788),
    .X(_1685_));
 sg13g2_mux4_1 _2608_ (.S0(net800),
    .A0(_1574_),
    .A1(_0019_),
    .A2(_0002_),
    .A3(_1578_),
    .S1(net817),
    .X(_1686_));
 sg13g2_mux4_1 _2609_ (.S0(net817),
    .A0(\cpu_instance.registers_instance.registers[0][2] ),
    .A1(\cpu_instance.registers_instance.registers[1][2] ),
    .A2(\cpu_instance.registers_instance.registers[2][2] ),
    .A3(uo_out[2]),
    .S1(net816),
    .X(_1687_));
 sg13g2_mux4_1 _2610_ (.S0(_1593_),
    .A0(_1571_),
    .A1(_1573_),
    .A2(_1577_),
    .A3(_1581_),
    .S1(net800),
    .X(_1688_));
 sg13g2_mux4_1 _2611_ (.S0(net817),
    .A0(\cpu_instance.registers_instance.registers[2][3] ),
    .A1(_1601_),
    .A2(_1602_),
    .A3(\cpu_instance.registers_instance.registers[1][3] ),
    .S1(_1592_),
    .X(_1689_));
 sg13g2_mux4_1 _2612_ (.S0(net817),
    .A0(_1572_),
    .A1(_0021_),
    .A2(_0020_),
    .A3(_1576_),
    .S1(_1592_),
    .X(_1690_));
 sg13g2_nor4_2 _2613_ (.A(net787),
    .B(net785),
    .C(net784),
    .Y(_1691_),
    .D(_1690_));
 sg13g2_mux4_1 _2614_ (.S0(net800),
    .A0(\cpu_instance.registers_instance.registers[2][0] ),
    .A1(\cpu_instance.registers_instance.registers[0][0] ),
    .A2(_1616_),
    .A3(\cpu_instance.registers_instance.registers[1][0] ),
    .S1(net818),
    .X(_1692_));
 sg13g2_nor4_2 _2615_ (.A(net786),
    .B(_1688_),
    .C(_1690_),
    .Y(_1693_),
    .D(net783));
 sg13g2_mux4_1 _2616_ (.S0(net800),
    .A0(\cpu_instance.registers_instance.registers[2][1] ),
    .A1(\cpu_instance.registers_instance.registers[0][1] ),
    .A2(_1617_),
    .A3(\cpu_instance.registers_instance.registers[1][1] ),
    .S1(net817),
    .X(_1694_));
 sg13g2_nor2_1 _2617_ (.A(net787),
    .B(_1694_),
    .Y(_1695_));
 sg13g2_nor4_2 _2618_ (.A(net787),
    .B(net784),
    .C(_1690_),
    .Y(_1696_),
    .D(net782));
 sg13g2_nor4_2 _2619_ (.A(net785),
    .B(net784),
    .C(_1689_),
    .Y(_1697_),
    .D(net783));
 sg13g2_nor4_2 _2620_ (.A(net787),
    .B(_1687_),
    .C(_1690_),
    .Y(_1698_),
    .D(net782));
 sg13g2_nor4_2 _2621_ (.A(net787),
    .B(net785),
    .C(_1687_),
    .Y(_1699_),
    .D(_1690_));
 sg13g2_nor4_2 _2622_ (.A(net788),
    .B(net785),
    .C(net784),
    .Y(_1700_),
    .D(_1689_));
 sg13g2_a21oi_1 _2623_ (.A1(net787),
    .A2(net783),
    .Y(_1701_),
    .B1(net785));
 sg13g2_nor4_2 _2624_ (.A(_1687_),
    .B(_1690_),
    .C(net783),
    .Y(_1702_),
    .D(net782));
 sg13g2_nor4_2 _2625_ (.A(net784),
    .B(_1690_),
    .C(net783),
    .Y(_1703_),
    .D(net782));
 sg13g2_nor4_2 _2626_ (.A(net784),
    .B(_1689_),
    .C(_1692_),
    .Y(_1704_),
    .D(net782));
 sg13g2_nor3_1 _2627_ (.A(net784),
    .B(net783),
    .C(net782),
    .Y(_1705_));
 sg13g2_nor4_1 _2628_ (.A(_1695_),
    .B(_1701_),
    .C(_1702_),
    .D(_1705_),
    .Y(_1706_));
 sg13g2_inv_1 _2629_ (.Y(_1707_),
    .A(net758));
 sg13g2_nor2b_1 _2630_ (.A(_0007_),
    .B_N(net758),
    .Y(_1708_));
 sg13g2_nor4_2 _2631_ (.A(net787),
    .B(_1687_),
    .C(_1689_),
    .Y(_1709_),
    .D(net782));
 sg13g2_a22oi_1 _2632_ (.Y(_1710_),
    .B1(_1709_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .A2(_1703_),
    .A1(\cpu_instance.registers_instance.register_bank[12][0] ));
 sg13g2_nor4_2 _2633_ (.A(net788),
    .B(net785),
    .C(_1687_),
    .Y(_1711_),
    .D(_1689_));
 sg13g2_nor4_2 _2634_ (.A(net787),
    .B(net784),
    .C(_1689_),
    .Y(_1712_),
    .D(net782));
 sg13g2_a22oi_1 _2635_ (.Y(_1713_),
    .B1(_1712_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ),
    .A2(_1711_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ));
 sg13g2_nor4_2 _2636_ (.A(net785),
    .B(_1687_),
    .C(_1689_),
    .Y(_1714_),
    .D(net783));
 sg13g2_nor4_2 _2637_ (.A(net785),
    .B(_1687_),
    .C(_1690_),
    .Y(_1715_),
    .D(net783));
 sg13g2_a22oi_1 _2638_ (.Y(_1716_),
    .B1(net764),
    .B2(\cpu_instance.registers_instance.register_bank[8][0] ),
    .A2(_1698_),
    .A1(\cpu_instance.registers_instance.register_bank[9][0] ));
 sg13g2_a21oi_1 _2639_ (.A1(\cpu_instance.registers_instance.register_bank[11][0] ),
    .A2(_1699_),
    .Y(_1717_),
    .B1(net799));
 sg13g2_a22oi_1 _2640_ (.Y(_1718_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][0] ),
    .A2(_1704_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ));
 sg13g2_nand4_1 _2641_ (.B(_1716_),
    .C(_1717_),
    .A(_1710_),
    .Y(_1719_),
    .D(_1718_));
 sg13g2_a22oi_1 _2642_ (.Y(_1720_),
    .B1(_1696_),
    .B2(\cpu_instance.registers_instance.register_bank[13][0] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][0] ));
 sg13g2_a22oi_1 _2643_ (.Y(_1721_),
    .B1(_1700_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ),
    .A2(_1697_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ));
 sg13g2_a22oi_1 _2644_ (.Y(_1722_),
    .B1(_1714_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ),
    .A2(_1693_),
    .A1(\cpu_instance.registers_instance.register_bank[14][0] ));
 sg13g2_nand4_1 _2645_ (.B(_1720_),
    .C(_1721_),
    .A(_1713_),
    .Y(_1723_),
    .D(_1722_));
 sg13g2_nor3_2 _2646_ (.A(_1708_),
    .B(_1719_),
    .C(_1723_),
    .Y(_1724_));
 sg13g2_nor2_2 _2647_ (.A(_1685_),
    .B(_1724_),
    .Y(_1725_));
 sg13g2_or2_1 _2648_ (.X(_1726_),
    .B(_1724_),
    .A(_1685_));
 sg13g2_nor2_1 _2649_ (.A(\cpu_instance.reg_2_out_sel[0] ),
    .B(\cpu_instance.reg_2_out_sel[1] ),
    .Y(_1727_));
 sg13g2_and2_2 _2650_ (.A(\cpu_instance.reg_2_out_sel[0] ),
    .B(\cpu_instance.reg_2_out_sel[1] ),
    .X(_1728_));
 sg13g2_nor2_2 _2651_ (.A(\cpu_instance.reg_2_out_sel[0] ),
    .B(net797),
    .Y(_1729_));
 sg13g2_mux4_1 _2652_ (.S0(net797),
    .A0(\cpu_instance.registers_instance.registers[2][0] ),
    .A1(_1600_),
    .A2(_1616_),
    .A3(\cpu_instance.registers_instance.registers[1][0] ),
    .S1(\cpu_instance.reg_2_out_sel[0] ),
    .X(_1730_));
 sg13g2_inv_1 _2653_ (.Y(_1731_),
    .A(_1730_));
 sg13g2_nor3_2 _2654_ (.A(_1685_),
    .B(_1724_),
    .C(_1731_),
    .Y(_1732_));
 sg13g2_nand2b_2 _2655_ (.Y(_1733_),
    .B(\cpu_instance.alu_instance.op[1] ),
    .A_N(\cpu_instance.alu_instance.op[0] ));
 sg13g2_nor2_2 _2656_ (.A(\cpu_instance.alu_instance.op[3] ),
    .B(\cpu_instance.alu_instance.op[2] ),
    .Y(_1734_));
 sg13g2_nor2b_2 _2657_ (.A(_1733_),
    .B_N(_1734_),
    .Y(_1735_));
 sg13g2_nand2b_1 _2658_ (.Y(_1736_),
    .B(_1734_),
    .A_N(_1733_));
 sg13g2_nand2b_2 _2659_ (.Y(_1737_),
    .B(\cpu_instance.alu_instance.op[0] ),
    .A_N(\cpu_instance.alu_instance.op[1] ));
 sg13g2_nor2_1 _2660_ (.A(\cpu_instance.alu_instance.op[2] ),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_nor2_1 _2661_ (.A(_1735_),
    .B(_1738_),
    .Y(_1739_));
 sg13g2_o21ai_1 _2662_ (.B1(_1679_),
    .Y(_1740_),
    .A1(_1732_),
    .A2(_1739_));
 sg13g2_o21ai_1 _2663_ (.B1(_1740_),
    .Y(_1741_),
    .A1(_1725_),
    .A2(_1730_));
 sg13g2_nor2_2 _2664_ (.A(_1676_),
    .B(_1733_),
    .Y(_1742_));
 sg13g2_or2_1 _2665_ (.X(_1743_),
    .B(_1733_),
    .A(_1676_));
 sg13g2_nand2_1 _2666_ (.Y(_1744_),
    .A(_1726_),
    .B(_1742_));
 sg13g2_and2_2 _2667_ (.A(_1677_),
    .B(_1734_),
    .X(_1745_));
 sg13g2_nand2_1 _2668_ (.Y(_1746_),
    .A(_1677_),
    .B(_1734_));
 sg13g2_and2_1 _2669_ (.A(net798),
    .B(net786),
    .X(_1747_));
 sg13g2_nand2_1 _2670_ (.Y(_1748_),
    .A(net798),
    .B(net786));
 sg13g2_a22oi_1 _2671_ (.Y(_1749_),
    .B1(_1711_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ),
    .A2(_1696_),
    .A1(\cpu_instance.registers_instance.register_bank[13][1] ));
 sg13g2_nor2b_1 _2672_ (.A(_0006_),
    .B_N(net758),
    .Y(_1750_));
 sg13g2_a22oi_1 _2673_ (.Y(_1751_),
    .B1(_1712_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ),
    .A2(_1704_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ));
 sg13g2_a22oi_1 _2674_ (.Y(_1752_),
    .B1(net764),
    .B2(\cpu_instance.registers_instance.register_bank[8][1] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][1] ));
 sg13g2_a22oi_1 _2675_ (.Y(_1753_),
    .B1(_1709_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .A2(_1700_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ));
 sg13g2_a22oi_1 _2676_ (.Y(_1754_),
    .B1(_1714_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ),
    .A2(_1693_),
    .A1(\cpu_instance.registers_instance.register_bank[14][1] ));
 sg13g2_a21oi_1 _2677_ (.A1(\cpu_instance.registers_instance.register_bank[9][1] ),
    .A2(_1698_),
    .Y(_1755_),
    .B1(net799));
 sg13g2_nand4_1 _2678_ (.B(_1752_),
    .C(_1754_),
    .A(_1749_),
    .Y(_1756_),
    .D(_1755_));
 sg13g2_a22oi_1 _2679_ (.Y(_1757_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][1] ),
    .A2(_1703_),
    .A1(\cpu_instance.registers_instance.register_bank[12][1] ));
 sg13g2_a22oi_1 _2680_ (.Y(_1758_),
    .B1(_1699_),
    .B2(\cpu_instance.registers_instance.register_bank[11][1] ),
    .A2(_1697_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ));
 sg13g2_nand4_1 _2681_ (.B(_1753_),
    .C(_1757_),
    .A(_1751_),
    .Y(_1759_),
    .D(_1758_));
 sg13g2_nor3_2 _2682_ (.A(_1750_),
    .B(_1756_),
    .C(_1759_),
    .Y(_1760_));
 sg13g2_or3_1 _2683_ (.A(_1750_),
    .B(_1756_),
    .C(_1759_),
    .X(_1761_));
 sg13g2_nor2_2 _2684_ (.A(_1747_),
    .B(_1760_),
    .Y(_1762_));
 sg13g2_nor2b_1 _2685_ (.A(\cpu_instance.alu_instance.op[3] ),
    .B_N(\cpu_instance.alu_instance.op[2] ),
    .Y(_1763_));
 sg13g2_nand2b_1 _2686_ (.Y(_1764_),
    .B(\cpu_instance.alu_instance.op[2] ),
    .A_N(\cpu_instance.alu_instance.op[3] ));
 sg13g2_nor2_1 _2687_ (.A(_1733_),
    .B(_1764_),
    .Y(_1765_));
 sg13g2_nor2_1 _2688_ (.A(_1737_),
    .B(_1764_),
    .Y(_1766_));
 sg13g2_a21oi_2 _2689_ (.B1(_1764_),
    .Y(_1767_),
    .A2(_1737_),
    .A1(_1733_));
 sg13g2_a22oi_1 _2690_ (.Y(_1768_),
    .B1(_1762_),
    .B2(_1767_),
    .A2(_1745_),
    .A1(_1725_));
 sg13g2_nand3_1 _2691_ (.B(\cpu_instance.alu_instance.op[0] ),
    .C(_1763_),
    .A(\cpu_instance.alu_instance.op[1] ),
    .Y(_1769_));
 sg13g2_inv_2 _2692_ (.Y(_1770_),
    .A(_1769_));
 sg13g2_a22oi_1 _2693_ (.Y(_1771_),
    .B1(_1714_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ),
    .A2(_1709_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ));
 sg13g2_nand2_1 _2694_ (.Y(_1772_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ),
    .B(_1700_));
 sg13g2_a22oi_1 _2695_ (.Y(_1773_),
    .B1(_1696_),
    .B2(\cpu_instance.registers_instance.register_bank[13][7] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][7] ));
 sg13g2_a22oi_1 _2696_ (.Y(_1774_),
    .B1(_1698_),
    .B2(\cpu_instance.registers_instance.register_bank[9][7] ),
    .A2(_1693_),
    .A1(\cpu_instance.registers_instance.register_bank[14][7] ));
 sg13g2_a22oi_1 _2697_ (.Y(_1775_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][7] ),
    .A2(_1699_),
    .A1(\cpu_instance.registers_instance.register_bank[11][7] ));
 sg13g2_a22oi_1 _2698_ (.Y(_1776_),
    .B1(_1703_),
    .B2(\cpu_instance.registers_instance.register_bank[12][7] ),
    .A2(net764),
    .A1(\cpu_instance.registers_instance.register_bank[8][7] ));
 sg13g2_nand4_1 _2699_ (.B(_1774_),
    .C(_1775_),
    .A(_1771_),
    .Y(_1777_),
    .D(_1776_));
 sg13g2_a22oi_1 _2700_ (.Y(_1778_),
    .B1(_1711_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ),
    .A2(_1704_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ));
 sg13g2_a22oi_1 _2701_ (.Y(_1779_),
    .B1(_1712_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ),
    .A2(_1697_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ));
 sg13g2_nand4_1 _2702_ (.B(_1773_),
    .C(_1778_),
    .A(_1772_),
    .Y(_1780_),
    .D(_1779_));
 sg13g2_nor3_2 _2703_ (.A(net757),
    .B(_1777_),
    .C(_1780_),
    .Y(_1781_));
 sg13g2_a21o_1 _2704_ (.A2(net758),
    .A1(_0014_),
    .B1(net798),
    .X(_1782_));
 sg13g2_a221oi_1 _2705_ (.B2(\cpu_instance.registers_instance.registers[2][7] ),
    .C1(_1683_),
    .B1(_1680_),
    .A1(\cpu_instance.registers_instance.registers[1][7] ),
    .Y(_1783_),
    .A2(net800));
 sg13g2_o21ai_1 _2706_ (.B1(_1783_),
    .Y(_1784_),
    .A1(_0013_),
    .A2(_1681_));
 sg13g2_a21oi_1 _2707_ (.A1(_0012_),
    .A2(_1683_),
    .Y(_1785_),
    .B1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ));
 sg13g2_nand2_2 _2708_ (.Y(_1786_),
    .A(_1784_),
    .B(_1785_));
 sg13g2_o21ai_1 _2709_ (.B1(_1786_),
    .Y(_1787_),
    .A1(_1781_),
    .A2(_1782_));
 sg13g2_nand2_1 _2710_ (.Y(_1788_),
    .A(_1677_),
    .B(_1763_));
 sg13g2_inv_1 _2711_ (.Y(_1789_),
    .A(_1788_));
 sg13g2_a22oi_1 _2712_ (.Y(_1790_),
    .B1(_1787_),
    .B2(_1789_),
    .A2(_1770_),
    .A1(_1732_));
 sg13g2_nand4_1 _2713_ (.B(_1744_),
    .C(_1768_),
    .A(_1741_),
    .Y(_1791_),
    .D(_1790_));
 sg13g2_nor2b_2 _2714_ (.A(\cpu_instance.mux_instance.sel[1] ),
    .B_N(\cpu_instance.mux_instance.sel[0] ),
    .Y(_1792_));
 sg13g2_a22oi_1 _2715_ (.Y(_1793_),
    .B1(_1792_),
    .B2(\cpu_instance.mem_instance.bus_data_out[0] ),
    .A2(_1791_),
    .A1(_1674_));
 sg13g2_nor2_1 _2716_ (.A(_1672_),
    .B(net717),
    .Y(_1794_));
 sg13g2_xnor2_1 _2717_ (.Y(_1795_),
    .A(net767),
    .B(net718));
 sg13g2_o21ai_1 _2718_ (.B1(_1667_),
    .Y(_1796_),
    .A1(net814),
    .A2(_1665_));
 sg13g2_a22oi_1 _2719_ (.Y(_1797_),
    .B1(_1796_),
    .B2(_1670_),
    .A2(_1795_),
    .A1(_1664_));
 sg13g2_a21oi_1 _2720_ (.A1(net802),
    .A2(_0017_),
    .Y(_1798_),
    .B1(_1797_));
 sg13g2_o21ai_1 _2721_ (.B1(_1663_),
    .Y(_1799_),
    .A1(net814),
    .A2(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ));
 sg13g2_a21oi_1 _2722_ (.A1(net814),
    .A2(net718),
    .Y(_1800_),
    .B1(_1799_));
 sg13g2_and2_1 _2723_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ),
    .B(_1669_),
    .X(_1801_));
 sg13g2_or3_2 _2724_ (.A(_1798_),
    .B(_1800_),
    .C(_1801_),
    .X(_1802_));
 sg13g2_o21ai_1 _2725_ (.B1(net876),
    .Y(_1803_),
    .A1(net842),
    .A2(_1802_));
 sg13g2_a21oi_1 _2726_ (.A1(_1590_),
    .A2(net842),
    .Y(_0034_),
    .B1(_1803_));
 sg13g2_o21ai_1 _2727_ (.B1(net905),
    .Y(_1804_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .A2(net801));
 sg13g2_nand3b_1 _2728_ (.B(net896),
    .C(_1804_),
    .Y(_1805_),
    .A_N(net671));
 sg13g2_nor2_1 _2729_ (.A(_1604_),
    .B(net762),
    .Y(_0035_));
 sg13g2_nand2b_1 _2730_ (.Y(_1806_),
    .B(_1728_),
    .A_N(_0013_));
 sg13g2_a221oi_1 _2731_ (.B2(\cpu_instance.registers_instance.registers[2][7] ),
    .C1(net794),
    .B1(_1729_),
    .A1(\cpu_instance.registers_instance.registers[1][7] ),
    .Y(_1807_),
    .A2(net797));
 sg13g2_a22oi_1 _2732_ (.Y(_1808_),
    .B1(_1806_),
    .B2(_1807_),
    .A2(net794),
    .A1(_0012_));
 sg13g2_inv_1 _2733_ (.Y(_1809_),
    .A(_1808_));
 sg13g2_nand2b_1 _2734_ (.Y(_1810_),
    .B(_1809_),
    .A_N(_1787_));
 sg13g2_nand2_1 _2735_ (.Y(_1811_),
    .A(_1787_),
    .B(_1808_));
 sg13g2_and2_1 _2736_ (.A(_1810_),
    .B(_1811_),
    .X(_1812_));
 sg13g2_nand2_1 _2737_ (.Y(_1813_),
    .A(_1810_),
    .B(_1811_));
 sg13g2_nand2_1 _2738_ (.Y(_1814_),
    .A(\cpu_instance.registers_instance.register_bank[12][6] ),
    .B(_1703_));
 sg13g2_a22oi_1 _2739_ (.Y(_1815_),
    .B1(_1700_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ),
    .A2(_1698_),
    .A1(\cpu_instance.registers_instance.register_bank[9][6] ));
 sg13g2_a22oi_1 _2740_ (.Y(_1816_),
    .B1(_1712_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ),
    .A2(_1699_),
    .A1(\cpu_instance.registers_instance.register_bank[11][6] ));
 sg13g2_a22oi_1 _2741_ (.Y(_1817_),
    .B1(_1697_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ),
    .A2(_1696_),
    .A1(\cpu_instance.registers_instance.register_bank[13][6] ));
 sg13g2_a22oi_1 _2742_ (.Y(_1818_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][6] ),
    .A2(_1714_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ));
 sg13g2_nand4_1 _2743_ (.B(_1816_),
    .C(_1817_),
    .A(_1815_),
    .Y(_1819_),
    .D(_1818_));
 sg13g2_a22oi_1 _2744_ (.Y(_1820_),
    .B1(_1709_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ),
    .A2(net764),
    .A1(\cpu_instance.registers_instance.register_bank[8][6] ));
 sg13g2_a22oi_1 _2745_ (.Y(_1821_),
    .B1(_1711_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ),
    .A2(_1693_),
    .A1(\cpu_instance.registers_instance.register_bank[14][6] ));
 sg13g2_a22oi_1 _2746_ (.Y(_1822_),
    .B1(_1704_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][6] ));
 sg13g2_nand4_1 _2747_ (.B(_1820_),
    .C(_1821_),
    .A(_1814_),
    .Y(_1823_),
    .D(_1822_));
 sg13g2_or3_2 _2748_ (.A(net757),
    .B(_1819_),
    .C(_1823_),
    .X(_1824_));
 sg13g2_a21oi_2 _2749_ (.B1(net798),
    .Y(_1825_),
    .A2(net757),
    .A1(_0011_));
 sg13g2_a221oi_1 _2750_ (.B2(\cpu_instance.registers_instance.registers[2][6] ),
    .C1(_1683_),
    .B1(_1680_),
    .A1(\cpu_instance.registers_instance.registers[1][6] ),
    .Y(_1826_),
    .A2(net800));
 sg13g2_o21ai_1 _2751_ (.B1(_1826_),
    .Y(_1827_),
    .A1(_0010_),
    .A2(_1681_));
 sg13g2_a21oi_1 _2752_ (.A1(_0009_),
    .A2(_1683_),
    .Y(_1828_),
    .B1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ));
 sg13g2_a22oi_1 _2753_ (.Y(_1829_),
    .B1(_1827_),
    .B2(_1828_),
    .A2(_1825_),
    .A1(_1824_));
 sg13g2_inv_1 _2754_ (.Y(_1830_),
    .A(_1829_));
 sg13g2_a21oi_1 _2755_ (.A1(\cpu_instance.registers_instance.registers[1][6] ),
    .A2(net797),
    .Y(_1831_),
    .B1(net794));
 sg13g2_a22oi_1 _2756_ (.Y(_1832_),
    .B1(_1729_),
    .B2(\cpu_instance.registers_instance.registers[2][6] ),
    .A2(_1728_),
    .A1(_1619_));
 sg13g2_a22oi_1 _2757_ (.Y(_1833_),
    .B1(_1831_),
    .B2(_1832_),
    .A2(net794),
    .A1(_0009_));
 sg13g2_nand2b_1 _2758_ (.Y(_1834_),
    .B(_1833_),
    .A_N(_1829_));
 sg13g2_inv_1 _2759_ (.Y(_1835_),
    .A(_1834_));
 sg13g2_nand2b_2 _2760_ (.Y(_1836_),
    .B(_1829_),
    .A_N(_1833_));
 sg13g2_nand2_1 _2761_ (.Y(_1837_),
    .A(_1834_),
    .B(_1836_));
 sg13g2_a22oi_1 _2762_ (.Y(_1838_),
    .B1(_1711_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][5] ));
 sg13g2_nand2_1 _2763_ (.Y(_1839_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ),
    .B(_1700_));
 sg13g2_a22oi_1 _2764_ (.Y(_1840_),
    .B1(_1698_),
    .B2(\cpu_instance.registers_instance.register_bank[9][5] ),
    .A2(_1697_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ));
 sg13g2_nand2_1 _2765_ (.Y(_1841_),
    .A(_1839_),
    .B(_1840_));
 sg13g2_a22oi_1 _2766_ (.Y(_1842_),
    .B1(_1712_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ),
    .A2(net764),
    .A1(\cpu_instance.registers_instance.register_bank[8][5] ));
 sg13g2_a22oi_1 _2767_ (.Y(_1843_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][5] ),
    .A2(_1699_),
    .A1(\cpu_instance.registers_instance.register_bank[11][5] ));
 sg13g2_nand3b_1 _2768_ (.B(_1842_),
    .C(_1843_),
    .Y(_1844_),
    .A_N(net757));
 sg13g2_a22oi_1 _2769_ (.Y(_1845_),
    .B1(_1709_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .A2(_1703_),
    .A1(\cpu_instance.registers_instance.register_bank[12][5] ));
 sg13g2_a22oi_1 _2770_ (.Y(_1846_),
    .B1(_1696_),
    .B2(\cpu_instance.registers_instance.register_bank[13][5] ),
    .A2(_1693_),
    .A1(\cpu_instance.registers_instance.register_bank[14][5] ));
 sg13g2_a22oi_1 _2771_ (.Y(_1847_),
    .B1(_1714_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ),
    .A2(_1704_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ));
 sg13g2_nand4_1 _2772_ (.B(_1845_),
    .C(_1846_),
    .A(_1838_),
    .Y(_1848_),
    .D(_1847_));
 sg13g2_nor3_2 _2773_ (.A(_1841_),
    .B(_1844_),
    .C(_1848_),
    .Y(_1849_));
 sg13g2_o21ai_1 _2774_ (.B1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .Y(_1850_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .A2(_1707_));
 sg13g2_nand3_1 _2775_ (.B(net816),
    .C(net817),
    .A(uo_out[5]),
    .Y(_1851_));
 sg13g2_a221oi_1 _2776_ (.B2(\cpu_instance.registers_instance.registers[1][5] ),
    .C1(_1683_),
    .B1(_1682_),
    .A1(\cpu_instance.registers_instance.registers[2][5] ),
    .Y(_1852_),
    .A2(_1593_));
 sg13g2_a221oi_1 _2777_ (.B2(_1852_),
    .C1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .B1(_1851_),
    .A1(_1580_),
    .Y(_1853_),
    .A2(_1683_));
 sg13g2_inv_1 _2778_ (.Y(_1854_),
    .A(_1853_));
 sg13g2_o21ai_1 _2779_ (.B1(_1854_),
    .Y(_1855_),
    .A1(_1849_),
    .A2(_1850_));
 sg13g2_inv_1 _2780_ (.Y(_1856_),
    .A(_1855_));
 sg13g2_a21oi_1 _2781_ (.A1(\cpu_instance.registers_instance.registers[1][5] ),
    .A2(net797),
    .Y(_1857_),
    .B1(net794));
 sg13g2_a22oi_1 _2782_ (.Y(_1858_),
    .B1(_1729_),
    .B2(\cpu_instance.registers_instance.registers[2][5] ),
    .A2(_1728_),
    .A1(uo_out[5]));
 sg13g2_a22oi_1 _2783_ (.Y(_1859_),
    .B1(_1857_),
    .B2(_1858_),
    .A2(net794),
    .A1(_0008_));
 sg13g2_inv_1 _2784_ (.Y(_1860_),
    .A(_1859_));
 sg13g2_nor2_1 _2785_ (.A(_1855_),
    .B(_1860_),
    .Y(_1861_));
 sg13g2_nand2_1 _2786_ (.Y(_1862_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .B(_1709_));
 sg13g2_a22oi_1 _2787_ (.Y(_1863_),
    .B1(_1703_),
    .B2(\cpu_instance.registers_instance.register_bank[12][4] ),
    .A2(_1698_),
    .A1(\cpu_instance.registers_instance.register_bank[9][4] ));
 sg13g2_a22oi_1 _2788_ (.Y(_1864_),
    .B1(net764),
    .B2(\cpu_instance.registers_instance.register_bank[8][4] ),
    .A2(_1693_),
    .A1(\cpu_instance.registers_instance.register_bank[14][4] ));
 sg13g2_a22oi_1 _2789_ (.Y(_1865_),
    .B1(_1712_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ),
    .A2(_1696_),
    .A1(\cpu_instance.registers_instance.register_bank[13][4] ));
 sg13g2_a22oi_1 _2790_ (.Y(_1866_),
    .B1(_1699_),
    .B2(\cpu_instance.registers_instance.register_bank[11][4] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][4] ));
 sg13g2_nand4_1 _2791_ (.B(_1864_),
    .C(_1865_),
    .A(_1863_),
    .Y(_1867_),
    .D(_1866_));
 sg13g2_a22oi_1 _2792_ (.Y(_1868_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][4] ),
    .A2(_1697_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ));
 sg13g2_a22oi_1 _2793_ (.Y(_1869_),
    .B1(_1711_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ),
    .A2(_1700_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ));
 sg13g2_a22oi_1 _2794_ (.Y(_1870_),
    .B1(_1714_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ),
    .A2(_1704_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ));
 sg13g2_nand4_1 _2795_ (.B(_1868_),
    .C(_1869_),
    .A(_1862_),
    .Y(_1871_),
    .D(_1870_));
 sg13g2_nor3_2 _2796_ (.A(net757),
    .B(_1867_),
    .C(_1871_),
    .Y(_1872_));
 sg13g2_o21ai_1 _2797_ (.B1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .Y(_1873_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .A2(_1707_));
 sg13g2_mux4_1 _2798_ (.S0(net817),
    .A0(\cpu_instance.registers_instance.registers[0][4] ),
    .A1(\cpu_instance.registers_instance.registers[1][4] ),
    .A2(\cpu_instance.registers_instance.registers[2][4] ),
    .A3(uo_out[4]),
    .S1(net816),
    .X(_1874_));
 sg13g2_nand2_1 _2799_ (.Y(_1875_),
    .A(net798),
    .B(_1874_));
 sg13g2_o21ai_1 _2800_ (.B1(_1875_),
    .Y(_1876_),
    .A1(_1872_),
    .A2(_1873_));
 sg13g2_nand2_1 _2801_ (.Y(_1877_),
    .A(\cpu_instance.registers_instance.registers[2][4] ),
    .B(_1729_));
 sg13g2_a221oi_1 _2802_ (.B2(uo_out[4]),
    .C1(net794),
    .B1(_1728_),
    .A1(\cpu_instance.registers_instance.registers[1][4] ),
    .Y(_1878_),
    .A2(net797));
 sg13g2_a22oi_1 _2803_ (.Y(_1879_),
    .B1(_1877_),
    .B2(_1878_),
    .A2(net794),
    .A1(_0003_));
 sg13g2_inv_1 _2804_ (.Y(_1880_),
    .A(_1879_));
 sg13g2_nand2_2 _2805_ (.Y(_1881_),
    .A(_1876_),
    .B(_1879_));
 sg13g2_nand2b_1 _2806_ (.Y(_1882_),
    .B(_1880_),
    .A_N(_1876_));
 sg13g2_and2_1 _2807_ (.A(_1881_),
    .B(_1882_),
    .X(_1883_));
 sg13g2_nand2_1 _2808_ (.Y(_1884_),
    .A(_1881_),
    .B(_1882_));
 sg13g2_nand2_1 _2809_ (.Y(_1885_),
    .A(\cpu_instance.registers_instance.register_bank[12][3] ),
    .B(_1703_));
 sg13g2_a22oi_1 _2810_ (.Y(_1886_),
    .B1(_1714_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ),
    .A2(_1693_),
    .A1(\cpu_instance.registers_instance.register_bank[14][3] ));
 sg13g2_nand2_1 _2811_ (.Y(_1887_),
    .A(_1885_),
    .B(_1886_));
 sg13g2_a22oi_1 _2812_ (.Y(_1888_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][3] ),
    .A2(_1712_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ));
 sg13g2_a22oi_1 _2813_ (.Y(_1889_),
    .B1(_1704_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ),
    .A2(_1697_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ));
 sg13g2_a22oi_1 _2814_ (.Y(_1890_),
    .B1(_1711_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ),
    .A2(_1709_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ));
 sg13g2_a22oi_1 _2815_ (.Y(_1891_),
    .B1(net764),
    .B2(\cpu_instance.registers_instance.register_bank[8][3] ),
    .A2(_1696_),
    .A1(\cpu_instance.registers_instance.register_bank[13][3] ));
 sg13g2_nand4_1 _2816_ (.B(_1889_),
    .C(_1890_),
    .A(_1888_),
    .Y(_1892_),
    .D(_1891_));
 sg13g2_a22oi_1 _2817_ (.Y(_1893_),
    .B1(_1699_),
    .B2(\cpu_instance.registers_instance.register_bank[11][3] ),
    .A2(_1698_),
    .A1(\cpu_instance.registers_instance.register_bank[9][3] ));
 sg13g2_a22oi_1 _2818_ (.Y(_1894_),
    .B1(_1700_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][3] ));
 sg13g2_nand2_1 _2819_ (.Y(_1895_),
    .A(_1893_),
    .B(_1894_));
 sg13g2_nor4_2 _2820_ (.A(net757),
    .B(_1887_),
    .C(_1892_),
    .Y(_1896_),
    .D(_1895_));
 sg13g2_o21ai_1 _2821_ (.B1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .Y(_1897_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .A2(_1707_));
 sg13g2_nand2_1 _2822_ (.Y(_1898_),
    .A(net799),
    .B(_1689_));
 sg13g2_o21ai_1 _2823_ (.B1(_1898_),
    .Y(_1899_),
    .A1(_1896_),
    .A2(_1897_));
 sg13g2_mux4_1 _2824_ (.S0(\cpu_instance.reg_2_out_sel[0] ),
    .A0(_1572_),
    .A1(_0021_),
    .A2(_0020_),
    .A3(_1576_),
    .S1(_1618_),
    .X(_1900_));
 sg13g2_inv_1 _2825_ (.Y(_1901_),
    .A(_1900_));
 sg13g2_and2_1 _2826_ (.A(net725),
    .B(_1900_),
    .X(_1902_));
 sg13g2_nand2b_1 _2827_ (.Y(_1903_),
    .B(_1900_),
    .A_N(net725));
 sg13g2_xnor2_1 _2828_ (.Y(_1904_),
    .A(net725),
    .B(_1900_));
 sg13g2_xnor2_1 _2829_ (.Y(_1905_),
    .A(net725),
    .B(_1901_));
 sg13g2_mux4_1 _2830_ (.S0(net797),
    .A0(_1574_),
    .A1(_0019_),
    .A2(_0002_),
    .A3(_1578_),
    .S1(\cpu_instance.reg_2_out_sel[0] ),
    .X(_1906_));
 sg13g2_inv_1 _2831_ (.Y(_1907_),
    .A(_1906_));
 sg13g2_nor3_2 _2832_ (.A(_1747_),
    .B(_1760_),
    .C(_1906_),
    .Y(_1908_));
 sg13g2_nand3_1 _2833_ (.B(_1761_),
    .C(_1907_),
    .A(_1748_),
    .Y(_1909_));
 sg13g2_a21oi_2 _2834_ (.B1(_1907_),
    .Y(_1910_),
    .A2(_1761_),
    .A1(_1748_));
 sg13g2_o21ai_1 _2835_ (.B1(_1906_),
    .Y(_0325_),
    .A1(_1747_),
    .A2(_1760_));
 sg13g2_o21ai_1 _2836_ (.B1(_1730_),
    .Y(_0326_),
    .A1(_1685_),
    .A2(_1724_));
 sg13g2_a22oi_1 _2837_ (.Y(_0327_),
    .B1(_1909_),
    .B2(_0325_),
    .A2(_1730_),
    .A1(_1726_));
 sg13g2_o21ai_1 _2838_ (.B1(_0326_),
    .Y(_0328_),
    .A1(_1908_),
    .A2(_1910_));
 sg13g2_nor3_1 _2839_ (.A(_1747_),
    .B(_1760_),
    .C(_1907_),
    .Y(_0329_));
 sg13g2_nand2_1 _2840_ (.Y(_0330_),
    .A(_1762_),
    .B(_1906_));
 sg13g2_nand2_1 _2841_ (.Y(_0331_),
    .A(net798),
    .B(_1687_));
 sg13g2_a22oi_1 _2842_ (.Y(_0332_),
    .B1(_1709_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ),
    .A2(_1700_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ));
 sg13g2_nand2_1 _2843_ (.Y(_0333_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ),
    .B(_1714_));
 sg13g2_a22oi_1 _2844_ (.Y(_0334_),
    .B1(_1693_),
    .B2(\cpu_instance.registers_instance.register_bank[14][2] ),
    .A2(_1691_),
    .A1(\cpu_instance.registers_instance.register_bank[15][2] ));
 sg13g2_a22oi_1 _2845_ (.Y(_0335_),
    .B1(_1712_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ),
    .A2(_1696_),
    .A1(\cpu_instance.registers_instance.register_bank[13][2] ));
 sg13g2_a22oi_1 _2846_ (.Y(_0336_),
    .B1(_1715_),
    .B2(\cpu_instance.registers_instance.register_bank[10][2] ),
    .A2(_1698_),
    .A1(\cpu_instance.registers_instance.register_bank[9][2] ));
 sg13g2_nand4_1 _2847_ (.B(_0334_),
    .C(_0335_),
    .A(_0332_),
    .Y(_0337_),
    .D(_0336_));
 sg13g2_a22oi_1 _2848_ (.Y(_0338_),
    .B1(_1711_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ),
    .A2(_1703_),
    .A1(\cpu_instance.registers_instance.register_bank[12][2] ));
 sg13g2_a22oi_1 _2849_ (.Y(_0339_),
    .B1(_1704_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ),
    .A2(_1697_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ));
 sg13g2_a22oi_1 _2850_ (.Y(_0340_),
    .B1(net764),
    .B2(\cpu_instance.registers_instance.register_bank[8][2] ),
    .A2(_1699_),
    .A1(\cpu_instance.registers_instance.register_bank[11][2] ));
 sg13g2_nand4_1 _2851_ (.B(_0338_),
    .C(_0339_),
    .A(_0333_),
    .Y(_0341_),
    .D(_0340_));
 sg13g2_nor3_2 _2852_ (.A(net757),
    .B(_0337_),
    .C(_0341_),
    .Y(_0342_));
 sg13g2_a21o_1 _2853_ (.A2(net757),
    .A1(_0004_),
    .B1(net799),
    .X(_0343_));
 sg13g2_o21ai_1 _2854_ (.B1(_0331_),
    .Y(_0344_),
    .A1(_0342_),
    .A2(_0343_));
 sg13g2_a21oi_1 _2855_ (.A1(_1573_),
    .A2(\cpu_instance.reg_2_out_sel[1] ),
    .Y(_0345_),
    .B1(\cpu_instance.reg_2_out_sel[0] ));
 sg13g2_a221oi_1 _2856_ (.B2(uo_out[2]),
    .C1(_0345_),
    .B1(_1728_),
    .A1(\cpu_instance.registers_instance.registers[1][2] ),
    .Y(_0346_),
    .A2(net797));
 sg13g2_a21oi_2 _2857_ (.B1(_0346_),
    .Y(_0347_),
    .A2(_1727_),
    .A1(_0005_));
 sg13g2_inv_1 _2858_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_nand2_1 _2859_ (.Y(_0349_),
    .A(net724),
    .B(_0347_));
 sg13g2_nand2b_1 _2860_ (.Y(_0350_),
    .B(_0348_),
    .A_N(net724));
 sg13g2_xnor2_1 _2861_ (.Y(_0351_),
    .A(net724),
    .B(_0347_));
 sg13g2_o21ai_1 _2862_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_0327_),
    .A2(_0329_));
 sg13g2_and2_1 _2863_ (.A(net724),
    .B(_0348_),
    .X(_0353_));
 sg13g2_a221oi_1 _2864_ (.B2(_0350_),
    .C1(_1904_),
    .B1(_0349_),
    .A1(_0328_),
    .Y(_0354_),
    .A2(_0330_));
 sg13g2_a21oi_1 _2865_ (.A1(_1905_),
    .A2(_0353_),
    .Y(_0355_),
    .B1(_0354_));
 sg13g2_a21o_1 _2866_ (.A2(_0353_),
    .A1(_1905_),
    .B1(_1902_),
    .X(_0356_));
 sg13g2_o21ai_1 _2867_ (.B1(_1884_),
    .Y(_0357_),
    .A1(_0354_),
    .A2(_0356_));
 sg13g2_nand2_1 _2868_ (.Y(_0358_),
    .A(_1876_),
    .B(_1880_));
 sg13g2_nand2_1 _2869_ (.Y(_0359_),
    .A(_0357_),
    .B(_0358_));
 sg13g2_a22oi_1 _2870_ (.Y(_0360_),
    .B1(_1876_),
    .B2(_1880_),
    .A2(_1860_),
    .A1(net726));
 sg13g2_a21oi_1 _2871_ (.A1(_0357_),
    .A2(_0360_),
    .Y(_0361_),
    .B1(_1861_));
 sg13g2_a221oi_1 _2872_ (.B2(_0360_),
    .C1(_1861_),
    .B1(_0357_),
    .A1(_1834_),
    .Y(_0362_),
    .A2(_1836_));
 sg13g2_nor2_1 _2873_ (.A(_1829_),
    .B(_1833_),
    .Y(_0363_));
 sg13g2_or3_1 _2874_ (.A(_1813_),
    .B(_0362_),
    .C(_0363_),
    .X(_0364_));
 sg13g2_o21ai_1 _2875_ (.B1(_1813_),
    .Y(_0365_),
    .A1(_0362_),
    .A2(_0363_));
 sg13g2_nand2_1 _2876_ (.Y(_0366_),
    .A(_1735_),
    .B(_0365_));
 sg13g2_nand3_1 _2877_ (.B(_0364_),
    .C(_0365_),
    .A(_1735_),
    .Y(_0367_));
 sg13g2_nor2_2 _2878_ (.A(_1676_),
    .B(_1737_),
    .Y(_0368_));
 sg13g2_nand3_1 _2879_ (.B(\cpu_instance.alu_instance.op[0] ),
    .C(_1734_),
    .A(\cpu_instance.alu_instance.op[1] ),
    .Y(_0369_));
 sg13g2_nand2_2 _2880_ (.Y(_0370_),
    .A(_1788_),
    .B(_0369_));
 sg13g2_and2_1 _2881_ (.A(_1678_),
    .B(_1810_),
    .X(_0371_));
 sg13g2_nand2_1 _2882_ (.Y(_0372_),
    .A(_1746_),
    .B(_1787_));
 sg13g2_o21ai_1 _2883_ (.B1(_0372_),
    .Y(_0373_),
    .A1(_1742_),
    .A2(_1787_));
 sg13g2_a221oi_1 _2884_ (.B2(_0370_),
    .C1(_0371_),
    .B1(_1830_),
    .A1(_1725_),
    .Y(_0374_),
    .A2(_1765_));
 sg13g2_o21ai_1 _2885_ (.B1(_0373_),
    .Y(_0375_),
    .A1(_1769_),
    .A2(_1811_));
 sg13g2_a21oi_1 _2886_ (.A1(_1812_),
    .A2(_0368_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_nand2_1 _2887_ (.Y(_0377_),
    .A(net726),
    .B(_1859_));
 sg13g2_nand2b_1 _2888_ (.Y(_0378_),
    .B(_1860_),
    .A_N(net726));
 sg13g2_nand3_1 _2889_ (.B(_1909_),
    .C(_0325_),
    .A(_1732_),
    .Y(_0379_));
 sg13g2_a21oi_1 _2890_ (.A1(_1732_),
    .A2(_0325_),
    .Y(_0380_),
    .B1(_1908_));
 sg13g2_or2_1 _2891_ (.X(_0381_),
    .B(_0380_),
    .A(_0351_));
 sg13g2_a22oi_1 _2892_ (.Y(_0382_),
    .B1(net724),
    .B2(_0347_),
    .A2(_1901_),
    .A1(net725));
 sg13g2_o21ai_1 _2893_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0351_),
    .A2(_0380_));
 sg13g2_nand3_1 _2894_ (.B(_1903_),
    .C(_0383_),
    .A(_1883_),
    .Y(_0384_));
 sg13g2_nand2_1 _2895_ (.Y(_0385_),
    .A(_1881_),
    .B(_0384_));
 sg13g2_and2_1 _2896_ (.A(_1881_),
    .B(_0377_),
    .X(_0386_));
 sg13g2_a22oi_1 _2897_ (.Y(_0387_),
    .B1(_0384_),
    .B2(_0386_),
    .A2(_1860_),
    .A1(_1856_));
 sg13g2_a221oi_1 _2898_ (.B2(_0386_),
    .C1(_1837_),
    .B1(_0384_),
    .A1(_1856_),
    .Y(_0388_),
    .A2(_1860_));
 sg13g2_or3_1 _2899_ (.A(_1812_),
    .B(_1835_),
    .C(_0388_),
    .X(_0389_));
 sg13g2_o21ai_1 _2900_ (.B1(_1812_),
    .Y(_0390_),
    .A1(_1835_),
    .A2(_0388_));
 sg13g2_nor3_2 _2901_ (.A(\cpu_instance.alu_instance.op[3] ),
    .B(\cpu_instance.alu_instance.op[2] ),
    .C(_1737_),
    .Y(_0391_));
 sg13g2_inv_1 _2902_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_nand3_1 _2903_ (.B(_0390_),
    .C(_0391_),
    .A(_0389_),
    .Y(_0393_));
 sg13g2_nand4_1 _2904_ (.B(_0374_),
    .C(_0376_),
    .A(_0367_),
    .Y(_0394_),
    .D(_0393_));
 sg13g2_and2_1 _2905_ (.A(\cpu_instance.mem_instance.bus_data_out[7] ),
    .B(_1792_),
    .X(_0395_));
 sg13g2_nor2b_2 _2906_ (.A(\cpu_instance.mux_instance.sel[0] ),
    .B_N(\cpu_instance.mux_instance.sel[1] ),
    .Y(_0396_));
 sg13g2_a221oi_1 _2907_ (.B2(net6),
    .C1(_0395_),
    .B1(_0396_),
    .A1(_1674_),
    .Y(_0397_),
    .A2(_0394_));
 sg13g2_xor2_1 _2908_ (.B(_0361_),
    .A(_1837_),
    .X(_0398_));
 sg13g2_nand2b_1 _2909_ (.Y(_0399_),
    .B(_1837_),
    .A_N(_0387_));
 sg13g2_nand3b_1 _2910_ (.B(_0391_),
    .C(_0399_),
    .Y(_0400_),
    .A_N(_0388_));
 sg13g2_a22oi_1 _2911_ (.Y(_0401_),
    .B1(net726),
    .B2(_0370_),
    .A2(_1787_),
    .A1(_1767_));
 sg13g2_nand3_1 _2912_ (.B(_1836_),
    .C(_0368_),
    .A(_1834_),
    .Y(_0402_));
 sg13g2_nand2_1 _2913_ (.Y(_0403_),
    .A(_1743_),
    .B(_1829_));
 sg13g2_o21ai_1 _2914_ (.B1(_0403_),
    .Y(_0404_),
    .A1(_1745_),
    .A2(_1829_));
 sg13g2_a22oi_1 _2915_ (.Y(_0405_),
    .B1(_1836_),
    .B2(_1678_),
    .A2(_1835_),
    .A1(_1770_));
 sg13g2_nand4_1 _2916_ (.B(_0402_),
    .C(_0404_),
    .A(_0401_),
    .Y(_0406_),
    .D(_0405_));
 sg13g2_a21oi_2 _2917_ (.B1(_0406_),
    .Y(_0407_),
    .A2(_0398_),
    .A1(_1735_));
 sg13g2_nand2_1 _2918_ (.Y(_0408_),
    .A(_0400_),
    .B(_0407_));
 sg13g2_a21oi_1 _2919_ (.A1(_0400_),
    .A2(_0407_),
    .Y(_0409_),
    .B1(_1675_));
 sg13g2_a221oi_1 _2920_ (.B2(net5),
    .C1(_0409_),
    .B1(_0396_),
    .A1(\cpu_instance.mem_instance.bus_data_out[6] ),
    .Y(_0410_),
    .A2(_1792_));
 sg13g2_inv_4 _2921_ (.A(net689),
    .Y(_0411_));
 sg13g2_nand2_2 _2922_ (.Y(_0412_),
    .A(_0377_),
    .B(_0378_));
 sg13g2_xor2_1 _2923_ (.B(_0412_),
    .A(_0359_),
    .X(_0413_));
 sg13g2_nor3_1 _2924_ (.A(_1676_),
    .B(_1737_),
    .C(_0412_),
    .Y(_0414_));
 sg13g2_nand3_1 _2925_ (.B(net726),
    .C(_1859_),
    .A(_1770_),
    .Y(_0415_));
 sg13g2_nand2_1 _2926_ (.Y(_0416_),
    .A(_1746_),
    .B(net726));
 sg13g2_o21ai_1 _2927_ (.B1(_0416_),
    .Y(_0417_),
    .A1(_1742_),
    .A2(net726));
 sg13g2_nand2_1 _2928_ (.Y(_0418_),
    .A(_1876_),
    .B(_0370_));
 sg13g2_a221oi_1 _2929_ (.B2(_1678_),
    .C1(_0414_),
    .B1(_0378_),
    .A1(_1767_),
    .Y(_0419_),
    .A2(_1830_));
 sg13g2_nand4_1 _2930_ (.B(_0417_),
    .C(_0418_),
    .A(_0415_),
    .Y(_0420_),
    .D(_0419_));
 sg13g2_xnor2_1 _2931_ (.Y(_0421_),
    .A(_0385_),
    .B(_0412_));
 sg13g2_a221oi_1 _2932_ (.B2(_0391_),
    .C1(_0420_),
    .B1(_0421_),
    .A1(_1735_),
    .Y(_0422_),
    .A2(_0413_));
 sg13g2_nor2_1 _2933_ (.A(_1675_),
    .B(_0422_),
    .Y(_0423_));
 sg13g2_a22oi_1 _2934_ (.Y(_0424_),
    .B1(_0396_),
    .B2(net4),
    .A2(_1792_),
    .A1(\cpu_instance.mem_instance.bus_data_out[5] ));
 sg13g2_nor2b_1 _2935_ (.A(_0423_),
    .B_N(_0424_),
    .Y(_0425_));
 sg13g2_o21ai_1 _2936_ (.B1(_0424_),
    .Y(_0426_),
    .A1(_1675_),
    .A2(_0422_));
 sg13g2_or3_1 _2937_ (.A(_1884_),
    .B(_0354_),
    .C(_0356_),
    .X(_0427_));
 sg13g2_nand3_1 _2938_ (.B(_0357_),
    .C(_0427_),
    .A(_1735_),
    .Y(_0428_));
 sg13g2_a21o_1 _2939_ (.A2(_0383_),
    .A1(_1903_),
    .B1(_1883_),
    .X(_0429_));
 sg13g2_nand3_1 _2940_ (.B(_0391_),
    .C(_0429_),
    .A(_0384_),
    .Y(_0430_));
 sg13g2_nor2_1 _2941_ (.A(_1769_),
    .B(_1881_),
    .Y(_0431_));
 sg13g2_nand2_1 _2942_ (.Y(_0432_),
    .A(_1745_),
    .B(_1876_));
 sg13g2_a221oi_1 _2943_ (.B2(_0370_),
    .C1(_0431_),
    .B1(net725),
    .A1(_1767_),
    .Y(_0433_),
    .A2(net726));
 sg13g2_o21ai_1 _2944_ (.B1(_0432_),
    .Y(_0434_),
    .A1(_1743_),
    .A2(_1876_));
 sg13g2_a221oi_1 _2945_ (.B2(_0368_),
    .C1(_0434_),
    .B1(_1883_),
    .A1(_1678_),
    .Y(_0435_),
    .A2(_1882_));
 sg13g2_nand4_1 _2946_ (.B(_0430_),
    .C(_0433_),
    .A(_0428_),
    .Y(_0436_),
    .D(_0435_));
 sg13g2_and2_1 _2947_ (.A(\cpu_instance.mem_instance.bus_data_out[4] ),
    .B(_1792_),
    .X(_0437_));
 sg13g2_a221oi_1 _2948_ (.B2(_1674_),
    .C1(_0437_),
    .B1(_0436_),
    .A1(net3),
    .Y(_0438_),
    .A2(_0396_));
 sg13g2_inv_4 _2949_ (.A(net702),
    .Y(_0439_));
 sg13g2_xnor2_1 _2950_ (.Y(_0440_),
    .A(\cpu_instance.ctrl_instance.flag_zero ),
    .B(net704));
 sg13g2_xor2_1 _2951_ (.B(_0426_),
    .A(\cpu_instance.ctrl_instance.flag_carry ),
    .X(_0441_));
 sg13g2_a21oi_2 _2952_ (.B1(net690),
    .Y(_0442_),
    .A2(_0441_),
    .A1(_0440_));
 sg13g2_nand2b_2 _2953_ (.Y(_0443_),
    .B(_0442_),
    .A_N(net693));
 sg13g2_nor2_2 _2954_ (.A(net693),
    .B(_0411_),
    .Y(_0444_));
 sg13g2_nand3_1 _2955_ (.B(net704),
    .C(_0444_),
    .A(_0426_),
    .Y(_0445_));
 sg13g2_nand2_1 _2956_ (.Y(_0446_),
    .A(_0443_),
    .B(_0445_));
 sg13g2_nor2_2 _2957_ (.A(\cpu_instance.ctrl_instance.state[3] ),
    .B(\cpu_instance.ctrl_instance.state[2] ),
    .Y(_0447_));
 sg13g2_nand3_1 _2958_ (.B(\cpu_instance.ctrl_instance.state[0] ),
    .C(_0447_),
    .A(_1597_),
    .Y(_0448_));
 sg13g2_nand2_2 _2959_ (.Y(_0449_),
    .A(net693),
    .B(net690));
 sg13g2_inv_2 _2960_ (.Y(_0450_),
    .A(_0449_));
 sg13g2_nor3_2 _2961_ (.A(net857),
    .B(_0448_),
    .C(_0450_),
    .Y(_0451_));
 sg13g2_nand2_1 _2962_ (.Y(_0452_),
    .A(_0446_),
    .B(_0451_));
 sg13g2_nor4_2 _2963_ (.A(\cpu_instance.ctrl_instance.state[3] ),
    .B(\cpu_instance.ctrl_instance.state[2] ),
    .C(_1597_),
    .Y(_0453_),
    .D(\cpu_instance.ctrl_instance.state[0] ));
 sg13g2_nand3_1 _2964_ (.B(_1598_),
    .C(_0447_),
    .A(\cpu_instance.ctrl_instance.state[1] ),
    .Y(_0454_));
 sg13g2_nor2b_2 _2965_ (.A(\cpu_instance.ctrl_instance.state[3] ),
    .B_N(\cpu_instance.ctrl_instance.state[2] ),
    .Y(_0455_));
 sg13g2_nor2_1 _2966_ (.A(_0453_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_a21oi_2 _2967_ (.B1(net857),
    .Y(_0457_),
    .A2(_0456_),
    .A1(net781));
 sg13g2_and2_1 _2968_ (.A(_1615_),
    .B(_0457_),
    .X(_0458_));
 sg13g2_nand2_1 _2969_ (.Y(_0459_),
    .A(_1615_),
    .B(_0457_));
 sg13g2_nor2_1 _2970_ (.A(\cpu_instance.ctrl_instance.state[1] ),
    .B(\cpu_instance.ctrl_instance.state[0] ),
    .Y(_0460_));
 sg13g2_and3_1 _2971_ (.X(_0461_),
    .A(net833),
    .B(_0447_),
    .C(_0460_));
 sg13g2_a221oi_1 _2972_ (.B2(_0457_),
    .C1(_0461_),
    .B1(_1615_),
    .A1(net660),
    .Y(_0462_),
    .A2(net855));
 sg13g2_a221oi_1 _2973_ (.B2(_0452_),
    .C1(net826),
    .B1(_0462_),
    .A1(_1598_),
    .Y(_0036_),
    .A2(_0458_));
 sg13g2_nor2_1 _2974_ (.A(net699),
    .B(_0439_),
    .Y(_0463_));
 sg13g2_nand2_2 _2975_ (.Y(_0464_),
    .A(_0444_),
    .B(_0463_));
 sg13g2_and2_1 _2976_ (.A(_0443_),
    .B(_0464_),
    .X(_0465_));
 sg13g2_nand2_1 _2977_ (.Y(_0466_),
    .A(_0443_),
    .B(_0464_));
 sg13g2_o21ai_1 _2978_ (.B1(_0451_),
    .Y(_0467_),
    .A1(net693),
    .A2(_0466_));
 sg13g2_a21oi_1 _2979_ (.A1(net655),
    .A2(net856),
    .Y(_0468_),
    .B1(_0458_));
 sg13g2_a221oi_1 _2980_ (.B2(_0468_),
    .C1(net825),
    .B1(_0467_),
    .A1(_1597_),
    .Y(_0037_),
    .A2(_0458_));
 sg13g2_nand2_1 _2981_ (.Y(_0469_),
    .A(net699),
    .B(_0439_));
 sg13g2_nand2_1 _2982_ (.Y(_0470_),
    .A(_0444_),
    .B(_0469_));
 sg13g2_nand2_1 _2983_ (.Y(_0471_),
    .A(_0443_),
    .B(_0470_));
 sg13g2_a221oi_1 _2984_ (.B2(_0471_),
    .C1(_0458_),
    .B1(_0451_),
    .A1(\cpu_instance.ctrl_instance.state[3] ),
    .Y(_0472_),
    .A2(net855));
 sg13g2_o21ai_1 _2985_ (.B1(net895),
    .Y(_0473_),
    .A1(net655),
    .A2(_0459_));
 sg13g2_nor2_1 _2986_ (.A(_0472_),
    .B(_0473_),
    .Y(_0038_));
 sg13g2_nor2_1 _2987_ (.A(_0457_),
    .B(_0461_),
    .Y(_0474_));
 sg13g2_nand2_1 _2988_ (.Y(_0475_),
    .A(net693),
    .B(_0411_));
 sg13g2_nor2_1 _2989_ (.A(_0442_),
    .B(net781),
    .Y(_0476_));
 sg13g2_nand3_1 _2990_ (.B(_0475_),
    .C(_0476_),
    .A(_0470_),
    .Y(_0477_));
 sg13g2_a21oi_1 _2991_ (.A1(_0456_),
    .A2(_0477_),
    .Y(_0478_),
    .B1(_0474_));
 sg13g2_a21oi_1 _2992_ (.A1(net500),
    .A2(net856),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_nor3_1 _2993_ (.A(net825),
    .B(_0458_),
    .C(_0479_),
    .Y(_0039_));
 sg13g2_nand2_1 _2994_ (.Y(_0480_),
    .A(net699),
    .B(_0450_));
 sg13g2_a21oi_1 _2995_ (.A1(_0464_),
    .A2(_0480_),
    .Y(_0481_),
    .B1(_0000_));
 sg13g2_nor2_1 _2996_ (.A(net781),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_and2_1 _2997_ (.A(_1597_),
    .B(_0455_),
    .X(_0483_));
 sg13g2_a21oi_1 _2998_ (.A1(_0447_),
    .A2(_0460_),
    .Y(_0484_),
    .B1(_0483_));
 sg13g2_nand3_1 _2999_ (.B(\cpu_instance.ctrl_instance.state[0] ),
    .C(_0455_),
    .A(\cpu_instance.ctrl_instance.state[1] ),
    .Y(_0485_));
 sg13g2_and2_1 _3000_ (.A(_0484_),
    .B(_0485_),
    .X(_0486_));
 sg13g2_nand2_1 _3001_ (.Y(_0487_),
    .A(_0454_),
    .B(_0485_));
 sg13g2_a21oi_1 _3002_ (.A1(_0000_),
    .A2(_0487_),
    .Y(_0488_),
    .B1(_0482_));
 sg13g2_nand2_1 _3003_ (.Y(_0489_),
    .A(_0484_),
    .B(_0488_));
 sg13g2_nor2_2 _3004_ (.A(net856),
    .B(_0454_),
    .Y(_0490_));
 sg13g2_a21o_2 _3005_ (.A2(_0454_),
    .A1(net781),
    .B1(net857),
    .X(_0491_));
 sg13g2_o21ai_1 _3006_ (.B1(_0491_),
    .Y(_0492_),
    .A1(net856),
    .A2(_0486_));
 sg13g2_a22oi_1 _3007_ (.Y(_0493_),
    .B1(_0489_),
    .B2(_0492_),
    .A2(net595),
    .A1(net862));
 sg13g2_nor2_1 _3008_ (.A(net829),
    .B(net596),
    .Y(_0040_));
 sg13g2_nor2_2 _3009_ (.A(_0000_),
    .B(net781),
    .Y(_0494_));
 sg13g2_or2_2 _3010_ (.X(_0495_),
    .B(net781),
    .A(_0000_));
 sg13g2_nor2_1 _3011_ (.A(_0480_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_nand3_1 _3012_ (.B(_0450_),
    .C(_0494_),
    .A(net699),
    .Y(_0497_));
 sg13g2_a22oi_1 _3013_ (.Y(_0498_),
    .B1(_0492_),
    .B2(_0496_),
    .A2(\cpu_instance.reg_2_out_sel[0] ),
    .A1(net862));
 sg13g2_nor2_1 _3014_ (.A(net829),
    .B(_0498_),
    .Y(_0041_));
 sg13g2_nand4_1 _3015_ (.B(_0330_),
    .C(_0349_),
    .A(_0328_),
    .Y(_0499_),
    .D(_0350_));
 sg13g2_nand3_1 _3016_ (.B(_0352_),
    .C(_0499_),
    .A(_1735_),
    .Y(_0500_));
 sg13g2_nand2b_1 _3017_ (.Y(_0501_),
    .B(_0368_),
    .A_N(_0351_));
 sg13g2_nand2_1 _3018_ (.Y(_0502_),
    .A(_1678_),
    .B(_0350_));
 sg13g2_a21oi_1 _3019_ (.A1(_1770_),
    .A2(_0347_),
    .Y(_0503_),
    .B1(_1745_));
 sg13g2_nand2_1 _3020_ (.Y(_0504_),
    .A(_0344_),
    .B(_0503_));
 sg13g2_o21ai_1 _3021_ (.B1(_0504_),
    .Y(_0505_),
    .A1(_1742_),
    .A2(net724));
 sg13g2_a22oi_1 _3022_ (.Y(_0506_),
    .B1(_0370_),
    .B2(_1762_),
    .A2(_1899_),
    .A1(_1767_));
 sg13g2_and4_1 _3023_ (.A(_0501_),
    .B(_0502_),
    .C(_0505_),
    .D(_0506_),
    .X(_0507_));
 sg13g2_nand2_1 _3024_ (.Y(_0508_),
    .A(_0351_),
    .B(_0380_));
 sg13g2_nand3_1 _3025_ (.B(_0391_),
    .C(_0508_),
    .A(_0381_),
    .Y(_0509_));
 sg13g2_nand3_1 _3026_ (.B(_0507_),
    .C(_0509_),
    .A(_0500_),
    .Y(_0510_));
 sg13g2_and2_1 _3027_ (.A(\cpu_instance.mem_instance.bus_data_out[2] ),
    .B(_1792_),
    .X(_0511_));
 sg13g2_a221oi_1 _3028_ (.B2(_1674_),
    .C1(_0511_),
    .B1(_0510_),
    .A1(net1),
    .Y(_0512_),
    .A2(_0396_));
 sg13g2_inv_2 _3029_ (.Y(_0513_),
    .A(net712));
 sg13g2_nor3_1 _3030_ (.A(_1908_),
    .B(_1910_),
    .C(_0326_),
    .Y(_0514_));
 sg13g2_nor3_1 _3031_ (.A(_1736_),
    .B(_0327_),
    .C(_0514_),
    .Y(_0515_));
 sg13g2_a21o_1 _3032_ (.A2(_0325_),
    .A1(_1909_),
    .B1(_1732_),
    .X(_0516_));
 sg13g2_and3_1 _3033_ (.X(_0517_),
    .A(_0379_),
    .B(_0391_),
    .C(_0516_));
 sg13g2_a22oi_1 _3034_ (.Y(_0518_),
    .B1(net724),
    .B2(_1767_),
    .A2(_1908_),
    .A1(_1770_));
 sg13g2_nand3_1 _3035_ (.B(_0325_),
    .C(_0368_),
    .A(_1909_),
    .Y(_0519_));
 sg13g2_nand2_1 _3036_ (.Y(_0520_),
    .A(_1725_),
    .B(_0370_));
 sg13g2_mux2_1 _3037_ (.A0(_1743_),
    .A1(_1746_),
    .S(_1762_),
    .X(_0521_));
 sg13g2_o21ai_1 _3038_ (.B1(_0519_),
    .Y(_0522_),
    .A1(_1679_),
    .A2(_1910_));
 sg13g2_nand3_1 _3039_ (.B(_0520_),
    .C(_0521_),
    .A(_0518_),
    .Y(_0523_));
 sg13g2_or4_2 _3040_ (.A(_0515_),
    .B(_0517_),
    .C(_0522_),
    .D(_0523_),
    .X(_0524_));
 sg13g2_a22oi_1 _3041_ (.Y(_0525_),
    .B1(_0524_),
    .B2(_1674_),
    .A2(_1792_),
    .A1(\cpu_instance.mem_instance.bus_data_out[1] ));
 sg13g2_nand3b_1 _3042_ (.B(_0469_),
    .C(net690),
    .Y(_0526_),
    .A_N(_0463_));
 sg13g2_nor3_1 _3043_ (.A(net694),
    .B(net716),
    .C(_0526_),
    .Y(_0527_));
 sg13g2_o21ai_1 _3044_ (.B1(_0454_),
    .Y(_0528_),
    .A1(_0480_),
    .A2(net713));
 sg13g2_nand2_1 _3045_ (.Y(_0529_),
    .A(_0349_),
    .B(_0381_));
 sg13g2_xnor2_1 _3046_ (.Y(_0530_),
    .A(_1904_),
    .B(_0529_));
 sg13g2_nand3_1 _3047_ (.B(net725),
    .C(_1901_),
    .A(_1770_),
    .Y(_0531_));
 sg13g2_nand2_1 _3048_ (.Y(_0532_),
    .A(_1678_),
    .B(_1903_));
 sg13g2_a22oi_1 _3049_ (.Y(_0533_),
    .B1(net724),
    .B2(_0370_),
    .A2(_1899_),
    .A1(_1745_));
 sg13g2_nor2_1 _3050_ (.A(_1743_),
    .B(net725),
    .Y(_0534_));
 sg13g2_a21oi_1 _3051_ (.A1(_1767_),
    .A2(_1876_),
    .Y(_0535_),
    .B1(_0534_));
 sg13g2_nand4_1 _3052_ (.B(_0532_),
    .C(_0533_),
    .A(_0531_),
    .Y(_0536_),
    .D(_0535_));
 sg13g2_nor2_1 _3053_ (.A(_1905_),
    .B(_0353_),
    .Y(_0537_));
 sg13g2_a21oi_1 _3054_ (.A1(_0352_),
    .A2(_0537_),
    .Y(_0538_),
    .B1(_1736_));
 sg13g2_a221oi_1 _3055_ (.B2(_0355_),
    .C1(_0536_),
    .B1(_0538_),
    .A1(_1904_),
    .Y(_0539_),
    .A2(_0368_));
 sg13g2_o21ai_1 _3056_ (.B1(_0539_),
    .Y(_0540_),
    .A1(_0392_),
    .A2(_0530_));
 sg13g2_and2_1 _3057_ (.A(\cpu_instance.mem_instance.bus_data_out[3] ),
    .B(_1792_),
    .X(_0541_));
 sg13g2_a221oi_1 _3058_ (.B2(_1674_),
    .C1(_0541_),
    .B1(_0540_),
    .A1(net2),
    .Y(_0542_),
    .A2(_0396_));
 sg13g2_nor2_1 _3059_ (.A(_0000_),
    .B(_0454_),
    .Y(_0543_));
 sg13g2_nor2_1 _3060_ (.A(net862),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_nand2_1 _3061_ (.Y(_0545_),
    .A(net835),
    .B(_0543_));
 sg13g2_a221oi_1 _3062_ (.B2(_0495_),
    .C1(net862),
    .B1(_0544_),
    .A1(_0453_),
    .Y(_0546_),
    .A2(_0542_));
 sg13g2_o21ai_1 _3063_ (.B1(_0546_),
    .Y(_0547_),
    .A1(_0527_),
    .A2(_0528_));
 sg13g2_nor2b_1 _3064_ (.A(net864),
    .B_N(\cpu_instance.ctrl_instance.use_register_bank_in ),
    .Y(_0548_));
 sg13g2_a22oi_1 _3065_ (.Y(_0549_),
    .B1(_0483_),
    .B2(_0548_),
    .A2(net863),
    .A1(net634));
 sg13g2_a21oi_1 _3066_ (.A1(_0547_),
    .A2(_0549_),
    .Y(_0042_),
    .B1(net829));
 sg13g2_and3_2 _3067_ (.X(_0550_),
    .A(\cpu_instance.ctrl_instance.state[1] ),
    .B(net834),
    .C(_0455_));
 sg13g2_a22oi_1 _3068_ (.Y(_0551_),
    .B1(_0550_),
    .B2(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .A2(net862),
    .A1(net675));
 sg13g2_nor2_1 _3069_ (.A(_0464_),
    .B(net716),
    .Y(_0552_));
 sg13g2_o21ai_1 _3070_ (.B1(_0454_),
    .Y(_0553_),
    .A1(net718),
    .A2(_0443_));
 sg13g2_nor2_1 _3071_ (.A(_0454_),
    .B(_0513_),
    .Y(_0554_));
 sg13g2_nor3_1 _3072_ (.A(_1615_),
    .B(_0491_),
    .C(_0554_),
    .Y(_0555_));
 sg13g2_o21ai_1 _3073_ (.B1(_0555_),
    .Y(_0556_),
    .A1(_0552_),
    .A2(_0553_));
 sg13g2_a21oi_1 _3074_ (.A1(net676),
    .A2(_0556_),
    .Y(_0043_),
    .B1(net829));
 sg13g2_nand4_1 _3075_ (.B(net694),
    .C(_0411_),
    .A(net835),
    .Y(_0557_),
    .D(_0494_));
 sg13g2_a22oi_1 _3076_ (.Y(_0558_),
    .B1(_0490_),
    .B2(net663),
    .A2(net864),
    .A1(net677));
 sg13g2_o21ai_1 _3077_ (.B1(_0558_),
    .Y(_0559_),
    .A1(net713),
    .A2(_0557_));
 sg13g2_and2_1 _3078_ (.A(net898),
    .B(_0559_),
    .X(_0044_));
 sg13g2_a22oi_1 _3079_ (.Y(_0560_),
    .B1(_0490_),
    .B2(net677),
    .A2(net864),
    .A1(net678));
 sg13g2_o21ai_1 _3080_ (.B1(_0560_),
    .Y(_0561_),
    .A1(_0542_),
    .A2(_0557_));
 sg13g2_and2_1 _3081_ (.A(net898),
    .B(_0561_),
    .X(_0045_));
 sg13g2_a22oi_1 _3082_ (.Y(_0562_),
    .B1(_0490_),
    .B2(net678),
    .A2(net864),
    .A1(\cpu_instance.alu_instance.op[3] ));
 sg13g2_o21ai_1 _3083_ (.B1(_0562_),
    .Y(_0563_),
    .A1(net704),
    .A2(_0557_));
 sg13g2_and2_1 _3084_ (.A(net898),
    .B(_0563_),
    .X(_0046_));
 sg13g2_a22oi_1 _3085_ (.Y(_0564_),
    .B1(_0490_),
    .B2(net906),
    .A2(net864),
    .A1(net815));
 sg13g2_o21ai_1 _3086_ (.B1(_0564_),
    .Y(_0565_),
    .A1(net688),
    .A2(_0557_));
 sg13g2_and2_1 _3087_ (.A(net903),
    .B(_0565_),
    .X(_0047_));
 sg13g2_a21oi_1 _3088_ (.A1(_1787_),
    .A2(_1809_),
    .Y(_0566_),
    .B1(_0366_));
 sg13g2_a21oi_1 _3089_ (.A1(_1811_),
    .A2(_0390_),
    .Y(_0567_),
    .B1(_0392_));
 sg13g2_nand2b_1 _3090_ (.Y(_0568_),
    .B(_1787_),
    .A_N(_0369_));
 sg13g2_a21oi_1 _3091_ (.A1(_1725_),
    .A2(_1766_),
    .Y(_0569_),
    .B1(_0545_));
 sg13g2_nand2_1 _3092_ (.Y(_0570_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_nor3_2 _3093_ (.A(_0566_),
    .B(_0567_),
    .C(_0570_),
    .Y(_0571_));
 sg13g2_nor3_1 _3094_ (.A(net615),
    .B(net862),
    .C(_0543_),
    .Y(_0572_));
 sg13g2_o21ai_1 _3095_ (.B1(net903),
    .Y(_0573_),
    .A1(net407),
    .A2(net835));
 sg13g2_nor3_1 _3096_ (.A(_0571_),
    .B(net616),
    .C(_0573_),
    .Y(_0048_));
 sg13g2_or2_1 _3097_ (.X(_0574_),
    .B(_0524_),
    .A(_1791_));
 sg13g2_nor4_1 _3098_ (.A(_0510_),
    .B(_0540_),
    .C(_0545_),
    .D(_0574_),
    .Y(_0575_));
 sg13g2_nand2_1 _3099_ (.Y(_0576_),
    .A(_0422_),
    .B(_0575_));
 sg13g2_nor4_1 _3100_ (.A(_0394_),
    .B(_0408_),
    .C(_0436_),
    .D(_0576_),
    .Y(_0577_));
 sg13g2_a221oi_1 _3101_ (.B2(net634),
    .C1(_0577_),
    .B1(_0544_),
    .A1(net615),
    .Y(_0578_),
    .A2(net862));
 sg13g2_nor2_1 _3102_ (.A(net829),
    .B(_0578_),
    .Y(_0049_));
 sg13g2_and2_1 _3103_ (.A(net834),
    .B(_0483_),
    .X(_0579_));
 sg13g2_inv_1 _3104_ (.Y(_0580_),
    .A(_0579_));
 sg13g2_o21ai_1 _3105_ (.B1(\cpu_instance.ctrl_instance.mem_op_done ),
    .Y(_0581_),
    .A1(_0453_),
    .A2(_0483_));
 sg13g2_a22oi_1 _3106_ (.Y(_0582_),
    .B1(_0581_),
    .B2(_0497_),
    .A2(_0580_),
    .A1(_0491_));
 sg13g2_a21oi_1 _3107_ (.A1(net663),
    .A2(net863),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_nor2_1 _3108_ (.A(net829),
    .B(_0583_),
    .Y(_0050_));
 sg13g2_nand2_1 _3109_ (.Y(_0584_),
    .A(\cpu_instance.ctrl_instance.mem_op_done ),
    .B(_0486_));
 sg13g2_a22oi_1 _3110_ (.Y(_0585_),
    .B1(_0492_),
    .B2(_0584_),
    .A2(net581),
    .A1(net856));
 sg13g2_nor2_1 _3111_ (.A(net826),
    .B(net582),
    .Y(_0051_));
 sg13g2_nand3_1 _3112_ (.B(_0463_),
    .C(_0494_),
    .A(_0444_),
    .Y(_0586_));
 sg13g2_nand3_1 _3113_ (.B(_1598_),
    .C(_0455_),
    .A(\cpu_instance.ctrl_instance.state[1] ),
    .Y(_0587_));
 sg13g2_a21oi_1 _3114_ (.A1(_0586_),
    .A2(_0587_),
    .Y(_0588_),
    .B1(_0474_));
 sg13g2_a21oi_1 _3115_ (.A1(net589),
    .A2(net855),
    .Y(_0589_),
    .B1(_0588_));
 sg13g2_nor2_1 _3116_ (.A(net826),
    .B(net590),
    .Y(_0052_));
 sg13g2_nor2_2 _3117_ (.A(_1615_),
    .B(net688),
    .Y(_0590_));
 sg13g2_nor2_2 _3118_ (.A(net856),
    .B(_0485_),
    .Y(_0591_));
 sg13g2_a22oi_1 _3119_ (.Y(_0592_),
    .B1(_0590_),
    .B2(_0591_),
    .A2(net657),
    .A1(net855));
 sg13g2_nor2_1 _3120_ (.A(net830),
    .B(_0592_),
    .Y(_0053_));
 sg13g2_nor2_2 _3121_ (.A(_1615_),
    .B(net690),
    .Y(_0593_));
 sg13g2_a22oi_1 _3122_ (.Y(_0594_),
    .B1(_0591_),
    .B2(_0593_),
    .A2(net444),
    .A1(net855));
 sg13g2_nor2_1 _3123_ (.A(net825),
    .B(_0594_),
    .Y(_0054_));
 sg13g2_nor2_1 _3124_ (.A(net693),
    .B(_0446_),
    .Y(_0595_));
 sg13g2_nand2_1 _3125_ (.Y(_0596_),
    .A(_0449_),
    .B(_0494_));
 sg13g2_nand3b_1 _3126_ (.B(_0460_),
    .C(\cpu_instance.ctrl_instance.state[3] ),
    .Y(_0597_),
    .A_N(\cpu_instance.ctrl_instance.state[2] ));
 sg13g2_o21ai_1 _3127_ (.B1(_0597_),
    .Y(_0598_),
    .A1(_0595_),
    .A2(_0596_));
 sg13g2_nand2_1 _3128_ (.Y(_0599_),
    .A(net835),
    .B(_0598_));
 sg13g2_nor2_2 _3129_ (.A(_1615_),
    .B(net693),
    .Y(_0600_));
 sg13g2_a22oi_1 _3130_ (.Y(_0601_),
    .B1(_0591_),
    .B2(_0600_),
    .A2(net662),
    .A1(net855));
 sg13g2_a21oi_1 _3131_ (.A1(_0599_),
    .A2(_0601_),
    .Y(_0055_),
    .B1(net825));
 sg13g2_or3_1 _3132_ (.A(net688),
    .B(_0495_),
    .C(net701),
    .X(_0602_));
 sg13g2_o21ai_1 _3133_ (.B1(_0449_),
    .Y(_0603_),
    .A1(net713),
    .A2(_0526_));
 sg13g2_nand3_1 _3134_ (.B(_0439_),
    .C(_0490_),
    .A(net651),
    .Y(_0604_));
 sg13g2_a21oi_1 _3135_ (.A1(_0596_),
    .A2(_0602_),
    .Y(_0605_),
    .B1(_0491_));
 sg13g2_a221oi_1 _3136_ (.B2(_0605_),
    .C1(_0579_),
    .B1(_0603_),
    .A1(net820),
    .Y(_0606_),
    .A2(net863));
 sg13g2_a221oi_1 _3137_ (.B2(_0606_),
    .C1(net828),
    .B1(_0604_),
    .A1(_1595_),
    .Y(_0056_),
    .A2(_0579_));
 sg13g2_o21ai_1 _3138_ (.B1(_0449_),
    .Y(_0607_),
    .A1(_0526_),
    .A2(net701));
 sg13g2_a21oi_1 _3139_ (.A1(_0450_),
    .A2(_0469_),
    .Y(_0608_),
    .B1(_0495_));
 sg13g2_a22oi_1 _3140_ (.Y(_0609_),
    .B1(_0607_),
    .B2(_0608_),
    .A2(_0590_),
    .A1(_0453_));
 sg13g2_a22oi_1 _3141_ (.Y(_0610_),
    .B1(_0579_),
    .B2(net820),
    .A2(net863),
    .A1(\cpu_instance.reg_op ));
 sg13g2_o21ai_1 _3142_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_0491_),
    .A2(_0609_));
 sg13g2_and2_1 _3143_ (.A(net899),
    .B(_0611_),
    .X(_0057_));
 sg13g2_nor3_2 _3144_ (.A(net862),
    .B(_0450_),
    .C(_0495_),
    .Y(_0612_));
 sg13g2_or2_1 _3145_ (.X(_0613_),
    .B(_0475_),
    .A(net718));
 sg13g2_o21ai_1 _3146_ (.B1(_0613_),
    .Y(_0614_),
    .A1(_0465_),
    .A2(net713));
 sg13g2_nor2_1 _3147_ (.A(_0490_),
    .B(_0550_),
    .Y(_0615_));
 sg13g2_a22oi_1 _3148_ (.Y(_0616_),
    .B1(_0612_),
    .B2(_0614_),
    .A2(net867),
    .A1(net816));
 sg13g2_o21ai_1 _3149_ (.B1(net899),
    .Y(_0617_),
    .A1(net819),
    .A2(_0615_));
 sg13g2_a21oi_1 _3150_ (.A1(_0615_),
    .A2(_0616_),
    .Y(_0058_),
    .B1(_0617_));
 sg13g2_or2_1 _3151_ (.X(_0618_),
    .B(net716),
    .A(_0475_));
 sg13g2_o21ai_1 _3152_ (.B1(_0618_),
    .Y(_0619_),
    .A1(_0465_),
    .A2(net701));
 sg13g2_a22oi_1 _3153_ (.Y(_0620_),
    .B1(_0612_),
    .B2(_0619_),
    .A2(net867),
    .A1(net821));
 sg13g2_o21ai_1 _3154_ (.B1(net899),
    .Y(_0621_),
    .A1(net816),
    .A2(_0615_));
 sg13g2_a21oi_1 _3155_ (.A1(_0615_),
    .A2(_0620_),
    .Y(_0059_),
    .B1(_0621_));
 sg13g2_nor2_1 _3156_ (.A(_1615_),
    .B(net699),
    .Y(_0622_));
 sg13g2_a21o_1 _3157_ (.A2(_0622_),
    .A1(_0444_),
    .B1(net781),
    .X(_0623_));
 sg13g2_a21oi_1 _3158_ (.A1(_1591_),
    .A2(\cpu_instance.ctrl_instance.mem_op_done ),
    .Y(_0624_),
    .B1(_0485_));
 sg13g2_o21ai_1 _3159_ (.B1(_0455_),
    .Y(_0625_),
    .A1(\cpu_instance.ctrl_instance.state[1] ),
    .A2(_1598_));
 sg13g2_a21oi_1 _3160_ (.A1(net781),
    .A2(_0625_),
    .Y(_0626_),
    .B1(net855));
 sg13g2_nor2b_1 _3161_ (.A(_0624_),
    .B_N(_0626_),
    .Y(_0627_));
 sg13g2_a221oi_1 _3162_ (.B2(_0627_),
    .C1(net825),
    .B1(_0623_),
    .A1(net855),
    .Y(_0060_),
    .A2(_1612_));
 sg13g2_or2_1 _3163_ (.X(_0628_),
    .B(net716),
    .A(net864));
 sg13g2_or3_1 _3164_ (.A(_0443_),
    .B(_0495_),
    .C(net710),
    .X(_0629_));
 sg13g2_a21oi_1 _3165_ (.A1(net865),
    .A2(\cpu_instance.mux_instance.sel[0] ),
    .Y(_0630_),
    .B1(_0591_));
 sg13g2_a221oi_1 _3166_ (.B2(_0630_),
    .C1(net829),
    .B1(_0629_),
    .A1(_1591_),
    .Y(_0061_),
    .A2(_0591_));
 sg13g2_nor2_1 _3167_ (.A(\cpu_instance.mem_instance.addr[24] ),
    .B(_1669_),
    .Y(_0631_));
 sg13g2_nor3_2 _3168_ (.A(\cpu_instance.mem_instance.addr[24] ),
    .B(net837),
    .C(_1669_),
    .Y(_0632_));
 sg13g2_nand2_2 _3169_ (.Y(_0633_),
    .A(net831),
    .B(_0631_));
 sg13g2_nor2_1 _3170_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ),
    .B(net813),
    .Y(_0634_));
 sg13g2_a21oi_2 _3171_ (.B1(_0634_),
    .Y(_0635_),
    .A2(_1590_),
    .A1(net813));
 sg13g2_nand2_1 _3172_ (.Y(_0636_),
    .A(net714),
    .B(_0635_));
 sg13g2_nor2b_1 _3173_ (.A(net714),
    .B_N(_0635_),
    .Y(_0637_));
 sg13g2_xnor2_1 _3174_ (.Y(_0638_),
    .A(net714),
    .B(_0635_));
 sg13g2_nor2_1 _3175_ (.A(_1612_),
    .B(_1665_),
    .Y(_0639_));
 sg13g2_nand2_2 _3176_ (.Y(_0640_),
    .A(\cpu_instance.addr_reg_op[0] ),
    .B(_1664_));
 sg13g2_xor2_1 _3177_ (.B(_0638_),
    .A(_1794_),
    .X(_0641_));
 sg13g2_nor2_1 _3178_ (.A(net767),
    .B(net717),
    .Y(_0642_));
 sg13g2_or2_1 _3179_ (.X(_0643_),
    .B(_0642_),
    .A(_0638_));
 sg13g2_nor2_2 _3180_ (.A(\cpu_instance.addr_reg_op[0] ),
    .B(_1665_),
    .Y(_0644_));
 sg13g2_nand2_2 _3181_ (.Y(_0645_),
    .A(_1612_),
    .B(_1664_));
 sg13g2_a21oi_1 _3182_ (.A1(_0638_),
    .A2(_0642_),
    .Y(_0646_),
    .B1(_0645_));
 sg13g2_a22oi_1 _3183_ (.Y(_0647_),
    .B1(_0643_),
    .B2(_0646_),
    .A2(_0641_),
    .A1(_0639_));
 sg13g2_and2_2 _3184_ (.A(net767),
    .B(_0635_),
    .X(_0648_));
 sg13g2_nand2_1 _3185_ (.Y(_0649_),
    .A(net765),
    .B(_0635_));
 sg13g2_nand2b_2 _3186_ (.Y(_0650_),
    .B(_1672_),
    .A_N(_0635_));
 sg13g2_and2_2 _3187_ (.A(_0649_),
    .B(_0650_),
    .X(_0651_));
 sg13g2_nand2_2 _3188_ (.Y(_0652_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_nand2_2 _3189_ (.Y(_0653_),
    .A(_1666_),
    .B(_0651_));
 sg13g2_a21oi_1 _3190_ (.A1(_0647_),
    .A2(_0653_),
    .Y(_0654_),
    .B1(\cpu_instance.mem_instance.addr[24] ));
 sg13g2_and2_1 _3191_ (.A(net813),
    .B(_1663_),
    .X(_0655_));
 sg13g2_nand2_1 _3192_ (.Y(_0656_),
    .A(net811),
    .B(_1663_));
 sg13g2_nor2_1 _3193_ (.A(net714),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_o21ai_1 _3194_ (.B1(_0632_),
    .Y(_0658_),
    .A1(_0654_),
    .A2(_0657_));
 sg13g2_nor2_1 _3195_ (.A(net837),
    .B(_0631_),
    .Y(_0659_));
 sg13g2_a22oi_1 _3196_ (.Y(_0660_),
    .B1(net743),
    .B2(net397),
    .A2(net841),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ));
 sg13g2_a21oi_1 _3197_ (.A1(_0658_),
    .A2(net398),
    .Y(_0062_),
    .B1(net824));
 sg13g2_mux2_2 _3198_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ),
    .S(net812),
    .X(_0661_));
 sg13g2_and2_1 _3199_ (.A(net712),
    .B(_0661_),
    .X(_0662_));
 sg13g2_nand2b_1 _3200_ (.Y(_0663_),
    .B(_0661_),
    .A_N(net711));
 sg13g2_xor2_1 _3201_ (.B(_0661_),
    .A(net712),
    .X(_0664_));
 sg13g2_o21ai_1 _3202_ (.B1(_0636_),
    .Y(_0665_),
    .A1(_0638_),
    .A2(_0642_));
 sg13g2_xor2_1 _3203_ (.B(_0665_),
    .A(_0664_),
    .X(_0666_));
 sg13g2_xnor2_1 _3204_ (.Y(_0667_),
    .A(_0648_),
    .B(_0661_));
 sg13g2_inv_2 _3205_ (.Y(_0668_),
    .A(net748));
 sg13g2_a21oi_1 _3206_ (.A1(_1794_),
    .A2(_0638_),
    .Y(_0669_),
    .B1(_0637_));
 sg13g2_or2_1 _3207_ (.X(_0670_),
    .B(_0669_),
    .A(_0664_));
 sg13g2_a21oi_1 _3208_ (.A1(_0664_),
    .A2(_0669_),
    .Y(_0671_),
    .B1(_0640_));
 sg13g2_a22oi_1 _3209_ (.Y(_0672_),
    .B1(_0670_),
    .B2(_0671_),
    .A2(_0666_),
    .A1(_0644_));
 sg13g2_o21ai_1 _3210_ (.B1(_0672_),
    .Y(_0673_),
    .A1(net789),
    .A2(net748));
 sg13g2_a22oi_1 _3211_ (.Y(_0674_),
    .B1(_0673_),
    .B2(_1584_),
    .A2(_0655_),
    .A1(_0513_));
 sg13g2_a22oi_1 _3212_ (.Y(_0675_),
    .B1(net743),
    .B2(net658),
    .A2(net841),
    .A1(net572));
 sg13g2_o21ai_1 _3213_ (.B1(_0675_),
    .Y(_0676_),
    .A1(_0633_),
    .A2(_0674_));
 sg13g2_and2_1 _3214_ (.A(net873),
    .B(_0676_),
    .X(_0063_));
 sg13g2_nor2_1 _3215_ (.A(net700),
    .B(_0656_),
    .Y(_0677_));
 sg13g2_o21ai_1 _3216_ (.B1(_0663_),
    .Y(_0678_),
    .A1(_0664_),
    .A2(_0669_));
 sg13g2_mux2_2 _3217_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ),
    .S(net812),
    .X(_0679_));
 sg13g2_nand2_1 _3218_ (.Y(_0680_),
    .A(net700),
    .B(_0679_));
 sg13g2_nor2b_1 _3219_ (.A(net700),
    .B_N(_0679_),
    .Y(_0681_));
 sg13g2_xnor2_1 _3220_ (.Y(_0682_),
    .A(net700),
    .B(_0679_));
 sg13g2_nand2_1 _3221_ (.Y(_0683_),
    .A(_0678_),
    .B(_0682_));
 sg13g2_nor2_1 _3222_ (.A(_0678_),
    .B(_0682_),
    .Y(_0684_));
 sg13g2_nor2_1 _3223_ (.A(_0640_),
    .B(_0684_),
    .Y(_0685_));
 sg13g2_a21oi_2 _3224_ (.B1(_0662_),
    .Y(_0686_),
    .A2(_0665_),
    .A1(_0664_));
 sg13g2_o21ai_1 _3225_ (.B1(_0644_),
    .Y(_0687_),
    .A1(_0682_),
    .A2(_0686_));
 sg13g2_a21oi_1 _3226_ (.A1(_0682_),
    .A2(_0686_),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_a21oi_1 _3227_ (.A1(_0683_),
    .A2(_0685_),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_nand3_1 _3228_ (.B(_0661_),
    .C(_0679_),
    .A(_0648_),
    .Y(_0690_));
 sg13g2_a21o_1 _3229_ (.A2(_0661_),
    .A1(_0648_),
    .B1(_0679_),
    .X(_0691_));
 sg13g2_and2_1 _3230_ (.A(_0690_),
    .B(_0691_),
    .X(_0692_));
 sg13g2_nand2_2 _3231_ (.Y(_0693_),
    .A(_1666_),
    .B(_0692_));
 sg13g2_a21oi_1 _3232_ (.A1(_0689_),
    .A2(_0693_),
    .Y(_0694_),
    .B1(\cpu_instance.mem_instance.addr[24] ));
 sg13g2_o21ai_1 _3233_ (.B1(_0632_),
    .Y(_0695_),
    .A1(_0677_),
    .A2(_0694_));
 sg13g2_a22oi_1 _3234_ (.Y(_0696_),
    .B1(net743),
    .B2(net572),
    .A2(net841),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ));
 sg13g2_a21oi_1 _3235_ (.A1(_0695_),
    .A2(net573),
    .Y(_0064_),
    .B1(net824));
 sg13g2_nand2_1 _3236_ (.Y(_0697_),
    .A(net812),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ));
 sg13g2_o21ai_1 _3237_ (.B1(_0697_),
    .Y(_0698_),
    .A1(_1583_),
    .A2(net812));
 sg13g2_nand2_1 _3238_ (.Y(_0699_),
    .A(net702),
    .B(_0698_));
 sg13g2_inv_1 _3239_ (.Y(_0700_),
    .A(_0699_));
 sg13g2_nand2_1 _3240_ (.Y(_0701_),
    .A(_0439_),
    .B(_0698_));
 sg13g2_xor2_1 _3241_ (.B(_0698_),
    .A(net702),
    .X(_0702_));
 sg13g2_a21oi_2 _3242_ (.B1(_0681_),
    .Y(_0703_),
    .A2(_0682_),
    .A1(_0678_));
 sg13g2_xnor2_1 _3243_ (.Y(_0704_),
    .A(_0702_),
    .B(_0703_));
 sg13g2_nand2b_1 _3244_ (.Y(_0705_),
    .B(_0698_),
    .A_N(_0690_));
 sg13g2_xnor2_1 _3245_ (.Y(_0706_),
    .A(_0690_),
    .B(_0698_));
 sg13g2_o21ai_1 _3246_ (.B1(_0680_),
    .Y(_0707_),
    .A1(_0682_),
    .A2(_0686_));
 sg13g2_nand2_1 _3247_ (.Y(_0708_),
    .A(_0702_),
    .B(_0707_));
 sg13g2_nor2_1 _3248_ (.A(_0702_),
    .B(_0707_),
    .Y(_0709_));
 sg13g2_nor2_1 _3249_ (.A(_0645_),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_a22oi_1 _3250_ (.Y(_0711_),
    .B1(_0708_),
    .B2(_0710_),
    .A2(_0706_),
    .A1(_1666_));
 sg13g2_o21ai_1 _3251_ (.B1(_0711_),
    .Y(_0712_),
    .A1(_0640_),
    .A2(_0704_));
 sg13g2_a22oi_1 _3252_ (.Y(_0713_),
    .B1(_0712_),
    .B2(_1584_),
    .A2(_0655_),
    .A1(_0439_));
 sg13g2_a22oi_1 _3253_ (.Y(_0714_),
    .B1(net743),
    .B2(net666),
    .A2(net841),
    .A1(net441));
 sg13g2_o21ai_1 _3254_ (.B1(_0714_),
    .Y(_0715_),
    .A1(_0633_),
    .A2(_0713_));
 sg13g2_and2_1 _3255_ (.A(net872),
    .B(_0715_),
    .X(_0065_));
 sg13g2_nor2_1 _3256_ (.A(net687),
    .B(_0656_),
    .Y(_0716_));
 sg13g2_mux2_2 _3257_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ),
    .S(net812),
    .X(_0717_));
 sg13g2_inv_2 _3258_ (.Y(_0718_),
    .A(_0717_));
 sg13g2_nand2_1 _3259_ (.Y(_0719_),
    .A(net687),
    .B(_0718_));
 sg13g2_xnor2_1 _3260_ (.Y(_0720_),
    .A(net699),
    .B(_0718_));
 sg13g2_o21ai_1 _3261_ (.B1(_0701_),
    .Y(_0721_),
    .A1(_0702_),
    .A2(_0703_));
 sg13g2_a21oi_1 _3262_ (.A1(_0720_),
    .A2(_0721_),
    .Y(_0722_),
    .B1(_0640_));
 sg13g2_o21ai_1 _3263_ (.B1(_0722_),
    .Y(_0723_),
    .A1(_0720_),
    .A2(_0721_));
 sg13g2_a21oi_1 _3264_ (.A1(_0702_),
    .A2(_0707_),
    .Y(_0724_),
    .B1(_0700_));
 sg13g2_a21oi_1 _3265_ (.A1(_0720_),
    .A2(_0724_),
    .Y(_0725_),
    .B1(_0645_));
 sg13g2_o21ai_1 _3266_ (.B1(_0725_),
    .Y(_0726_),
    .A1(_0720_),
    .A2(_0724_));
 sg13g2_and2_1 _3267_ (.A(_0723_),
    .B(_0726_),
    .X(_0727_));
 sg13g2_nand2b_1 _3268_ (.Y(_0728_),
    .B(_0717_),
    .A_N(_0705_));
 sg13g2_a21oi_1 _3269_ (.A1(_0705_),
    .A2(_0718_),
    .Y(_0729_),
    .B1(net789));
 sg13g2_nand2_2 _3270_ (.Y(_0730_),
    .A(_0728_),
    .B(_0729_));
 sg13g2_a21oi_1 _3271_ (.A1(_0727_),
    .A2(_0730_),
    .Y(_0731_),
    .B1(\cpu_instance.mem_instance.addr[24] ));
 sg13g2_o21ai_1 _3272_ (.B1(net749),
    .Y(_0732_),
    .A1(_0716_),
    .A2(_0731_));
 sg13g2_a22oi_1 _3273_ (.Y(_0733_),
    .B1(net743),
    .B2(net441),
    .A2(net838),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ));
 sg13g2_a21oi_1 _3274_ (.A1(_0732_),
    .A2(net442),
    .Y(_0066_),
    .B1(net824));
 sg13g2_nand2_1 _3275_ (.Y(_0734_),
    .A(net811),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ));
 sg13g2_o21ai_1 _3276_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_1582_),
    .A2(net811));
 sg13g2_nand2_1 _3277_ (.Y(_0736_),
    .A(net689),
    .B(_0735_));
 sg13g2_nand2_1 _3278_ (.Y(_0737_),
    .A(_0411_),
    .B(_0735_));
 sg13g2_xnor2_1 _3279_ (.Y(_0738_),
    .A(net689),
    .B(_0735_));
 sg13g2_nand2_1 _3280_ (.Y(_0739_),
    .A(net687),
    .B(_0717_));
 sg13g2_o21ai_1 _3281_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0720_),
    .A2(_0724_));
 sg13g2_nand2b_1 _3282_ (.Y(_0741_),
    .B(_0738_),
    .A_N(_0740_));
 sg13g2_nand2b_1 _3283_ (.Y(_0742_),
    .B(_0740_),
    .A_N(_0738_));
 sg13g2_nand3_1 _3284_ (.B(_0741_),
    .C(_0742_),
    .A(_0644_),
    .Y(_0743_));
 sg13g2_nand2b_1 _3285_ (.Y(_0744_),
    .B(_0735_),
    .A_N(_0728_));
 sg13g2_nand2b_1 _3286_ (.Y(_0745_),
    .B(_0728_),
    .A_N(_0735_));
 sg13g2_nand3_1 _3287_ (.B(_0744_),
    .C(_0745_),
    .A(_1666_),
    .Y(_0746_));
 sg13g2_a22oi_1 _3288_ (.Y(_0747_),
    .B1(_0717_),
    .B2(net699),
    .A2(_0698_),
    .A1(_0439_));
 sg13g2_o21ai_1 _3289_ (.B1(_0747_),
    .Y(_0748_),
    .A1(_0702_),
    .A2(_0703_));
 sg13g2_a21o_1 _3290_ (.A2(_0748_),
    .A1(_0719_),
    .B1(_0738_),
    .X(_0749_));
 sg13g2_nand3_1 _3291_ (.B(_0738_),
    .C(_0748_),
    .A(_0719_),
    .Y(_0750_));
 sg13g2_nand3_1 _3292_ (.B(_0749_),
    .C(_0750_),
    .A(net780),
    .Y(_0751_));
 sg13g2_nand3_1 _3293_ (.B(_0746_),
    .C(_0751_),
    .A(_0743_),
    .Y(_0752_));
 sg13g2_a22oi_1 _3294_ (.Y(_0753_),
    .B1(_0752_),
    .B2(_1584_),
    .A2(_0655_),
    .A1(_0411_));
 sg13g2_a22oi_1 _3295_ (.Y(_0754_),
    .B1(net743),
    .B2(net650),
    .A2(net838),
    .A1(net422));
 sg13g2_o21ai_1 _3296_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0633_),
    .A2(_0753_));
 sg13g2_and2_1 _3297_ (.A(net872),
    .B(_0755_),
    .X(_0067_));
 sg13g2_or2_1 _3298_ (.X(_0756_),
    .B(net691),
    .A(net841));
 sg13g2_nor2_1 _3299_ (.A(_0656_),
    .B(net681),
    .Y(_0757_));
 sg13g2_nor2_1 _3300_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ),
    .B(net811),
    .Y(_0758_));
 sg13g2_a21oi_2 _3301_ (.B1(_0758_),
    .Y(_0759_),
    .A2(_1589_),
    .A1(net811));
 sg13g2_inv_1 _3302_ (.Y(_0760_),
    .A(_0759_));
 sg13g2_nor2_1 _3303_ (.A(net691),
    .B(_0759_),
    .Y(_0761_));
 sg13g2_xnor2_1 _3304_ (.Y(_0762_),
    .A(net693),
    .B(_0760_));
 sg13g2_inv_1 _3305_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_a21oi_1 _3306_ (.A1(_0736_),
    .A2(_0742_),
    .Y(_0764_),
    .B1(_0763_));
 sg13g2_nand3_1 _3307_ (.B(_0742_),
    .C(_0763_),
    .A(_0736_),
    .Y(_0765_));
 sg13g2_nor2_1 _3308_ (.A(_0645_),
    .B(_0764_),
    .Y(_0766_));
 sg13g2_nand2b_2 _3309_ (.Y(_0767_),
    .B(_0759_),
    .A_N(_0744_));
 sg13g2_xnor2_1 _3310_ (.Y(_0768_),
    .A(_0744_),
    .B(_0759_));
 sg13g2_inv_2 _3311_ (.Y(_0769_),
    .A(_0768_));
 sg13g2_nand3_1 _3312_ (.B(_0750_),
    .C(_0762_),
    .A(_0737_),
    .Y(_0770_));
 sg13g2_a21o_2 _3313_ (.A2(_0750_),
    .A1(_0737_),
    .B1(_0762_),
    .X(_0771_));
 sg13g2_nand3_1 _3314_ (.B(_0770_),
    .C(_0771_),
    .A(net780),
    .Y(_0772_));
 sg13g2_o21ai_1 _3315_ (.B1(_0772_),
    .Y(_0773_),
    .A1(net789),
    .A2(_0769_));
 sg13g2_a21oi_2 _3316_ (.B1(_0773_),
    .Y(_0774_),
    .A2(_0766_),
    .A1(_0765_));
 sg13g2_a22oi_1 _3317_ (.Y(_0775_),
    .B1(net749),
    .B2(_0774_),
    .A2(net837),
    .A1(_1588_));
 sg13g2_o21ai_1 _3318_ (.B1(net875),
    .Y(_0776_),
    .A1(_0757_),
    .A2(_0775_));
 sg13g2_a21oi_1 _3319_ (.A1(_1589_),
    .A2(net743),
    .Y(_0068_),
    .B1(_0776_));
 sg13g2_nor2_1 _3320_ (.A(net802),
    .B(_1588_),
    .Y(_0777_));
 sg13g2_a21oi_2 _3321_ (.B1(_0777_),
    .Y(_0778_),
    .A2(net802),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ));
 sg13g2_nor2_1 _3322_ (.A(_0736_),
    .B(_0761_),
    .Y(_0779_));
 sg13g2_nor2b_1 _3323_ (.A(_0738_),
    .B_N(_0762_),
    .Y(_0780_));
 sg13g2_a221oi_1 _3324_ (.B2(_0740_),
    .C1(_0779_),
    .B1(_0780_),
    .A1(net691),
    .Y(_0781_),
    .A2(_0759_));
 sg13g2_nand2_1 _3325_ (.Y(_0782_),
    .A(net761),
    .B(_0781_));
 sg13g2_xnor2_1 _3326_ (.Y(_0783_),
    .A(_0778_),
    .B(_0781_));
 sg13g2_nand2b_2 _3327_ (.Y(_0784_),
    .B(_0759_),
    .A_N(net691));
 sg13g2_nand3_1 _3328_ (.B(net761),
    .C(_0784_),
    .A(_0771_),
    .Y(_0785_));
 sg13g2_a21oi_1 _3329_ (.A1(_0771_),
    .A2(_0784_),
    .Y(_0786_),
    .B1(net761));
 sg13g2_nand2_1 _3330_ (.Y(_0787_),
    .A(net780),
    .B(_0785_));
 sg13g2_or2_1 _3331_ (.X(_0788_),
    .B(net761),
    .A(_0767_));
 sg13g2_a21oi_1 _3332_ (.A1(_0767_),
    .A2(net761),
    .Y(_0789_),
    .B1(net789));
 sg13g2_a22oi_1 _3333_ (.Y(_0790_),
    .B1(_0788_),
    .B2(_0789_),
    .A2(_0783_),
    .A1(net779));
 sg13g2_o21ai_1 _3334_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_0786_),
    .A2(_0787_));
 sg13g2_nand2_1 _3335_ (.Y(_0792_),
    .A(net749),
    .B(_0791_));
 sg13g2_a22oi_1 _3336_ (.Y(_0793_),
    .B1(net742),
    .B2(net366),
    .A2(net840),
    .A1(net364));
 sg13g2_a21oi_1 _3337_ (.A1(_0792_),
    .A2(_0793_),
    .Y(_0069_),
    .B1(net822));
 sg13g2_nor2b_1 _3338_ (.A(net810),
    .B_N(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ),
    .Y(_0794_));
 sg13g2_a21oi_2 _3339_ (.B1(_0794_),
    .Y(_0795_),
    .A2(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ),
    .A1(net810));
 sg13g2_a21o_2 _3340_ (.A2(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ),
    .A1(net810),
    .B1(_0794_),
    .X(_0796_));
 sg13g2_nand3_1 _3341_ (.B(_0781_),
    .C(_0795_),
    .A(net761),
    .Y(_0797_));
 sg13g2_xnor2_1 _3342_ (.Y(_0798_),
    .A(_0782_),
    .B(_0796_));
 sg13g2_nand2b_1 _3343_ (.Y(_0799_),
    .B(_0796_),
    .A_N(net761));
 sg13g2_a21oi_2 _3344_ (.B1(_0799_),
    .Y(_0800_),
    .A2(_0784_),
    .A1(_0771_));
 sg13g2_nor2_1 _3345_ (.A(_0640_),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_o21ai_1 _3346_ (.B1(_0801_),
    .Y(_0802_),
    .A1(_0786_),
    .A2(_0796_));
 sg13g2_nand2b_2 _3347_ (.Y(_0803_),
    .B(_0796_),
    .A_N(_0788_));
 sg13g2_a21oi_1 _3348_ (.A1(_0788_),
    .A2(_0795_),
    .Y(_0804_),
    .B1(net789));
 sg13g2_a22oi_1 _3349_ (.Y(_0805_),
    .B1(_0803_),
    .B2(_0804_),
    .A2(_0798_),
    .A1(net779));
 sg13g2_nand2_1 _3350_ (.Y(_0806_),
    .A(_0802_),
    .B(_0805_));
 sg13g2_nand2_1 _3351_ (.Y(_0807_),
    .A(net364),
    .B(net742));
 sg13g2_a22oi_1 _3352_ (.Y(_0808_),
    .B1(net749),
    .B2(_0806_),
    .A2(net840),
    .A1(net361));
 sg13g2_a21oi_1 _3353_ (.A1(_0807_),
    .A2(_0808_),
    .Y(_0070_),
    .B1(net823));
 sg13g2_nor2b_1 _3354_ (.A(net810),
    .B_N(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][10] ),
    .Y(_0809_));
 sg13g2_a21oi_2 _3355_ (.B1(_0809_),
    .Y(_0810_),
    .A2(net361),
    .A1(net810));
 sg13g2_a21o_2 _3356_ (.A2(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ),
    .A1(net809),
    .B1(_0809_),
    .X(_0811_));
 sg13g2_nor2_1 _3357_ (.A(_0800_),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_a21o_1 _3358_ (.A2(_0811_),
    .A1(_0800_),
    .B1(_0640_),
    .X(_0813_));
 sg13g2_xnor2_1 _3359_ (.Y(_0814_),
    .A(_0803_),
    .B(_0811_));
 sg13g2_xnor2_1 _3360_ (.Y(_0815_),
    .A(_0797_),
    .B(_0811_));
 sg13g2_or3_1 _3361_ (.A(_0645_),
    .B(_0797_),
    .C(_0811_),
    .X(_0816_));
 sg13g2_a22oi_1 _3362_ (.Y(_0817_),
    .B1(_0815_),
    .B2(net779),
    .A2(_0814_),
    .A1(_1666_));
 sg13g2_o21ai_1 _3363_ (.B1(_0817_),
    .Y(_0818_),
    .A1(_0812_),
    .A2(_0813_));
 sg13g2_nand2_1 _3364_ (.Y(_0819_),
    .A(net749),
    .B(_0818_));
 sg13g2_a22oi_1 _3365_ (.Y(_0820_),
    .B1(net742),
    .B2(net361),
    .A2(net840),
    .A1(net603));
 sg13g2_a21oi_1 _3366_ (.A1(_0819_),
    .A2(_0820_),
    .Y(_0071_),
    .B1(net823));
 sg13g2_o21ai_1 _3367_ (.B1(net779),
    .Y(_0821_),
    .A1(_0797_),
    .A2(_0811_));
 sg13g2_nor2b_1 _3368_ (.A(net809),
    .B_N(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ),
    .Y(_0822_));
 sg13g2_a21oi_2 _3369_ (.B1(_0822_),
    .Y(_0823_),
    .A2(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ),
    .A1(net809));
 sg13g2_a21o_2 _3370_ (.A2(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ),
    .A1(net809),
    .B1(_0822_),
    .X(_0824_));
 sg13g2_nand3_1 _3371_ (.B(_0821_),
    .C(_0824_),
    .A(_0813_),
    .Y(_0825_));
 sg13g2_nand3_1 _3372_ (.B(_0800_),
    .C(_0811_),
    .A(net780),
    .Y(_0826_));
 sg13g2_nand3_1 _3373_ (.B(_0823_),
    .C(_0826_),
    .A(_0816_),
    .Y(_0827_));
 sg13g2_o21ai_1 _3374_ (.B1(_0823_),
    .Y(_0828_),
    .A1(_0803_),
    .A2(_0810_));
 sg13g2_nand3b_1 _3375_ (.B(_0811_),
    .C(_0824_),
    .Y(_0829_),
    .A_N(_0799_));
 sg13g2_nor4_1 _3376_ (.A(_0767_),
    .B(_0799_),
    .C(_0810_),
    .D(_0823_),
    .Y(_0830_));
 sg13g2_nor2_1 _3377_ (.A(net789),
    .B(_0830_),
    .Y(_0831_));
 sg13g2_a22oi_1 _3378_ (.Y(_0832_),
    .B1(_0828_),
    .B2(_0831_),
    .A2(_0827_),
    .A1(_0825_));
 sg13g2_a22oi_1 _3379_ (.Y(_0833_),
    .B1(net742),
    .B2(net603),
    .A2(net836),
    .A1(net549));
 sg13g2_o21ai_1 _3380_ (.B1(_0833_),
    .Y(_0834_),
    .A1(_0633_),
    .A2(_0832_));
 sg13g2_and2_1 _3381_ (.A(net872),
    .B(_0834_),
    .X(_0072_));
 sg13g2_and2_1 _3382_ (.A(net809),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ),
    .X(_0835_));
 sg13g2_a21oi_1 _3383_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ),
    .A2(net802),
    .Y(_0836_),
    .B1(_0835_));
 sg13g2_and4_2 _3384_ (.A(net761),
    .B(_0795_),
    .C(_0810_),
    .D(_0823_),
    .X(_0837_));
 sg13g2_nand3_1 _3385_ (.B(net778),
    .C(_0837_),
    .A(_0781_),
    .Y(_0838_));
 sg13g2_a21o_1 _3386_ (.A2(_0837_),
    .A1(_0781_),
    .B1(net777),
    .X(_0839_));
 sg13g2_a21o_1 _3387_ (.A2(_0839_),
    .A1(_0838_),
    .B1(_0645_),
    .X(_0840_));
 sg13g2_o21ai_1 _3388_ (.B1(net777),
    .Y(_0841_),
    .A1(_0767_),
    .A2(_0829_));
 sg13g2_nand2b_1 _3389_ (.Y(_0842_),
    .B(_0830_),
    .A_N(net778));
 sg13g2_nand3_1 _3390_ (.B(_0841_),
    .C(_0842_),
    .A(_1666_),
    .Y(_0843_));
 sg13g2_a21oi_2 _3391_ (.B1(_0829_),
    .Y(_0844_),
    .A2(_0784_),
    .A1(_0771_));
 sg13g2_nand2b_1 _3392_ (.Y(_0845_),
    .B(_0844_),
    .A_N(net777));
 sg13g2_nand2b_1 _3393_ (.Y(_0846_),
    .B(net777),
    .A_N(_0844_));
 sg13g2_nand3_1 _3394_ (.B(_0845_),
    .C(_0846_),
    .A(net780),
    .Y(_0847_));
 sg13g2_nand3_1 _3395_ (.B(_0843_),
    .C(_0847_),
    .A(_0840_),
    .Y(_0848_));
 sg13g2_nand2_1 _3396_ (.Y(_0849_),
    .A(net749),
    .B(_0848_));
 sg13g2_a22oi_1 _3397_ (.Y(_0850_),
    .B1(net742),
    .B2(net549),
    .A2(net836),
    .A1(net401));
 sg13g2_a21oi_1 _3398_ (.A1(_0849_),
    .A2(_0850_),
    .Y(_0073_),
    .B1(net822));
 sg13g2_and2_1 _3399_ (.A(net809),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ),
    .X(_0851_));
 sg13g2_a21oi_2 _3400_ (.B1(_0851_),
    .Y(_0852_),
    .A2(net802),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ));
 sg13g2_inv_1 _3401_ (.Y(_0853_),
    .A(_0852_));
 sg13g2_nand4_1 _3402_ (.B(net777),
    .C(_0837_),
    .A(_0781_),
    .Y(_0854_),
    .D(_0852_));
 sg13g2_xnor2_1 _3403_ (.Y(_0855_),
    .A(_0838_),
    .B(_0853_));
 sg13g2_nor2_1 _3404_ (.A(net777),
    .B(_0852_),
    .Y(_0856_));
 sg13g2_a221oi_1 _3405_ (.B2(_0844_),
    .C1(_0640_),
    .B1(_0856_),
    .A1(_0845_),
    .Y(_0857_),
    .A2(_0852_));
 sg13g2_nand2_1 _3406_ (.Y(_0858_),
    .A(_0842_),
    .B(_0852_));
 sg13g2_nor4_1 _3407_ (.A(_0767_),
    .B(_0829_),
    .C(net777),
    .D(_0852_),
    .Y(_0859_));
 sg13g2_nor2_1 _3408_ (.A(net789),
    .B(_0859_),
    .Y(_0860_));
 sg13g2_a22oi_1 _3409_ (.Y(_0861_),
    .B1(_0858_),
    .B2(_0860_),
    .A2(_0855_),
    .A1(net779));
 sg13g2_nand2b_1 _3410_ (.Y(_0862_),
    .B(_0861_),
    .A_N(_0857_));
 sg13g2_nand2_1 _3411_ (.Y(_0863_),
    .A(net749),
    .B(_0862_));
 sg13g2_a22oi_1 _3412_ (.Y(_0864_),
    .B1(net742),
    .B2(net401),
    .A2(net836),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ));
 sg13g2_a21oi_1 _3413_ (.A1(_0863_),
    .A2(net402),
    .Y(_0074_),
    .B1(net822));
 sg13g2_mux2_2 _3414_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ),
    .S(net809),
    .X(_0865_));
 sg13g2_a21oi_1 _3415_ (.A1(_0844_),
    .A2(_0856_),
    .Y(_0866_),
    .B1(net793));
 sg13g2_nand3_1 _3416_ (.B(_0856_),
    .C(net793),
    .A(_0844_),
    .Y(_0867_));
 sg13g2_nor2b_1 _3417_ (.A(_0866_),
    .B_N(_0867_),
    .Y(_0868_));
 sg13g2_nand3_1 _3418_ (.B(_0854_),
    .C(net793),
    .A(net779),
    .Y(_0869_));
 sg13g2_nor2_1 _3419_ (.A(_0853_),
    .B(net793),
    .Y(_0870_));
 sg13g2_nor2_1 _3420_ (.A(_0854_),
    .B(net793),
    .Y(_0871_));
 sg13g2_nand4_1 _3421_ (.B(net777),
    .C(_0837_),
    .A(_0781_),
    .Y(_0872_),
    .D(_0870_));
 sg13g2_o21ai_1 _3422_ (.B1(_1666_),
    .Y(_0873_),
    .A1(_0859_),
    .A2(net793));
 sg13g2_nand3b_1 _3423_ (.B(_0853_),
    .C(net793),
    .Y(_0874_),
    .A_N(_0842_));
 sg13g2_inv_1 _3424_ (.Y(_0875_),
    .A(_0874_));
 sg13g2_o21ai_1 _3425_ (.B1(_0869_),
    .Y(_0876_),
    .A1(_0873_),
    .A2(_0875_));
 sg13g2_a221oi_1 _3426_ (.B2(net779),
    .C1(_0876_),
    .B1(_0871_),
    .A1(net780),
    .Y(_0877_),
    .A2(_0868_));
 sg13g2_a22oi_1 _3427_ (.Y(_0878_),
    .B1(net742),
    .B2(net664),
    .A2(net836),
    .A1(net423));
 sg13g2_o21ai_1 _3428_ (.B1(_0878_),
    .Y(_0879_),
    .A1(_0633_),
    .A2(_0877_));
 sg13g2_and2_1 _3429_ (.A(net872),
    .B(_0879_),
    .X(_0075_));
 sg13g2_nand4_1 _3430_ (.B(_0844_),
    .C(_0856_),
    .A(net780),
    .Y(_0880_),
    .D(net793));
 sg13g2_and2_1 _3431_ (.A(net809),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ),
    .X(_0881_));
 sg13g2_a21oi_2 _3432_ (.B1(_0881_),
    .Y(_0882_),
    .A2(net802),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ));
 sg13g2_o21ai_1 _3433_ (.B1(_0882_),
    .Y(_0883_),
    .A1(_0645_),
    .A2(_0872_));
 sg13g2_nor2b_1 _3434_ (.A(_0883_),
    .B_N(_0880_),
    .Y(_0884_));
 sg13g2_a221oi_1 _3435_ (.B2(net779),
    .C1(_0882_),
    .B1(_0872_),
    .A1(net780),
    .Y(_0885_),
    .A2(_0867_));
 sg13g2_a21oi_1 _3436_ (.A1(_0874_),
    .A2(_0882_),
    .Y(_0886_),
    .B1(net789));
 sg13g2_o21ai_1 _3437_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0874_),
    .A2(_0882_));
 sg13g2_o21ai_1 _3438_ (.B1(_0887_),
    .Y(_0888_),
    .A1(_0884_),
    .A2(_0885_));
 sg13g2_nand2_1 _3439_ (.Y(_0889_),
    .A(net749),
    .B(_0888_));
 sg13g2_a22oi_1 _3440_ (.Y(_0890_),
    .B1(net742),
    .B2(net423),
    .A2(net837),
    .A1(net415));
 sg13g2_a21oi_1 _3441_ (.A1(_0889_),
    .A2(_0890_),
    .Y(_0076_),
    .B1(net823));
 sg13g2_nand2b_2 _3442_ (.Y(_0891_),
    .B(_1650_),
    .A_N(net763));
 sg13g2_and2_2 _3443_ (.A(net806),
    .B(_1633_),
    .X(_0892_));
 sg13g2_nand2_2 _3444_ (.Y(_0893_),
    .A(net806),
    .B(_1633_));
 sg13g2_nand2_1 _3445_ (.Y(_0894_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ),
    .B(net796));
 sg13g2_a21oi_1 _3446_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ),
    .A2(net796),
    .Y(_0895_),
    .B1(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ));
 sg13g2_nor2_1 _3447_ (.A(net429),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ),
    .Y(_0896_));
 sg13g2_nor3_2 _3448_ (.A(net384),
    .B(net429),
    .C(net553),
    .Y(_0897_));
 sg13g2_nand2_2 _3449_ (.Y(_0898_),
    .A(_1587_),
    .B(_0896_));
 sg13g2_and2_1 _3450_ (.A(_0025_),
    .B(net796),
    .X(_0899_));
 sg13g2_nand2_1 _3451_ (.Y(_0900_),
    .A(net807),
    .B(net795));
 sg13g2_o21ai_1 _3452_ (.B1(net795),
    .Y(_0901_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ),
    .A2(_0025_));
 sg13g2_nor2_1 _3453_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .Y(_0902_));
 sg13g2_nor2_1 _3454_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_a21oi_2 _3455_ (.B1(_0903_),
    .Y(_0904_),
    .A2(_0901_),
    .A1(_0024_));
 sg13g2_nand2_1 _3456_ (.Y(_0905_),
    .A(_0897_),
    .B(_0904_));
 sg13g2_nand2_1 _3457_ (.Y(_0906_),
    .A(net806),
    .B(_1648_));
 sg13g2_a21oi_1 _3458_ (.A1(_0894_),
    .A2(_0906_),
    .Y(_0907_),
    .B1(_0905_));
 sg13g2_nand2b_1 _3459_ (.Y(_0908_),
    .B(_0907_),
    .A_N(_0895_));
 sg13g2_o21ai_1 _3460_ (.B1(_1609_),
    .Y(_0909_),
    .A1(_0905_),
    .A2(_0906_));
 sg13g2_a21oi_1 _3461_ (.A1(_0908_),
    .A2(_0909_),
    .Y(_0910_),
    .B1(net776));
 sg13g2_o21ai_1 _3462_ (.B1(net776),
    .Y(_0911_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .A2(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ));
 sg13g2_nor4_1 _3463_ (.A(net804),
    .B(net665),
    .C(net659),
    .D(_0893_),
    .Y(_0912_));
 sg13g2_a21oi_1 _3464_ (.A1(net467),
    .A2(_0912_),
    .Y(_0913_),
    .B1(_0891_));
 sg13g2_o21ai_1 _3465_ (.B1(_0913_),
    .Y(_0914_),
    .A1(net567),
    .A2(_0911_));
 sg13g2_nor2_1 _3466_ (.A(_0910_),
    .B(_0914_),
    .Y(_0915_));
 sg13g2_a21oi_1 _3467_ (.A1(_1609_),
    .A2(_0891_),
    .Y(_0077_),
    .B1(_0915_));
 sg13g2_nand2_1 _3468_ (.Y(_0916_),
    .A(net388),
    .B(_0907_));
 sg13g2_nand3b_1 _3469_ (.B(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .C(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ),
    .Y(_0917_),
    .A_N(_0907_));
 sg13g2_nor2b_1 _3470_ (.A(_0891_),
    .B_N(_0917_),
    .Y(_0918_));
 sg13g2_a22oi_1 _3471_ (.Y(_0078_),
    .B1(_0916_),
    .B2(_0918_),
    .A2(_0891_),
    .A1(_1610_));
 sg13g2_nor4_1 _3472_ (.A(net804),
    .B(net659),
    .C(_1628_),
    .D(_0905_),
    .Y(_0919_));
 sg13g2_nor2_1 _3473_ (.A(_0912_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nor2_1 _3474_ (.A(_0891_),
    .B(_0920_),
    .Y(_0079_));
 sg13g2_a21oi_2 _3475_ (.B1(_1651_),
    .Y(_0921_),
    .A2(_1608_),
    .A1(_1585_));
 sg13g2_nor2_1 _3476_ (.A(_1650_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_nor3_1 _3477_ (.A(_1649_),
    .B(net776),
    .C(_0904_),
    .Y(_0923_));
 sg13g2_or2_1 _3478_ (.X(_0924_),
    .B(_0923_),
    .A(_0922_));
 sg13g2_nand2_2 _3479_ (.Y(_0925_),
    .A(_0893_),
    .B(_0897_));
 sg13g2_nor3_1 _3480_ (.A(net805),
    .B(net795),
    .C(_0925_),
    .Y(_0926_));
 sg13g2_nor3_1 _3481_ (.A(net806),
    .B(net805),
    .C(_0898_),
    .Y(_0927_));
 sg13g2_nor3_2 _3482_ (.A(net776),
    .B(_0924_),
    .C(_0927_),
    .Y(_0928_));
 sg13g2_and2_1 _3483_ (.A(_1650_),
    .B(_0928_),
    .X(_0929_));
 sg13g2_and2_1 _3484_ (.A(net553),
    .B(_0929_),
    .X(_0930_));
 sg13g2_nor2_1 _3485_ (.A(net553),
    .B(_0928_),
    .Y(_0931_));
 sg13g2_nor3_1 _3486_ (.A(net762),
    .B(_0930_),
    .C(_0931_),
    .Y(_0080_));
 sg13g2_a21oi_1 _3487_ (.A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .A2(net801),
    .Y(_0932_),
    .B1(_1641_));
 sg13g2_nand2b_1 _3488_ (.Y(_0933_),
    .B(_1628_),
    .A_N(_1639_));
 sg13g2_o21ai_1 _3489_ (.B1(_1587_),
    .Y(_0934_),
    .A1(_0932_),
    .A2(_0933_));
 sg13g2_nand3_1 _3490_ (.B(_0929_),
    .C(_0934_),
    .A(_0896_),
    .Y(_0935_));
 sg13g2_nand2b_1 _3491_ (.Y(_0936_),
    .B(_0928_),
    .A_N(_0930_));
 sg13g2_nand2_1 _3492_ (.Y(_0937_),
    .A(net429),
    .B(_0936_));
 sg13g2_a21oi_1 _3493_ (.A1(_0935_),
    .A2(_0937_),
    .Y(_0081_),
    .B1(net762));
 sg13g2_o21ai_1 _3494_ (.B1(_0928_),
    .Y(_0938_),
    .A1(net790),
    .A2(_0896_));
 sg13g2_nor3_2 _3495_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ),
    .B(_1632_),
    .C(_0898_),
    .Y(_0939_));
 sg13g2_a21o_1 _3496_ (.A2(net790),
    .A1(net815),
    .B1(_0939_),
    .X(_0940_));
 sg13g2_a22oi_1 _3497_ (.Y(_0941_),
    .B1(_0940_),
    .B2(_0928_),
    .A2(_0938_),
    .A1(net384));
 sg13g2_nor2_1 _3498_ (.A(net762),
    .B(net385),
    .Y(_0082_));
 sg13g2_nand3_1 _3499_ (.B(_1629_),
    .C(_0897_),
    .A(net803),
    .Y(_0942_));
 sg13g2_nor3_1 _3500_ (.A(net763),
    .B(_0904_),
    .C(_0942_),
    .Y(_0083_));
 sg13g2_and4_2 _3501_ (.A(_1586_),
    .B(_1609_),
    .C(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .D(net776),
    .X(_0943_));
 sg13g2_mux2_1 _3502_ (.A0(net334),
    .A1(net8),
    .S(_0943_),
    .X(_0084_));
 sg13g2_mux2_1 _3503_ (.A0(net349),
    .A1(net9),
    .S(_0943_),
    .X(_0085_));
 sg13g2_mux2_1 _3504_ (.A0(net337),
    .A1(net10),
    .S(_0943_),
    .X(_0086_));
 sg13g2_mux2_1 _3505_ (.A0(net338),
    .A1(net11),
    .S(_0943_),
    .X(_0087_));
 sg13g2_and4_1 _3506_ (.A(_1650_),
    .B(_0893_),
    .C(_0898_),
    .D(_0904_),
    .X(_0944_));
 sg13g2_a21oi_1 _3507_ (.A1(_0900_),
    .A2(_0944_),
    .Y(_0945_),
    .B1(_0924_));
 sg13g2_and2_2 _3508_ (.A(_0911_),
    .B(_0945_),
    .X(_0946_));
 sg13g2_a21oi_1 _3509_ (.A1(_0016_),
    .A2(_1641_),
    .Y(_0947_),
    .B1(_0932_));
 sg13g2_a21oi_1 _3510_ (.A1(_0015_),
    .A2(net795),
    .Y(_0948_),
    .B1(_0925_));
 sg13g2_o21ai_1 _3511_ (.B1(_0948_),
    .Y(_0949_),
    .A1(net795),
    .A2(_0947_));
 sg13g2_nand2_1 _3512_ (.Y(_0950_),
    .A(_1650_),
    .B(_0949_));
 sg13g2_o21ai_1 _3513_ (.B1(_0950_),
    .Y(_0951_),
    .A1(_1584_),
    .A2(_1650_));
 sg13g2_mux2_1 _3514_ (.A0(net808),
    .A1(_0951_),
    .S(_0946_),
    .X(_0952_));
 sg13g2_nor2b_1 _3515_ (.A(net762),
    .B_N(_0952_),
    .Y(_0088_));
 sg13g2_o21ai_1 _3516_ (.B1(net805),
    .Y(_0953_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .A2(net803));
 sg13g2_and2_1 _3517_ (.A(_1633_),
    .B(_0953_),
    .X(_0954_));
 sg13g2_or3_1 _3518_ (.A(net795),
    .B(_1631_),
    .C(_0954_),
    .X(_0955_));
 sg13g2_nand3_1 _3519_ (.B(net388),
    .C(net776),
    .A(_1586_),
    .Y(_0956_));
 sg13g2_a22oi_1 _3520_ (.Y(_0957_),
    .B1(_0948_),
    .B2(_0955_),
    .A2(net790),
    .A1(net815));
 sg13g2_nand3_1 _3521_ (.B(_0956_),
    .C(_0957_),
    .A(_0946_),
    .Y(_0958_));
 sg13g2_o21ai_1 _3522_ (.B1(_0958_),
    .Y(_0959_),
    .A1(net807),
    .A2(_0946_));
 sg13g2_nor2_1 _3523_ (.A(net763),
    .B(_0959_),
    .Y(_0089_));
 sg13g2_a21oi_1 _3524_ (.A1(net807),
    .A2(net808),
    .Y(_0960_),
    .B1(net805));
 sg13g2_nor3_1 _3525_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .B(net803),
    .C(net808),
    .Y(_0961_));
 sg13g2_nor2_1 _3526_ (.A(_1639_),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_nor4_1 _3527_ (.A(net795),
    .B(_0925_),
    .C(_0960_),
    .D(_0962_),
    .Y(_0963_));
 sg13g2_o21ai_1 _3528_ (.B1(_0946_),
    .Y(_0964_),
    .A1(net790),
    .A2(_0963_));
 sg13g2_o21ai_1 _3529_ (.B1(_0964_),
    .Y(_0965_),
    .A1(net806),
    .A2(_0946_));
 sg13g2_nor2_1 _3530_ (.A(net763),
    .B(_0965_),
    .Y(_0090_));
 sg13g2_nand2_2 _3531_ (.Y(_0966_),
    .A(net790),
    .B(_0921_));
 sg13g2_a21oi_1 _3532_ (.A1(net790),
    .A2(_0921_),
    .Y(_0967_),
    .B1(net803));
 sg13g2_a21oi_1 _3533_ (.A1(net802),
    .A2(_1607_),
    .Y(_0968_),
    .B1(_0966_));
 sg13g2_nor3_1 _3534_ (.A(net762),
    .B(_0967_),
    .C(_0968_),
    .Y(_0091_));
 sg13g2_a22oi_1 _3535_ (.Y(_0969_),
    .B1(_0966_),
    .B2(net326),
    .A2(_1652_),
    .A1(net815));
 sg13g2_nand2b_1 _3536_ (.Y(_0092_),
    .B(_0969_),
    .A_N(net762));
 sg13g2_a21oi_1 _3537_ (.A1(net627),
    .A2(_0966_),
    .Y(_0970_),
    .B1(net762));
 sg13g2_o21ai_1 _3538_ (.B1(_0970_),
    .Y(_0093_),
    .A1(_1584_),
    .A2(_0966_));
 sg13g2_a21oi_1 _3539_ (.A1(_1650_),
    .A2(_0893_),
    .Y(_0971_),
    .B1(net399));
 sg13g2_nor2b_1 _3540_ (.A(_0922_),
    .B_N(net399),
    .Y(_0972_));
 sg13g2_nor3_1 _3541_ (.A(net763),
    .B(_0971_),
    .C(_0972_),
    .Y(_0094_));
 sg13g2_o21ai_1 _3542_ (.B1(_0025_),
    .Y(_0973_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .A2(net803));
 sg13g2_a21oi_1 _3543_ (.A1(_1640_),
    .A2(_0973_),
    .Y(_0974_),
    .B1(net795));
 sg13g2_nor2_1 _3544_ (.A(_0925_),
    .B(_0974_),
    .Y(_0975_));
 sg13g2_o21ai_1 _3545_ (.B1(_0904_),
    .Y(_0976_),
    .A1(_0939_),
    .A2(_0975_));
 sg13g2_nor2_1 _3546_ (.A(_0926_),
    .B(_0944_),
    .Y(_0977_));
 sg13g2_nand3_1 _3547_ (.B(_0976_),
    .C(_0977_),
    .A(_0928_),
    .Y(_0978_));
 sg13g2_mux2_1 _3548_ (.A0(net790),
    .A1(net638),
    .S(_0978_),
    .X(_0979_));
 sg13g2_nor2b_1 _3549_ (.A(net763),
    .B_N(_0979_),
    .Y(_0095_));
 sg13g2_nor2_2 _3550_ (.A(_0892_),
    .B(_0897_),
    .Y(_0980_));
 sg13g2_nand3_1 _3551_ (.B(_1630_),
    .C(_0980_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .Y(_0981_));
 sg13g2_a21oi_1 _3552_ (.A1(_0024_),
    .A2(_0893_),
    .Y(_0982_),
    .B1(_0025_));
 sg13g2_a22oi_1 _3553_ (.Y(_0983_),
    .B1(_0981_),
    .B2(_0982_),
    .A2(_0902_),
    .A1(_0899_));
 sg13g2_and2_2 _3554_ (.A(_1629_),
    .B(_0902_),
    .X(_0984_));
 sg13g2_nand2b_1 _3555_ (.Y(_0985_),
    .B(net334),
    .A_N(_0984_));
 sg13g2_a21oi_1 _3556_ (.A1(net8),
    .A2(_0984_),
    .Y(_0986_),
    .B1(net804));
 sg13g2_o21ai_1 _3557_ (.B1(\cpu_instance.ctrl_instance.scan_in ),
    .Y(_0987_),
    .A1(_0892_),
    .A2(_0897_));
 sg13g2_a21oi_1 _3558_ (.A1(net8),
    .A2(_0980_),
    .Y(_0988_),
    .B1(net801));
 sg13g2_a22oi_1 _3559_ (.Y(_0989_),
    .B1(_0987_),
    .B2(_0988_),
    .A2(_0986_),
    .A1(_0985_));
 sg13g2_mux2_1 _3560_ (.A0(_0989_),
    .A1(net461),
    .S(net745),
    .X(_0096_));
 sg13g2_nand2b_1 _3561_ (.Y(_0990_),
    .B(net349),
    .A_N(_0984_));
 sg13g2_a21oi_1 _3562_ (.A1(net9),
    .A2(_0984_),
    .Y(_0991_),
    .B1(net803));
 sg13g2_o21ai_1 _3563_ (.B1(net432),
    .Y(_0992_),
    .A1(_0892_),
    .A2(_0897_));
 sg13g2_a21oi_1 _3564_ (.A1(net9),
    .A2(_0980_),
    .Y(_0993_),
    .B1(net801));
 sg13g2_a22oi_1 _3565_ (.Y(_0994_),
    .B1(_0992_),
    .B2(_0993_),
    .A2(_0991_),
    .A1(_0990_));
 sg13g2_mux2_1 _3566_ (.A0(_0994_),
    .A1(net517),
    .S(net746),
    .X(_0097_));
 sg13g2_nand2b_1 _3567_ (.Y(_0995_),
    .B(net337),
    .A_N(_0984_));
 sg13g2_a21oi_1 _3568_ (.A1(net10),
    .A2(_0984_),
    .Y(_0996_),
    .B1(net803));
 sg13g2_o21ai_1 _3569_ (.B1(net420),
    .Y(_0997_),
    .A1(net776),
    .A2(_0897_));
 sg13g2_a21oi_1 _3570_ (.A1(net10),
    .A2(_0980_),
    .Y(_0998_),
    .B1(net801));
 sg13g2_a22oi_1 _3571_ (.Y(_0999_),
    .B1(_0997_),
    .B2(_0998_),
    .A2(_0996_),
    .A1(_0995_));
 sg13g2_mux2_1 _3572_ (.A0(_0999_),
    .A1(net511),
    .S(net746),
    .X(_0098_));
 sg13g2_nand2b_1 _3573_ (.Y(_1000_),
    .B(net338),
    .A_N(_0984_));
 sg13g2_a21oi_1 _3574_ (.A1(net11),
    .A2(_0984_),
    .Y(_1001_),
    .B1(net803));
 sg13g2_o21ai_1 _3575_ (.B1(net450),
    .Y(_1002_),
    .A1(net776),
    .A2(_0897_));
 sg13g2_a21oi_1 _3576_ (.A1(net11),
    .A2(_0980_),
    .Y(_1003_),
    .B1(net801));
 sg13g2_a22oi_1 _3577_ (.Y(_1004_),
    .B1(_1002_),
    .B2(_1003_),
    .A2(_1001_),
    .A1(_1000_));
 sg13g2_mux2_1 _3578_ (.A0(_1004_),
    .A1(net599),
    .S(net746),
    .X(_0099_));
 sg13g2_nor2_2 _3579_ (.A(net801),
    .B(_0980_),
    .Y(_1005_));
 sg13g2_nor2b_1 _3580_ (.A(_1005_),
    .B_N(net461),
    .Y(_1006_));
 sg13g2_a21oi_1 _3581_ (.A1(net424),
    .A2(_1005_),
    .Y(_1007_),
    .B1(_1006_));
 sg13g2_nand2_1 _3582_ (.Y(_1008_),
    .A(net484),
    .B(net745));
 sg13g2_o21ai_1 _3583_ (.B1(_1008_),
    .Y(_0100_),
    .A1(net745),
    .A2(_1007_));
 sg13g2_nor2b_1 _3584_ (.A(_1005_),
    .B_N(\cpu_instance.mem_instance.data_qo_mi[1] ),
    .Y(_1009_));
 sg13g2_a21oi_1 _3585_ (.A1(net443),
    .A2(_1005_),
    .Y(_1010_),
    .B1(_1009_));
 sg13g2_nand2_1 _3586_ (.Y(_1011_),
    .A(net446),
    .B(net745));
 sg13g2_o21ai_1 _3587_ (.B1(_1011_),
    .Y(_0101_),
    .A1(net746),
    .A2(_1010_));
 sg13g2_mux2_1 _3588_ (.A0(net511),
    .A1(net396),
    .S(_1005_),
    .X(_1012_));
 sg13g2_nor2_1 _3589_ (.A(net745),
    .B(_1012_),
    .Y(_1013_));
 sg13g2_a21oi_1 _3590_ (.A1(_1626_),
    .A2(net745),
    .Y(_0102_),
    .B1(_1013_));
 sg13g2_nor2b_1 _3591_ (.A(_1005_),
    .B_N(\cpu_instance.mem_instance.data_qo_mi[3] ),
    .Y(_1014_));
 sg13g2_a21oi_1 _3592_ (.A1(net372),
    .A2(_1005_),
    .Y(_1015_),
    .B1(_1014_));
 sg13g2_nand2_1 _3593_ (.Y(_1016_),
    .A(net518),
    .B(net745));
 sg13g2_o21ai_1 _3594_ (.B1(_1016_),
    .Y(_0103_),
    .A1(net745),
    .A2(_1015_));
 sg13g2_nand2b_1 _3595_ (.Y(_0104_),
    .B(net895),
    .A_N(net326));
 sg13g2_nand2_1 _3596_ (.Y(_1017_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ));
 sg13g2_nand2b_1 _3597_ (.Y(_1018_),
    .B(\cpu_instance.mem_ctrl_op[1] ),
    .A_N(\cpu_instance.mem_ctrl_op[0] ));
 sg13g2_nor2_1 _3598_ (.A(_1017_),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_nor3_2 _3599_ (.A(\cpu_instance.mem_instance.data_req ),
    .B(_1017_),
    .C(_1018_),
    .Y(_1020_));
 sg13g2_nor2b_1 _3600_ (.A(net581),
    .B_N(\cpu_instance.mem_ctrl_op[0] ),
    .Y(_1021_));
 sg13g2_nand2b_2 _3601_ (.Y(_1022_),
    .B(\cpu_instance.mem_ctrl_op[0] ),
    .A_N(\cpu_instance.mem_ctrl_op[1] ));
 sg13g2_nand2_1 _3602_ (.Y(_1023_),
    .A(_1017_),
    .B(_1021_));
 sg13g2_nor2_1 _3603_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .Y(_1024_));
 sg13g2_nor3_1 _3604_ (.A(net857),
    .B(_1020_),
    .C(_1024_),
    .Y(_1025_));
 sg13g2_a22oi_1 _3605_ (.Y(_1026_),
    .B1(_1023_),
    .B2(_1025_),
    .A2(net659),
    .A1(net854));
 sg13g2_nor2_1 _3606_ (.A(net825),
    .B(_1026_),
    .Y(_0105_));
 sg13g2_mux2_1 _3607_ (.A0(net8),
    .A1(net467),
    .S(net896),
    .X(_0106_));
 sg13g2_mux2_1 _3608_ (.A0(net9),
    .A1(net388),
    .S(net896),
    .X(_0107_));
 sg13g2_a22oi_1 _3609_ (.Y(_1027_),
    .B1(net766),
    .B2(net770),
    .A2(net759),
    .A1(net333));
 sg13g2_inv_1 _3610_ (.Y(_0108_),
    .A(_1027_));
 sg13g2_a22oi_1 _3611_ (.Y(_1028_),
    .B1(_0635_),
    .B2(net769),
    .A2(net760),
    .A1(net330));
 sg13g2_inv_1 _3612_ (.Y(_0109_),
    .A(_1028_));
 sg13g2_a22oi_1 _3613_ (.Y(_1029_),
    .B1(_0661_),
    .B2(net770),
    .A2(net760),
    .A1(net331));
 sg13g2_inv_1 _3614_ (.Y(_0110_),
    .A(_1029_));
 sg13g2_a22oi_1 _3615_ (.Y(_1030_),
    .B1(_0679_),
    .B2(net769),
    .A2(net759),
    .A1(net329));
 sg13g2_inv_1 _3616_ (.Y(_0111_),
    .A(_1030_));
 sg13g2_nor2_1 _3617_ (.A(net342),
    .B(_1655_),
    .Y(_1031_));
 sg13g2_nor2_1 _3618_ (.A(_1653_),
    .B(_0698_),
    .Y(_1032_));
 sg13g2_nor2_1 _3619_ (.A(net333),
    .B(_1647_),
    .Y(_1033_));
 sg13g2_nor3_1 _3620_ (.A(_1031_),
    .B(_1032_),
    .C(_1033_),
    .Y(_0112_));
 sg13g2_nor2_1 _3621_ (.A(net330),
    .B(_1647_),
    .Y(_1034_));
 sg13g2_a221oi_1 _3622_ (.B2(net769),
    .C1(_1034_),
    .B1(_0718_),
    .A1(_1620_),
    .Y(_0113_),
    .A2(net759));
 sg13g2_nor2_1 _3623_ (.A(net357),
    .B(_1655_),
    .Y(_1035_));
 sg13g2_nor2_1 _3624_ (.A(net331),
    .B(_1647_),
    .Y(_1036_));
 sg13g2_nor2_1 _3625_ (.A(_1653_),
    .B(_0735_),
    .Y(_1037_));
 sg13g2_nor3_1 _3626_ (.A(_1035_),
    .B(_1036_),
    .C(_1037_),
    .Y(_0114_));
 sg13g2_nor2_1 _3627_ (.A(net329),
    .B(_1647_),
    .Y(_1038_));
 sg13g2_a221oi_1 _3628_ (.B2(net770),
    .C1(_1038_),
    .B1(_0760_),
    .A1(_1621_),
    .Y(_0115_),
    .A2(net759));
 sg13g2_nor2_1 _3629_ (.A(net342),
    .B(_1647_),
    .Y(_1039_));
 sg13g2_a221oi_1 _3630_ (.B2(net769),
    .C1(_1039_),
    .B1(_0778_),
    .A1(_1622_),
    .Y(_0116_),
    .A2(net759));
 sg13g2_nor2_1 _3631_ (.A(_1653_),
    .B(_0796_),
    .Y(_1040_));
 sg13g2_a221oi_1 _3632_ (.B2(_1623_),
    .C1(_1040_),
    .B1(net759),
    .A1(_1620_),
    .Y(_0117_),
    .A2(net772));
 sg13g2_nor2_1 _3633_ (.A(net357),
    .B(_1647_),
    .Y(_1041_));
 sg13g2_a221oi_1 _3634_ (.B2(net769),
    .C1(_1041_),
    .B1(net362),
    .A1(_1624_),
    .Y(_0118_),
    .A2(net759));
 sg13g2_nor2_1 _3635_ (.A(_1653_),
    .B(_0824_),
    .Y(_1042_));
 sg13g2_a221oi_1 _3636_ (.B2(_1625_),
    .C1(_1042_),
    .B1(net759),
    .A1(_1621_),
    .Y(_0119_),
    .A2(net772));
 sg13g2_nor2_1 _3637_ (.A(net352),
    .B(_1655_),
    .Y(_1043_));
 sg13g2_a221oi_1 _3638_ (.B2(net778),
    .C1(_1043_),
    .B1(net769),
    .A1(_1622_),
    .Y(_0120_),
    .A2(net772));
 sg13g2_nor2_1 _3639_ (.A(net323),
    .B(_1655_),
    .Y(_1044_));
 sg13g2_a221oi_1 _3640_ (.B2(_0852_),
    .C1(_1044_),
    .B1(net769),
    .A1(_1623_),
    .Y(_0121_),
    .A2(net772));
 sg13g2_or2_1 _3641_ (.X(_1045_),
    .B(_0865_),
    .A(_1653_));
 sg13g2_o21ai_1 _3642_ (.B1(_1045_),
    .Y(_1046_),
    .A1(net320),
    .A2(_1655_));
 sg13g2_a21oi_1 _3643_ (.A1(_1624_),
    .A2(net772),
    .Y(_0122_),
    .B1(_1046_));
 sg13g2_nor2_1 _3644_ (.A(net312),
    .B(_1655_),
    .Y(_1047_));
 sg13g2_a221oi_1 _3645_ (.B2(net351),
    .C1(_1047_),
    .B1(net769),
    .A1(_1625_),
    .Y(_0123_),
    .A2(net772));
 sg13g2_nor2b_1 _3646_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ),
    .B_N(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .Y(_1048_));
 sg13g2_o21ai_1 _3647_ (.B1(net895),
    .Y(_1049_),
    .A1(net854),
    .A2(_1048_));
 sg13g2_a21oi_1 _3648_ (.A1(net854),
    .A2(_1606_),
    .Y(_0124_),
    .B1(_1049_));
 sg13g2_nand2b_1 _3649_ (.Y(_1050_),
    .B(_1024_),
    .A_N(_1018_));
 sg13g2_and2_1 _3650_ (.A(net833),
    .B(_1050_),
    .X(_1051_));
 sg13g2_nand2b_1 _3651_ (.Y(_1052_),
    .B(net895),
    .A_N(_1051_));
 sg13g2_a21oi_1 _3652_ (.A1(net854),
    .A2(_1607_),
    .Y(_0125_),
    .B1(net756));
 sg13g2_o21ai_1 _3653_ (.B1(net897),
    .Y(_1053_),
    .A1(net833),
    .A2(net651));
 sg13g2_a21oi_1 _3654_ (.A1(_1021_),
    .A2(_1024_),
    .Y(_1054_),
    .B1(net854));
 sg13g2_nor2_1 _3655_ (.A(_1053_),
    .B(_1054_),
    .Y(_0126_));
 sg13g2_nand2_1 _3656_ (.Y(_1055_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ),
    .B(\cpu_instance.mem_instance.data_ready ));
 sg13g2_nor2_1 _3657_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .B(_1055_),
    .Y(_1056_));
 sg13g2_o21ai_1 _3658_ (.B1(net833),
    .Y(_1057_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .A2(_1055_));
 sg13g2_nor2_1 _3659_ (.A(\cpu_instance.mem_instance.addr[24] ),
    .B(_1022_),
    .Y(_1058_));
 sg13g2_and3_1 _3660_ (.X(_1059_),
    .A(net778),
    .B(_0882_),
    .C(_1058_));
 sg13g2_nand3_1 _3661_ (.B(_0870_),
    .C(_1059_),
    .A(_0837_),
    .Y(_1060_));
 sg13g2_nor4_1 _3662_ (.A(_0679_),
    .B(_0698_),
    .C(_0717_),
    .D(_0735_),
    .Y(_1061_));
 sg13g2_nor2_1 _3663_ (.A(_0760_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_nor4_2 _3664_ (.A(_0692_),
    .B(_0769_),
    .C(_1060_),
    .Y(_1063_),
    .D(_1062_));
 sg13g2_a221oi_1 _3665_ (.B2(_1063_),
    .C1(_1057_),
    .B1(_1024_),
    .A1(net576),
    .Y(_1064_),
    .A2(_1019_));
 sg13g2_o21ai_1 _3666_ (.B1(net895),
    .Y(_1065_),
    .A1(net833),
    .A2(net647));
 sg13g2_nor2_1 _3667_ (.A(_1064_),
    .B(_1065_),
    .Y(_0127_));
 sg13g2_a221oi_1 _3668_ (.B2(_1050_),
    .C1(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .B1(_1022_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ),
    .Y(_1066_),
    .A2(\cpu_instance.mem_instance.data_ready ));
 sg13g2_nor2_1 _3669_ (.A(_1020_),
    .B(_1066_),
    .Y(_1067_));
 sg13g2_nor2b_1 _3670_ (.A(_1022_),
    .B_N(_1048_),
    .Y(_1068_));
 sg13g2_nor3_1 _3671_ (.A(_1020_),
    .B(_1056_),
    .C(_1068_),
    .Y(_1069_));
 sg13g2_and2_1 _3672_ (.A(_1050_),
    .B(_1069_),
    .X(_1070_));
 sg13g2_nor4_2 _3673_ (.A(_1614_),
    .B(_1020_),
    .C(_1066_),
    .Y(_1071_),
    .D(_1070_));
 sg13g2_nand2_1 _3674_ (.Y(_1072_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ),
    .B(_0768_));
 sg13g2_nor2_2 _3675_ (.A(_0652_),
    .B(_0769_),
    .Y(_1073_));
 sg13g2_nor2b_1 _3676_ (.A(net744),
    .B_N(_1063_),
    .Y(_1074_));
 sg13g2_nand2b_2 _3677_ (.Y(_1075_),
    .B(_1063_),
    .A_N(net744));
 sg13g2_mux2_1 _3678_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ),
    .S(net766),
    .X(_1076_));
 sg13g2_nand2_1 _3679_ (.Y(_1077_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .B(net766));
 sg13g2_nand2_1 _3680_ (.Y(_1078_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .B(_1672_));
 sg13g2_a21oi_1 _3681_ (.A1(_1077_),
    .A2(_1078_),
    .Y(_1079_),
    .B1(_0769_));
 sg13g2_a22oi_1 _3682_ (.Y(_1080_),
    .B1(_1079_),
    .B2(_0652_),
    .A2(_1076_),
    .A1(_1073_));
 sg13g2_o21ai_1 _3683_ (.B1(_0768_),
    .Y(_1081_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ),
    .A2(net765));
 sg13g2_a21oi_1 _3684_ (.A1(_1570_),
    .A2(net765),
    .Y(_1082_),
    .B1(_1081_));
 sg13g2_a21oi_1 _3685_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ),
    .A2(_0768_),
    .Y(_1083_),
    .B1(_1672_));
 sg13g2_a21oi_1 _3686_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .A2(_0768_),
    .Y(_1084_),
    .B1(net765));
 sg13g2_or2_1 _3687_ (.X(_1085_),
    .B(_1084_),
    .A(_1083_));
 sg13g2_a21oi_1 _3688_ (.A1(_0651_),
    .A2(_1085_),
    .Y(_1086_),
    .B1(_0668_));
 sg13g2_o21ai_1 _3689_ (.B1(_1086_),
    .Y(_1087_),
    .A1(_0651_),
    .A2(_1082_));
 sg13g2_o21ai_1 _3690_ (.B1(_1087_),
    .Y(_1088_),
    .A1(net747),
    .A2(_1080_));
 sg13g2_a221oi_1 _3691_ (.B2(_1088_),
    .C1(net858),
    .B1(_1074_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[0] ),
    .Y(_1089_),
    .A2(_1071_));
 sg13g2_nor2_1 _3692_ (.A(net854),
    .B(_1067_),
    .Y(_1090_));
 sg13g2_nor2_1 _3693_ (.A(net854),
    .B(_1070_),
    .Y(_1091_));
 sg13g2_a21oi_1 _3694_ (.A1(_1614_),
    .A2(_1091_),
    .Y(_1092_),
    .B1(_1090_));
 sg13g2_nor2_1 _3695_ (.A(_1063_),
    .B(_1092_),
    .Y(_1093_));
 sg13g2_or2_1 _3696_ (.X(_1094_),
    .B(_1092_),
    .A(_1063_));
 sg13g2_nor2_1 _3697_ (.A(net564),
    .B(net834),
    .Y(_1095_));
 sg13g2_nand2_1 _3698_ (.Y(_1096_),
    .A(net669),
    .B(_1093_));
 sg13g2_o21ai_1 _3699_ (.B1(_1096_),
    .Y(_1097_),
    .A1(_1089_),
    .A2(_1095_));
 sg13g2_and2_1 _3700_ (.A(net897),
    .B(_1097_),
    .X(_0128_));
 sg13g2_nand2_1 _3701_ (.Y(_1098_),
    .A(net517),
    .B(_1071_));
 sg13g2_a21oi_1 _3702_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ),
    .A2(_0768_),
    .Y(_1099_),
    .B1(_0650_));
 sg13g2_mux2_1 _3703_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .S(net765),
    .X(_1100_));
 sg13g2_nand2_1 _3704_ (.Y(_1101_),
    .A(_0768_),
    .B(_1100_));
 sg13g2_a221oi_1 _3705_ (.B2(_0651_),
    .C1(_1099_),
    .B1(_1101_),
    .A1(_0648_),
    .Y(_1102_),
    .A2(_1072_));
 sg13g2_mux2_1 _3706_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .S(net765),
    .X(_1103_));
 sg13g2_nor2_2 _3707_ (.A(_0651_),
    .B(_0769_),
    .Y(_1104_));
 sg13g2_mux2_1 _3708_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .S(net765),
    .X(_1105_));
 sg13g2_a22oi_1 _3709_ (.Y(_1106_),
    .B1(_1105_),
    .B2(_1073_),
    .A2(_1104_),
    .A1(_1103_));
 sg13g2_a21oi_1 _3710_ (.A1(_0668_),
    .A2(_1106_),
    .Y(_1107_),
    .B1(_1075_));
 sg13g2_o21ai_1 _3711_ (.B1(_1107_),
    .Y(_1108_),
    .A1(_0668_),
    .A2(_1102_));
 sg13g2_a21oi_1 _3712_ (.A1(_1098_),
    .A2(_1108_),
    .Y(_1109_),
    .B1(net858));
 sg13g2_a21oi_1 _3713_ (.A1(net597),
    .A2(net859),
    .Y(_1110_),
    .B1(_1109_));
 sg13g2_o21ai_1 _3714_ (.B1(net897),
    .Y(_1111_),
    .A1(net564),
    .A2(net707));
 sg13g2_a21oi_1 _3715_ (.A1(net707),
    .A2(_1110_),
    .Y(_0129_),
    .B1(_1111_));
 sg13g2_nor2_1 _3716_ (.A(net610),
    .B(net834),
    .Y(_1112_));
 sg13g2_mux2_1 _3717_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .S(net765),
    .X(_1113_));
 sg13g2_a22oi_1 _3718_ (.Y(_1114_),
    .B1(_1113_),
    .B2(_1073_),
    .A2(_1104_),
    .A1(_1076_));
 sg13g2_a21oi_1 _3719_ (.A1(_0652_),
    .A2(_1085_),
    .Y(_1115_),
    .B1(_0668_));
 sg13g2_o21ai_1 _3720_ (.B1(_1115_),
    .Y(_1116_),
    .A1(_0652_),
    .A2(_1079_));
 sg13g2_o21ai_1 _3721_ (.B1(_1116_),
    .Y(_1117_),
    .A1(net747),
    .A2(_1114_));
 sg13g2_a221oi_1 _3722_ (.B2(_1117_),
    .C1(net858),
    .B1(_1074_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[2] ),
    .Y(_1118_),
    .A2(net744));
 sg13g2_o21ai_1 _3723_ (.B1(net707),
    .Y(_1119_),
    .A1(_1112_),
    .A2(_1118_));
 sg13g2_o21ai_1 _3724_ (.B1(net897),
    .Y(_1120_),
    .A1(net597),
    .A2(net707));
 sg13g2_nor2b_1 _3725_ (.A(_1120_),
    .B_N(_1119_),
    .Y(_0130_));
 sg13g2_a21oi_1 _3726_ (.A1(_1073_),
    .A2(_1103_),
    .Y(_1121_),
    .B1(_0668_));
 sg13g2_o21ai_1 _3727_ (.B1(_1121_),
    .Y(_1122_),
    .A1(_0651_),
    .A2(_1101_));
 sg13g2_mux2_1 _3728_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .S(net767),
    .X(_1123_));
 sg13g2_mux2_1 _3729_ (.A0(_1105_),
    .A1(_1123_),
    .S(_0651_),
    .X(_1124_));
 sg13g2_a21oi_1 _3730_ (.A1(_0768_),
    .A2(_1124_),
    .Y(_1125_),
    .B1(net748));
 sg13g2_nor2_2 _3731_ (.A(_1075_),
    .B(_1125_),
    .Y(_1126_));
 sg13g2_a22oi_1 _3732_ (.Y(_1127_),
    .B1(_1122_),
    .B2(_1126_),
    .A2(net744),
    .A1(\cpu_instance.mem_instance.data_qo_mi[3] ));
 sg13g2_or2_1 _3733_ (.X(_1128_),
    .B(_1127_),
    .A(net856));
 sg13g2_a21oi_1 _3734_ (.A1(net570),
    .A2(net859),
    .Y(_1129_),
    .B1(_1093_));
 sg13g2_o21ai_1 _3735_ (.B1(net895),
    .Y(_1130_),
    .A1(\cpu_instance.mem_instance.bus_data_out[3] ),
    .A2(net707));
 sg13g2_a21oi_1 _3736_ (.A1(_1128_),
    .A2(_1129_),
    .Y(_0131_),
    .B1(_1130_));
 sg13g2_mux2_1 _3737_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ),
    .S(net767),
    .X(_1131_));
 sg13g2_a22oi_1 _3738_ (.Y(_1132_),
    .B1(_1131_),
    .B2(_1073_),
    .A2(_1113_),
    .A1(_1104_));
 sg13g2_nand2_2 _3739_ (.Y(_1133_),
    .A(_0668_),
    .B(_1132_));
 sg13g2_a21oi_2 _3740_ (.B1(_1075_),
    .Y(_1134_),
    .A2(_1080_),
    .A1(net747));
 sg13g2_a22oi_1 _3741_ (.Y(_1135_),
    .B1(_1133_),
    .B2(_1134_),
    .A2(net744),
    .A1(net484));
 sg13g2_a21oi_1 _3742_ (.A1(net575),
    .A2(net858),
    .Y(_1136_),
    .B1(_1093_));
 sg13g2_o21ai_1 _3743_ (.B1(_1136_),
    .Y(_1137_),
    .A1(net858),
    .A2(_1135_));
 sg13g2_o21ai_1 _3744_ (.B1(_1137_),
    .Y(_1138_),
    .A1(net570),
    .A2(net708));
 sg13g2_nor2_1 _3745_ (.A(net826),
    .B(_1138_),
    .Y(_0132_));
 sg13g2_mux2_1 _3746_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ),
    .S(net767),
    .X(_1139_));
 sg13g2_a221oi_1 _3747_ (.B2(_1073_),
    .C1(net747),
    .B1(_1139_),
    .A1(_1104_),
    .Y(_1140_),
    .A2(_1123_));
 sg13g2_nor2_1 _3748_ (.A(net563),
    .B(net834),
    .Y(_1141_));
 sg13g2_a21oi_2 _3749_ (.B1(_1140_),
    .Y(_1142_),
    .A2(_1106_),
    .A1(net747));
 sg13g2_a221oi_1 _3750_ (.B2(_1142_),
    .C1(net858),
    .B1(_1074_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[5] ),
    .Y(_1143_),
    .A2(net744));
 sg13g2_o21ai_1 _3751_ (.B1(net708),
    .Y(_1144_),
    .A1(_1141_),
    .A2(_1143_));
 sg13g2_o21ai_1 _3752_ (.B1(_1144_),
    .Y(_1145_),
    .A1(net575),
    .A2(net707));
 sg13g2_nor2_1 _3753_ (.A(net826),
    .B(_1145_),
    .Y(_0133_));
 sg13g2_mux2_1 _3754_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .S(net767),
    .X(_1146_));
 sg13g2_a221oi_1 _3755_ (.B2(_1073_),
    .C1(net747),
    .B1(_1146_),
    .A1(_1104_),
    .Y(_1147_),
    .A2(_1131_));
 sg13g2_a21o_1 _3756_ (.A2(_1114_),
    .A1(net747),
    .B1(_1075_),
    .X(_1148_));
 sg13g2_a21oi_1 _3757_ (.A1(net548),
    .A2(net744),
    .Y(_1149_),
    .B1(net858));
 sg13g2_o21ai_1 _3758_ (.B1(_1149_),
    .Y(_1150_),
    .A1(_1147_),
    .A2(_1148_));
 sg13g2_o21ai_1 _3759_ (.B1(_1150_),
    .Y(_1151_),
    .A1(net489),
    .A2(net833));
 sg13g2_o21ai_1 _3760_ (.B1(net895),
    .Y(_1152_),
    .A1(net563),
    .A2(net707));
 sg13g2_a21oi_1 _3761_ (.A1(net707),
    .A2(_1151_),
    .Y(_0134_),
    .B1(_1152_));
 sg13g2_mux2_1 _3762_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .S(net767),
    .X(_1153_));
 sg13g2_nand2_1 _3763_ (.Y(_1154_),
    .A(_0651_),
    .B(_1153_));
 sg13g2_nand2_1 _3764_ (.Y(_1155_),
    .A(_0652_),
    .B(_1139_));
 sg13g2_a21oi_1 _3765_ (.A1(_1154_),
    .A2(_1155_),
    .Y(_1156_),
    .B1(net747));
 sg13g2_a21oi_2 _3766_ (.B1(_1156_),
    .Y(_1157_),
    .A2(_1124_),
    .A1(net748));
 sg13g2_a21oi_1 _3767_ (.A1(\cpu_instance.mem_instance.data_qo_mi[7] ),
    .A2(net744),
    .Y(_1158_),
    .B1(net858));
 sg13g2_o21ai_1 _3768_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_1075_),
    .A2(_1157_));
 sg13g2_o21ai_1 _3769_ (.B1(_1159_),
    .Y(_1160_),
    .A1(net833),
    .A2(net321));
 sg13g2_o21ai_1 _3770_ (.B1(net897),
    .Y(_1161_),
    .A1(net489),
    .A2(net708));
 sg13g2_a21oi_1 _3771_ (.A1(net708),
    .A2(_1160_),
    .Y(_0135_),
    .B1(_1161_));
 sg13g2_a21oi_1 _3772_ (.A1(net854),
    .A2(net613),
    .Y(_1162_),
    .B1(_1090_));
 sg13g2_nor2_1 _3773_ (.A(net825),
    .B(_1162_),
    .Y(_0136_));
 sg13g2_a21oi_1 _3774_ (.A1(net857),
    .A2(_1802_),
    .Y(_1163_),
    .B1(_1091_));
 sg13g2_nor2_1 _3775_ (.A(net825),
    .B(_1163_),
    .Y(_0137_));
 sg13g2_a22oi_1 _3776_ (.Y(_1164_),
    .B1(_0490_),
    .B2(_0593_),
    .A2(net607),
    .A1(net859));
 sg13g2_nor2_1 _3777_ (.A(net828),
    .B(_1164_),
    .Y(_0138_));
 sg13g2_a22oi_1 _3778_ (.Y(_1165_),
    .B1(_0490_),
    .B2(_0600_),
    .A2(net859),
    .A1(net819));
 sg13g2_nor2_1 _3779_ (.A(net828),
    .B(_1165_),
    .Y(_0139_));
 sg13g2_nand2_1 _3780_ (.Y(_1166_),
    .A(net895),
    .B(_1051_));
 sg13g2_a21oi_2 _3781_ (.B1(_1166_),
    .Y(_1167_),
    .A2(_1069_),
    .A1(_1067_));
 sg13g2_or2_2 _3782_ (.X(_1168_),
    .B(net718),
    .A(net865));
 sg13g2_nand2_1 _3783_ (.Y(_1169_),
    .A(net432),
    .B(net860));
 sg13g2_a21oi_1 _3784_ (.A1(net706),
    .A2(_1169_),
    .Y(_1170_),
    .B1(_1052_));
 sg13g2_a21o_1 _3785_ (.A2(_1167_),
    .A1(net500),
    .B1(_1170_),
    .X(_0140_));
 sg13g2_nand2_1 _3786_ (.Y(_1171_),
    .A(net420),
    .B(net860));
 sg13g2_a21oi_1 _3787_ (.A1(net710),
    .A2(_1171_),
    .Y(_1172_),
    .B1(net756));
 sg13g2_a21o_1 _3788_ (.A2(_1167_),
    .A1(net432),
    .B1(_1172_),
    .X(_0141_));
 sg13g2_nand2_2 _3789_ (.Y(_1173_),
    .A(net832),
    .B(_0513_));
 sg13g2_nand2_1 _3790_ (.Y(_1174_),
    .A(\cpu_instance.mem_instance.data_qi_mo[3] ),
    .B(net860));
 sg13g2_a21oi_1 _3791_ (.A1(net698),
    .A2(_1174_),
    .Y(_1175_),
    .B1(net756));
 sg13g2_a21o_1 _3792_ (.A2(_1167_),
    .A1(net420),
    .B1(_1175_),
    .X(_0142_));
 sg13g2_or2_1 _3793_ (.X(_1176_),
    .B(net701),
    .A(net842));
 sg13g2_nand2_1 _3794_ (.Y(_1177_),
    .A(net424),
    .B(net861));
 sg13g2_a21oi_1 _3795_ (.A1(net696),
    .A2(_1177_),
    .Y(_1178_),
    .B1(net756));
 sg13g2_a21o_1 _3796_ (.A2(_1167_),
    .A1(net450),
    .B1(_1178_),
    .X(_0143_));
 sg13g2_nand2_2 _3797_ (.Y(_1179_),
    .A(net832),
    .B(_0439_));
 sg13g2_nand2_1 _3798_ (.Y(_1180_),
    .A(\cpu_instance.mem_instance.data_qi_mo[5] ),
    .B(net860));
 sg13g2_a21oi_1 _3799_ (.A1(net686),
    .A2(_1180_),
    .Y(_1181_),
    .B1(net756));
 sg13g2_a21o_1 _3800_ (.A2(_1167_),
    .A1(net424),
    .B1(_1181_),
    .X(_0144_));
 sg13g2_nand2_1 _3801_ (.Y(_1182_),
    .A(_1603_),
    .B(net699));
 sg13g2_nand2_1 _3802_ (.Y(_1183_),
    .A(net396),
    .B(net860));
 sg13g2_a21oi_1 _3803_ (.A1(net684),
    .A2(_1183_),
    .Y(_1184_),
    .B1(net756));
 sg13g2_a21o_1 _3804_ (.A2(_1167_),
    .A1(net443),
    .B1(_1184_),
    .X(_0145_));
 sg13g2_nand2_2 _3805_ (.Y(_1185_),
    .A(net832),
    .B(_0411_));
 sg13g2_nand2_1 _3806_ (.Y(_1186_),
    .A(net372),
    .B(net860));
 sg13g2_a21oi_1 _3807_ (.A1(net680),
    .A2(_1186_),
    .Y(_1187_),
    .B1(net756));
 sg13g2_a21o_1 _3808_ (.A2(_1167_),
    .A1(net396),
    .B1(_1187_),
    .X(_0146_));
 sg13g2_nand2_1 _3809_ (.Y(_1188_),
    .A(\cpu_instance.mem_instance.bus_data_out[0] ),
    .B(net861));
 sg13g2_a21oi_1 _3810_ (.A1(net682),
    .A2(_1188_),
    .Y(_1189_),
    .B1(net756));
 sg13g2_a21o_1 _3811_ (.A2(_1167_),
    .A1(net372),
    .B1(_1189_),
    .X(_0147_));
 sg13g2_nor2_1 _3812_ (.A(net811),
    .B(_1669_),
    .Y(_1190_));
 sg13g2_nor2_1 _3813_ (.A(net837),
    .B(_1190_),
    .Y(_1191_));
 sg13g2_o21ai_1 _3814_ (.B1(net831),
    .Y(_1192_),
    .A1(net811),
    .A2(_1669_));
 sg13g2_nor2_2 _3815_ (.A(net837),
    .B(_1191_),
    .Y(_1193_));
 sg13g2_o21ai_1 _3816_ (.B1(_1193_),
    .Y(_1194_),
    .A1(net768),
    .A2(net717));
 sg13g2_a221oi_1 _3817_ (.B2(_1664_),
    .C1(_1194_),
    .B1(_1795_),
    .A1(_1666_),
    .Y(_1195_),
    .A2(_1672_));
 sg13g2_o21ai_1 _3818_ (.B1(net872),
    .Y(_1196_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ),
    .A2(net831));
 sg13g2_nor2_1 _3819_ (.A(net415),
    .B(_1192_),
    .Y(_1197_));
 sg13g2_nor3_1 _3820_ (.A(_1195_),
    .B(_1196_),
    .C(_1197_),
    .Y(_0148_));
 sg13g2_nand2_2 _3821_ (.Y(_1198_),
    .A(net831),
    .B(_1668_));
 sg13g2_and2_1 _3822_ (.A(_0653_),
    .B(_1193_),
    .X(_1199_));
 sg13g2_o21ai_1 _3823_ (.B1(_1199_),
    .Y(_1200_),
    .A1(net768),
    .A2(net714));
 sg13g2_o21ai_1 _3824_ (.B1(_1200_),
    .Y(_1201_),
    .A1(net346),
    .A2(net831));
 sg13g2_o21ai_1 _3825_ (.B1(_1201_),
    .Y(_1202_),
    .A1(_0647_),
    .A2(_1198_));
 sg13g2_o21ai_1 _3826_ (.B1(_1202_),
    .Y(_1203_),
    .A1(net637),
    .A2(_1192_));
 sg13g2_nor2_1 _3827_ (.A(net824),
    .B(_1203_),
    .Y(_0149_));
 sg13g2_o21ai_1 _3828_ (.B1(_1193_),
    .Y(_1204_),
    .A1(net768),
    .A2(net712));
 sg13g2_nor2_1 _3829_ (.A(_0673_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_o21ai_1 _3830_ (.B1(net874),
    .Y(_1206_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ),
    .A2(net831));
 sg13g2_nor2_1 _3831_ (.A(net346),
    .B(_1192_),
    .Y(_1207_));
 sg13g2_nor3_1 _3832_ (.A(_1205_),
    .B(_1206_),
    .C(_1207_),
    .Y(_0150_));
 sg13g2_nor2_1 _3833_ (.A(_0689_),
    .B(_1198_),
    .Y(_1208_));
 sg13g2_a22oi_1 _3834_ (.Y(_1209_),
    .B1(_0693_),
    .B2(_1193_),
    .A2(net841),
    .A1(_1583_));
 sg13g2_nor2_1 _3835_ (.A(net768),
    .B(net695),
    .Y(_1210_));
 sg13g2_nor3_1 _3836_ (.A(_1208_),
    .B(_1209_),
    .C(_1210_),
    .Y(_1211_));
 sg13g2_o21ai_1 _3837_ (.B1(net874),
    .Y(_1212_),
    .A1(net498),
    .A2(_1192_));
 sg13g2_nor2_1 _3838_ (.A(_1211_),
    .B(_1212_),
    .Y(_0151_));
 sg13g2_o21ai_1 _3839_ (.B1(_1193_),
    .Y(_1213_),
    .A1(net768),
    .A2(net702));
 sg13g2_nor2_1 _3840_ (.A(_0712_),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_o21ai_1 _3841_ (.B1(net874),
    .Y(_1215_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ),
    .A2(net831));
 sg13g2_nor2_1 _3842_ (.A(net340),
    .B(_1192_),
    .Y(_1216_));
 sg13g2_nor3_1 _3843_ (.A(_1214_),
    .B(_1215_),
    .C(_1216_),
    .Y(_0152_));
 sg13g2_nor2_1 _3844_ (.A(_0727_),
    .B(_1198_),
    .Y(_1217_));
 sg13g2_a22oi_1 _3845_ (.Y(_1218_),
    .B1(_0730_),
    .B2(_1193_),
    .A2(net838),
    .A1(_1582_));
 sg13g2_nor2_1 _3846_ (.A(net768),
    .B(net683),
    .Y(_1219_));
 sg13g2_nor3_1 _3847_ (.A(_1217_),
    .B(_1218_),
    .C(_1219_),
    .Y(_1220_));
 sg13g2_o21ai_1 _3848_ (.B1(net874),
    .Y(_1221_),
    .A1(net547),
    .A2(_1192_));
 sg13g2_nor2_1 _3849_ (.A(_1220_),
    .B(_1221_),
    .Y(_0153_));
 sg13g2_o21ai_1 _3850_ (.B1(_1193_),
    .Y(_1222_),
    .A1(net768),
    .A2(net689));
 sg13g2_nor2_1 _3851_ (.A(_0752_),
    .B(_1222_),
    .Y(_1223_));
 sg13g2_o21ai_1 _3852_ (.B1(net872),
    .Y(_1224_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ),
    .A2(net831));
 sg13g2_nor2_1 _3853_ (.A(net344),
    .B(_1192_),
    .Y(_1225_));
 sg13g2_nor3_1 _3854_ (.A(_1223_),
    .B(_1224_),
    .C(_1225_),
    .Y(_0154_));
 sg13g2_nor2_2 _3855_ (.A(net811),
    .B(_1198_),
    .Y(_1226_));
 sg13g2_inv_1 _3856_ (.Y(_1227_),
    .A(_1226_));
 sg13g2_nand2b_1 _3857_ (.Y(_1228_),
    .B(_1192_),
    .A_N(net681));
 sg13g2_a22oi_1 _3858_ (.Y(_1229_),
    .B1(_1227_),
    .B2(_1228_),
    .A2(_0774_),
    .A1(net768));
 sg13g2_a221oi_1 _3859_ (.B2(net608),
    .C1(_1229_),
    .B1(net741),
    .A1(net522),
    .Y(_1230_),
    .A2(net837));
 sg13g2_nor2_1 _3860_ (.A(net823),
    .B(_1230_),
    .Y(_0155_));
 sg13g2_nand2_1 _3861_ (.Y(_1231_),
    .A(_0791_),
    .B(_1226_));
 sg13g2_a22oi_1 _3862_ (.Y(_1232_),
    .B1(net741),
    .B2(net522),
    .A2(net836),
    .A1(net363));
 sg13g2_a21oi_1 _3863_ (.A1(_1231_),
    .A2(_1232_),
    .Y(_0156_),
    .B1(net822));
 sg13g2_nand2_1 _3864_ (.Y(_1233_),
    .A(net363),
    .B(net741));
 sg13g2_a22oi_1 _3865_ (.Y(_1234_),
    .B1(_0806_),
    .B2(_1226_),
    .A2(net840),
    .A1(net354));
 sg13g2_a21oi_1 _3866_ (.A1(_1233_),
    .A2(_1234_),
    .Y(_0157_),
    .B1(net822));
 sg13g2_nand2_1 _3867_ (.Y(_1235_),
    .A(net354),
    .B(net741));
 sg13g2_a22oi_1 _3868_ (.Y(_1236_),
    .B1(_0818_),
    .B2(_1226_),
    .A2(net836),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ));
 sg13g2_a21oi_1 _3869_ (.A1(_1235_),
    .A2(_1236_),
    .Y(_0158_),
    .B1(net822));
 sg13g2_a22oi_1 _3870_ (.Y(_1237_),
    .B1(net741),
    .B2(net668),
    .A2(net839),
    .A1(net359));
 sg13g2_o21ai_1 _3871_ (.B1(_1237_),
    .Y(_1238_),
    .A1(_0832_),
    .A2(_1227_));
 sg13g2_and2_1 _3872_ (.A(net872),
    .B(_1238_),
    .X(_0159_));
 sg13g2_nand2_1 _3873_ (.Y(_1239_),
    .A(net359),
    .B(net741));
 sg13g2_a22oi_1 _3874_ (.Y(_1240_),
    .B1(_0848_),
    .B2(_1226_),
    .A2(net839),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ));
 sg13g2_a21oi_1 _3875_ (.A1(_1239_),
    .A2(_1240_),
    .Y(_0160_),
    .B1(net822));
 sg13g2_nand2_1 _3876_ (.Y(_1241_),
    .A(_0862_),
    .B(_1226_));
 sg13g2_a22oi_1 _3877_ (.Y(_1242_),
    .B1(net741),
    .B2(net543),
    .A2(net836),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ));
 sg13g2_a21oi_1 _3878_ (.A1(_1241_),
    .A2(net544),
    .Y(_0161_),
    .B1(net822));
 sg13g2_a22oi_1 _3879_ (.Y(_1243_),
    .B1(net741),
    .B2(net640),
    .A2(net836),
    .A1(net350));
 sg13g2_o21ai_1 _3880_ (.B1(_1243_),
    .Y(_1244_),
    .A1(_0877_),
    .A2(_1227_));
 sg13g2_and2_1 _3881_ (.A(net872),
    .B(_1244_),
    .X(_0162_));
 sg13g2_nand2_1 _3882_ (.Y(_1245_),
    .A(_0888_),
    .B(_1226_));
 sg13g2_a22oi_1 _3883_ (.Y(_1246_),
    .B1(_1191_),
    .B2(net350),
    .A2(net837),
    .A1(net540));
 sg13g2_a21oi_1 _3884_ (.A1(_1245_),
    .A2(_1246_),
    .Y(_0163_),
    .B1(net823));
 sg13g2_a22oi_1 _3885_ (.Y(_1247_),
    .B1(net760),
    .B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ),
    .A2(net771),
    .A1(net327));
 sg13g2_inv_1 _3886_ (.Y(_0164_),
    .A(net328));
 sg13g2_nor2_2 _3887_ (.A(\cpu_instance.reg_in_sel[1] ),
    .B(net821),
    .Y(_1248_));
 sg13g2_inv_1 _3888_ (.Y(_1249_),
    .A(_1248_));
 sg13g2_nand2_1 _3889_ (.Y(_1250_),
    .A(net820),
    .B(\cpu_instance.reg_in_sel[0] ));
 sg13g2_nand2b_1 _3890_ (.Y(_1251_),
    .B(_1601_),
    .A_N(_1250_));
 sg13g2_a21oi_1 _3891_ (.A1(_1576_),
    .A2(net821),
    .Y(_1252_),
    .B1(net820));
 sg13g2_a21oi_1 _3892_ (.A1(\cpu_instance.registers_instance.registers[2][3] ),
    .A2(_1595_),
    .Y(_1253_),
    .B1(_1252_));
 sg13g2_a22oi_1 _3893_ (.Y(_1254_),
    .B1(_1251_),
    .B2(_1253_),
    .A2(_1248_),
    .A1(_0020_));
 sg13g2_nor2_1 _3894_ (.A(_1594_),
    .B(net821),
    .Y(_1255_));
 sg13g2_mux4_1 _3895_ (.S0(net821),
    .A0(\cpu_instance.registers_instance.registers[0][2] ),
    .A1(\cpu_instance.registers_instance.registers[1][2] ),
    .A2(\cpu_instance.registers_instance.registers[2][2] ),
    .A3(uo_out[2]),
    .S1(net820),
    .X(_1256_));
 sg13g2_nand2_2 _3896_ (.Y(_1257_),
    .A(_1254_),
    .B(_1256_));
 sg13g2_nand2_2 _3897_ (.Y(_1258_),
    .A(\cpu_instance.ctrl_instance.use_register_bank_in ),
    .B(\cpu_instance.reg_op ));
 sg13g2_nand3_1 _3898_ (.B(net820),
    .C(net821),
    .A(uo_out[1]),
    .Y(_1259_));
 sg13g2_nor2_1 _3899_ (.A(\cpu_instance.reg_in_sel[1] ),
    .B(_1595_),
    .Y(_1260_));
 sg13g2_a221oi_1 _3900_ (.B2(\cpu_instance.registers_instance.registers[1][1] ),
    .C1(_1248_),
    .B1(_1260_),
    .A1(\cpu_instance.registers_instance.registers[2][1] ),
    .Y(_1261_),
    .A2(_1595_));
 sg13g2_a22oi_1 _3901_ (.Y(_1262_),
    .B1(_1259_),
    .B2(_1261_),
    .A2(_1248_),
    .A1(_0019_));
 sg13g2_nand3_1 _3902_ (.B(net820),
    .C(net821),
    .A(uo_out[0]),
    .Y(_1263_));
 sg13g2_a221oi_1 _3903_ (.B2(\cpu_instance.registers_instance.registers[2][0] ),
    .C1(_1248_),
    .B1(_1255_),
    .A1(\cpu_instance.registers_instance.registers[1][0] ),
    .Y(_1264_),
    .A2(_1594_));
 sg13g2_a22oi_1 _3904_ (.Y(_1265_),
    .B1(_1263_),
    .B2(_1264_),
    .A2(_1248_),
    .A1(_0018_));
 sg13g2_nand2_1 _3905_ (.Y(_1266_),
    .A(_1262_),
    .B(_1265_));
 sg13g2_nor3_1 _3906_ (.A(_1257_),
    .B(_1258_),
    .C(_1266_),
    .Y(_1267_));
 sg13g2_o21ai_1 _3907_ (.B1(net886),
    .Y(_1268_),
    .A1(net392),
    .A2(net739));
 sg13g2_a21oi_1 _3908_ (.A1(net718),
    .A2(net739),
    .Y(_0165_),
    .B1(_1268_));
 sg13g2_o21ai_1 _3909_ (.B1(net879),
    .Y(_1269_),
    .A1(net458),
    .A2(net740));
 sg13g2_a21oi_1 _3910_ (.A1(net715),
    .A2(net740),
    .Y(_0166_),
    .B1(_1269_));
 sg13g2_o21ai_1 _3911_ (.B1(net882),
    .Y(_1270_),
    .A1(net368),
    .A2(net739));
 sg13g2_a21oi_1 _3912_ (.A1(net711),
    .A2(net739),
    .Y(_0167_),
    .B1(_1270_));
 sg13g2_o21ai_1 _3913_ (.B1(net881),
    .Y(_1271_),
    .A1(net413),
    .A2(net740));
 sg13g2_a21oi_1 _3914_ (.A1(net701),
    .A2(net740),
    .Y(_0168_),
    .B1(_1271_));
 sg13g2_o21ai_1 _3915_ (.B1(net882),
    .Y(_1272_),
    .A1(net414),
    .A2(net739));
 sg13g2_a21oi_1 _3916_ (.A1(net703),
    .A2(net739),
    .Y(_0169_),
    .B1(_1272_));
 sg13g2_o21ai_1 _3917_ (.B1(net890),
    .Y(_1273_),
    .A1(net463),
    .A2(_1267_));
 sg13g2_a21oi_1 _3918_ (.A1(net688),
    .A2(net740),
    .Y(_0170_),
    .B1(_1273_));
 sg13g2_o21ai_1 _3919_ (.B1(net890),
    .Y(_1274_),
    .A1(net403),
    .A2(net740));
 sg13g2_a21oi_1 _3920_ (.A1(net690),
    .A2(net740),
    .Y(_0171_),
    .B1(_1274_));
 sg13g2_o21ai_1 _3921_ (.B1(net883),
    .Y(_1275_),
    .A1(net437),
    .A2(net739));
 sg13g2_a21oi_1 _3922_ (.A1(net692),
    .A2(net739),
    .Y(_0172_),
    .B1(_1275_));
 sg13g2_nor2b_2 _3923_ (.A(_0022_),
    .B_N(_0548_),
    .Y(_1276_));
 sg13g2_a21oi_2 _3924_ (.B1(_1276_),
    .Y(_1277_),
    .A2(net834),
    .A1(_1599_));
 sg13g2_a21o_2 _3925_ (.A2(net834),
    .A1(_1599_),
    .B1(_1276_),
    .X(_1278_));
 sg13g2_nor3_2 _3926_ (.A(\cpu_instance.ctrl_instance.use_register_bank_in ),
    .B(net867),
    .C(_0022_),
    .Y(_1279_));
 sg13g2_or3_1 _3927_ (.A(\cpu_instance.ctrl_instance.use_register_bank_in ),
    .B(net867),
    .C(_0022_),
    .X(_1280_));
 sg13g2_a21oi_2 _3928_ (.B1(_1278_),
    .Y(_1281_),
    .A2(_1279_),
    .A1(_1249_));
 sg13g2_o21ai_1 _3929_ (.B1(_1277_),
    .Y(_1282_),
    .A1(_1248_),
    .A2(_1280_));
 sg13g2_a21oi_1 _3930_ (.A1(\cpu_instance.registers_instance.registers[0][1] ),
    .A2(net870),
    .Y(_1283_),
    .B1(net755));
 sg13g2_o21ai_1 _3931_ (.B1(net900),
    .Y(_1284_),
    .A1(net520),
    .A2(_1281_));
 sg13g2_a21oi_1 _3932_ (.A1(net706),
    .A2(_1283_),
    .Y(_0173_),
    .B1(_1284_));
 sg13g2_a21oi_1 _3933_ (.A1(net552),
    .A2(net869),
    .Y(_1285_),
    .B1(net755));
 sg13g2_o21ai_1 _3934_ (.B1(net902),
    .Y(_1286_),
    .A1(net624),
    .A2(_1281_));
 sg13g2_a21oi_1 _3935_ (.A1(net710),
    .A2(_1285_),
    .Y(_0174_),
    .B1(_1286_));
 sg13g2_a21oi_1 _3936_ (.A1(net435),
    .A2(net869),
    .Y(_1287_),
    .B1(_1282_));
 sg13g2_a221oi_1 _3937_ (.B2(net698),
    .C1(net827),
    .B1(_1287_),
    .A1(_1581_),
    .Y(_0175_),
    .A2(net755));
 sg13g2_a21oi_1 _3938_ (.A1(\cpu_instance.registers_instance.registers[0][4] ),
    .A2(net869),
    .Y(_1288_),
    .B1(_1282_));
 sg13g2_o21ai_1 _3939_ (.B1(net901),
    .Y(_1289_),
    .A1(net435),
    .A2(_1281_));
 sg13g2_a21oi_1 _3940_ (.A1(net696),
    .A2(_1288_),
    .Y(_0176_),
    .B1(_1289_));
 sg13g2_a21oi_1 _3941_ (.A1(net374),
    .A2(net868),
    .Y(_1290_),
    .B1(net755));
 sg13g2_o21ai_1 _3942_ (.B1(net901),
    .Y(_1291_),
    .A1(net473),
    .A2(_1281_));
 sg13g2_a21oi_1 _3943_ (.A1(net686),
    .A2(_1290_),
    .Y(_0177_),
    .B1(_1291_));
 sg13g2_a21oi_1 _3944_ (.A1(\cpu_instance.registers_instance.registers[0][6] ),
    .A2(net870),
    .Y(_1292_),
    .B1(net755));
 sg13g2_a221oi_1 _3945_ (.B2(net684),
    .C1(net827),
    .B1(_1292_),
    .A1(_1580_),
    .Y(_0178_),
    .A2(net755));
 sg13g2_a21oi_1 _3946_ (.A1(net418),
    .A2(net868),
    .Y(_1293_),
    .B1(net755));
 sg13g2_o21ai_1 _3947_ (.B1(net900),
    .Y(_1294_),
    .A1(net499),
    .A2(_1281_));
 sg13g2_a21oi_1 _3948_ (.A1(net680),
    .A2(_1293_),
    .Y(_0179_),
    .B1(_1294_));
 sg13g2_a21oi_1 _3949_ (.A1(net869),
    .A2(net7),
    .Y(_1295_),
    .B1(net755));
 sg13g2_o21ai_1 _3950_ (.B1(net901),
    .Y(_1296_),
    .A1(net418),
    .A2(_1281_));
 sg13g2_a21oi_1 _3951_ (.A1(net682),
    .A2(_1295_),
    .Y(_0180_),
    .B1(_1296_));
 sg13g2_nor2_1 _3952_ (.A(_1260_),
    .B(_1280_),
    .Y(_1297_));
 sg13g2_nor2_2 _3953_ (.A(_1278_),
    .B(_1297_),
    .Y(_1298_));
 sg13g2_nand2b_1 _3954_ (.Y(_1299_),
    .B(_1277_),
    .A_N(_1297_));
 sg13g2_a21oi_1 _3955_ (.A1(\cpu_instance.registers_instance.registers[1][1] ),
    .A2(net870),
    .Y(_1300_),
    .B1(net753));
 sg13g2_a221oi_1 _3956_ (.B2(net706),
    .C1(net827),
    .B1(_1300_),
    .A1(_1579_),
    .Y(_0181_),
    .A2(net753));
 sg13g2_a21oi_1 _3957_ (.A1(net646),
    .A2(net869),
    .Y(_1301_),
    .B1(net753));
 sg13g2_a221oi_1 _3958_ (.B2(net710),
    .C1(net828),
    .B1(_1301_),
    .A1(_1578_),
    .Y(_0182_),
    .A2(net753));
 sg13g2_a21oi_1 _3959_ (.A1(net587),
    .A2(net869),
    .Y(_1302_),
    .B1(net753));
 sg13g2_a221oi_1 _3960_ (.B2(net698),
    .C1(net828),
    .B1(_1302_),
    .A1(_1577_),
    .Y(_0183_),
    .A2(net753));
 sg13g2_a21oi_1 _3961_ (.A1(net641),
    .A2(net868),
    .Y(_1303_),
    .B1(net754));
 sg13g2_a221oi_1 _3962_ (.B2(net696),
    .C1(net827),
    .B1(_1303_),
    .A1(_1576_),
    .Y(_0184_),
    .A2(net753));
 sg13g2_a21oi_1 _3963_ (.A1(net605),
    .A2(net868),
    .Y(_1304_),
    .B1(net754));
 sg13g2_o21ai_1 _3964_ (.B1(net900),
    .Y(_1305_),
    .A1(\cpu_instance.registers_instance.registers[1][4] ),
    .A2(_1298_));
 sg13g2_a21oi_1 _3965_ (.A1(net686),
    .A2(_1304_),
    .Y(_0185_),
    .B1(_1305_));
 sg13g2_a21oi_1 _3966_ (.A1(net530),
    .A2(net868),
    .Y(_1306_),
    .B1(net754));
 sg13g2_o21ai_1 _3967_ (.B1(net900),
    .Y(_1307_),
    .A1(\cpu_instance.registers_instance.registers[1][5] ),
    .A2(_1298_));
 sg13g2_a21oi_1 _3968_ (.A1(net684),
    .A2(_1306_),
    .Y(_0186_),
    .B1(_1307_));
 sg13g2_a21oi_1 _3969_ (.A1(net559),
    .A2(net870),
    .Y(_1308_),
    .B1(net754));
 sg13g2_o21ai_1 _3970_ (.B1(net900),
    .Y(_1309_),
    .A1(net530),
    .A2(_1298_));
 sg13g2_a21oi_1 _3971_ (.A1(net680),
    .A2(_1308_),
    .Y(_0187_),
    .B1(_1309_));
 sg13g2_a21oi_1 _3972_ (.A1(net520),
    .A2(net870),
    .Y(_1310_),
    .B1(net753));
 sg13g2_o21ai_1 _3973_ (.B1(net900),
    .Y(_1311_),
    .A1(net559),
    .A2(_1298_));
 sg13g2_a21oi_1 _3974_ (.A1(net682),
    .A2(_1310_),
    .Y(_0188_),
    .B1(_1311_));
 sg13g2_nor2_1 _3975_ (.A(_1255_),
    .B(_1280_),
    .Y(_1312_));
 sg13g2_nor2_2 _3976_ (.A(_1278_),
    .B(_1312_),
    .Y(_1313_));
 sg13g2_nand2b_1 _3977_ (.Y(_1314_),
    .B(_1277_),
    .A_N(_1312_));
 sg13g2_a21oi_1 _3978_ (.A1(net579),
    .A2(net867),
    .Y(_1315_),
    .B1(net751));
 sg13g2_a221oi_1 _3979_ (.B2(net706),
    .C1(net827),
    .B1(_1315_),
    .A1(_1575_),
    .Y(_0189_),
    .A2(net751));
 sg13g2_a21oi_1 _3980_ (.A1(net629),
    .A2(net867),
    .Y(_1316_),
    .B1(net751));
 sg13g2_a221oi_1 _3981_ (.B2(net710),
    .C1(net827),
    .B1(_1316_),
    .A1(_1574_),
    .Y(_0190_),
    .A2(net751));
 sg13g2_a21oi_1 _3982_ (.A1(net617),
    .A2(net869),
    .Y(_1317_),
    .B1(net751));
 sg13g2_a221oi_1 _3983_ (.B2(net698),
    .C1(net827),
    .B1(_1317_),
    .A1(_1573_),
    .Y(_0191_),
    .A2(net751));
 sg13g2_a21oi_1 _3984_ (.A1(net601),
    .A2(net870),
    .Y(_1318_),
    .B1(net752));
 sg13g2_a221oi_1 _3985_ (.B2(net696),
    .C1(net827),
    .B1(_1318_),
    .A1(_1572_),
    .Y(_0192_),
    .A2(net751));
 sg13g2_a21oi_1 _3986_ (.A1(net574),
    .A2(net868),
    .Y(_1319_),
    .B1(net752));
 sg13g2_o21ai_1 _3987_ (.B1(net901),
    .Y(_1320_),
    .A1(net601),
    .A2(_1313_));
 sg13g2_a21oi_1 _3988_ (.A1(net686),
    .A2(_1319_),
    .Y(_0193_),
    .B1(_1320_));
 sg13g2_a21oi_1 _3989_ (.A1(net557),
    .A2(net868),
    .Y(_1321_),
    .B1(net752));
 sg13g2_o21ai_1 _3990_ (.B1(net901),
    .Y(_1322_),
    .A1(net574),
    .A2(_1313_));
 sg13g2_a21oi_1 _3991_ (.A1(net684),
    .A2(_1321_),
    .Y(_0194_),
    .B1(_1322_));
 sg13g2_a21oi_1 _3992_ (.A1(\cpu_instance.registers_instance.registers[2][7] ),
    .A2(net868),
    .Y(_1323_),
    .B1(net752));
 sg13g2_o21ai_1 _3993_ (.B1(net900),
    .Y(_1324_),
    .A1(net557),
    .A2(_1313_));
 sg13g2_a21oi_1 _3994_ (.A1(net680),
    .A2(_1323_),
    .Y(_0195_),
    .B1(_1324_));
 sg13g2_a21oi_1 _3995_ (.A1(net318),
    .A2(net870),
    .Y(_1325_),
    .B1(net751));
 sg13g2_o21ai_1 _3996_ (.B1(net900),
    .Y(_1326_),
    .A1(\cpu_instance.registers_instance.registers[2][7] ),
    .A2(_1313_));
 sg13g2_a21oi_1 _3997_ (.A1(net682),
    .A2(_1325_),
    .Y(_0196_),
    .B1(_1326_));
 sg13g2_a21oi_2 _3998_ (.B1(_1278_),
    .Y(_1327_),
    .A2(_1279_),
    .A1(_1250_));
 sg13g2_a21o_1 _3999_ (.A2(_1279_),
    .A1(_1250_),
    .B1(_1278_),
    .X(_1328_));
 sg13g2_a21oi_1 _4000_ (.A1(net653),
    .A2(net866),
    .Y(_1329_),
    .B1(net750));
 sg13g2_o21ai_1 _4001_ (.B1(net899),
    .Y(_1330_),
    .A1(uo_out[0]),
    .A2(_1327_));
 sg13g2_a21oi_1 _4002_ (.A1(net706),
    .A2(_1329_),
    .Y(_0197_),
    .B1(_1330_));
 sg13g2_a21oi_1 _4003_ (.A1(net609),
    .A2(net866),
    .Y(_1331_),
    .B1(_1328_));
 sg13g2_o21ai_1 _4004_ (.B1(net899),
    .Y(_1332_),
    .A1(net653),
    .A2(_1327_));
 sg13g2_a21oi_1 _4005_ (.A1(net710),
    .A2(_1331_),
    .Y(_0198_),
    .B1(_1332_));
 sg13g2_a21oi_1 _4006_ (.A1(net583),
    .A2(net866),
    .Y(_1333_),
    .B1(net750));
 sg13g2_a221oi_1 _4007_ (.B2(net698),
    .C1(net828),
    .B1(_1333_),
    .A1(_1571_),
    .Y(_0199_),
    .A2(net750));
 sg13g2_a21oi_1 _4008_ (.A1(uo_out[4]),
    .A2(net866),
    .Y(_1334_),
    .B1(net750));
 sg13g2_o21ai_1 _4009_ (.B1(net899),
    .Y(_1335_),
    .A1(net583),
    .A2(_1327_));
 sg13g2_a21oi_1 _4010_ (.A1(net696),
    .A2(_1334_),
    .Y(_0200_),
    .B1(_1335_));
 sg13g2_a21oi_1 _4011_ (.A1(net633),
    .A2(net866),
    .Y(_1336_),
    .B1(net750));
 sg13g2_o21ai_1 _4012_ (.B1(net899),
    .Y(_1337_),
    .A1(net648),
    .A2(_1327_));
 sg13g2_a21oi_1 _4013_ (.A1(net686),
    .A2(_1336_),
    .Y(_0201_),
    .B1(_1337_));
 sg13g2_a21oi_1 _4014_ (.A1(net619),
    .A2(net866),
    .Y(_1338_),
    .B1(net750));
 sg13g2_o21ai_1 _4015_ (.B1(net899),
    .Y(_1339_),
    .A1(net633),
    .A2(_1327_));
 sg13g2_a21oi_1 _4016_ (.A1(net684),
    .A2(_1338_),
    .Y(_0202_),
    .B1(_1339_));
 sg13g2_a21oi_1 _4017_ (.A1(uo_out[7]),
    .A2(net866),
    .Y(_1340_),
    .B1(net750));
 sg13g2_o21ai_1 _4018_ (.B1(net902),
    .Y(_1341_),
    .A1(net619),
    .A2(_1327_));
 sg13g2_a21oi_1 _4019_ (.A1(net680),
    .A2(_1340_),
    .Y(_0203_),
    .B1(_1341_));
 sg13g2_a21oi_1 _4020_ (.A1(\cpu_instance.registers_instance.registers[2][0] ),
    .A2(net866),
    .Y(_1342_),
    .B1(net750));
 sg13g2_o21ai_1 _4021_ (.B1(net902),
    .Y(_1343_),
    .A1(net631),
    .A2(_1327_));
 sg13g2_a21oi_1 _4022_ (.A1(net682),
    .A2(_1342_),
    .Y(_0204_),
    .B1(_1343_));
 sg13g2_nor2_1 _4023_ (.A(_1262_),
    .B(_1265_),
    .Y(_1344_));
 sg13g2_nor2_2 _4024_ (.A(_1254_),
    .B(_1256_),
    .Y(_1345_));
 sg13g2_nand2_1 _4025_ (.Y(_1346_),
    .A(_1344_),
    .B(_1345_));
 sg13g2_a21oi_2 _4026_ (.B1(net846),
    .Y(_1347_),
    .A2(\cpu_instance.reg_op ),
    .A1(\cpu_instance.ctrl_instance.use_register_bank_in ));
 sg13g2_a21oi_2 _4027_ (.B1(net791),
    .Y(_1348_),
    .A2(_1346_),
    .A1(net775));
 sg13g2_a21o_2 _4028_ (.A2(_1346_),
    .A1(net775),
    .B1(net791),
    .X(_1349_));
 sg13g2_a21oi_1 _4029_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ),
    .A2(net846),
    .Y(_1350_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4030_ (.B1(net887),
    .Y(_1351_),
    .A1(net568),
    .A2(_1348_));
 sg13g2_a21oi_1 _4031_ (.A1(net705),
    .A2(_1350_),
    .Y(_0205_),
    .B1(_1351_));
 sg13g2_a21oi_1 _4032_ (.A1(net577),
    .A2(net846),
    .Y(_1352_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4033_ (.B1(net887),
    .Y(_1353_),
    .A1(net594),
    .A2(_1348_));
 sg13g2_a21oi_1 _4034_ (.A1(net709),
    .A2(_1352_),
    .Y(_0206_),
    .B1(_1353_));
 sg13g2_a21oi_1 _4035_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .A2(net846),
    .Y(_1354_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4036_ (.B1(net887),
    .Y(_1355_),
    .A1(net577),
    .A2(_1348_));
 sg13g2_a21oi_1 _4037_ (.A1(net697),
    .A2(_1354_),
    .Y(_0207_),
    .B1(_1355_));
 sg13g2_a21oi_1 _4038_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .A2(net846),
    .Y(_1356_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4039_ (.B1(net898),
    .Y(_1357_),
    .A1(net643),
    .A2(_1348_));
 sg13g2_a21oi_1 _4040_ (.A1(net696),
    .A2(_1356_),
    .Y(_0208_),
    .B1(_1357_));
 sg13g2_a21oi_1 _4041_ (.A1(net614),
    .A2(net846),
    .Y(_1358_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4042_ (.B1(net898),
    .Y(_1359_),
    .A1(net649),
    .A2(_1348_));
 sg13g2_a21oi_1 _4043_ (.A1(net685),
    .A2(_1358_),
    .Y(_0209_),
    .B1(_1359_));
 sg13g2_a21oi_1 _4044_ (.A1(net585),
    .A2(net846),
    .Y(_1360_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4045_ (.B1(net898),
    .Y(_1361_),
    .A1(net614),
    .A2(_1348_));
 sg13g2_a21oi_1 _4046_ (.A1(net683),
    .A2(_1360_),
    .Y(_0210_),
    .B1(_1361_));
 sg13g2_a21oi_1 _4047_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .A2(net846),
    .Y(_1362_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4048_ (.B1(net898),
    .Y(_1363_),
    .A1(net585),
    .A2(_1348_));
 sg13g2_a21oi_1 _4049_ (.A1(net679),
    .A2(_1362_),
    .Y(_0211_),
    .B1(_1363_));
 sg13g2_a21oi_1 _4050_ (.A1(uo_out[0]),
    .A2(net865),
    .Y(_1364_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4051_ (.B1(net898),
    .Y(_1365_),
    .A1(net625),
    .A2(_1348_));
 sg13g2_a21oi_1 _4052_ (.A1(net682),
    .A2(_1364_),
    .Y(_0212_),
    .B1(_1365_));
 sg13g2_nor2b_1 _4053_ (.A(_1262_),
    .B_N(_1265_),
    .Y(_1366_));
 sg13g2_nand2b_1 _4054_ (.Y(_1367_),
    .B(_1265_),
    .A_N(_1262_));
 sg13g2_nand2_1 _4055_ (.Y(_1368_),
    .A(_1345_),
    .B(_1366_));
 sg13g2_a21oi_2 _4056_ (.B1(net791),
    .Y(_1369_),
    .A2(_1368_),
    .A1(net773));
 sg13g2_a21o_2 _4057_ (.A2(_1368_),
    .A1(net773),
    .B1(net791),
    .X(_1370_));
 sg13g2_a21oi_1 _4058_ (.A1(net642),
    .A2(net842),
    .Y(_1371_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4059_ (.B1(net876),
    .Y(_1372_),
    .A1(net566),
    .A2(_1369_));
 sg13g2_a21oi_1 _4060_ (.A1(net705),
    .A2(_1371_),
    .Y(_0213_),
    .B1(_1372_));
 sg13g2_a21oi_1 _4061_ (.A1(net611),
    .A2(net853),
    .Y(_1373_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4062_ (.B1(net876),
    .Y(_1374_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .A2(_1369_));
 sg13g2_a21oi_1 _4063_ (.A1(net709),
    .A2(_1373_),
    .Y(_0214_),
    .B1(_1374_));
 sg13g2_a21oi_1 _4064_ (.A1(net630),
    .A2(net842),
    .Y(_1375_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4065_ (.B1(net876),
    .Y(_1376_),
    .A1(net611),
    .A2(_1369_));
 sg13g2_a21oi_1 _4066_ (.A1(net697),
    .A2(_1375_),
    .Y(_0215_),
    .B1(_1376_));
 sg13g2_a21oi_1 _4067_ (.A1(net592),
    .A2(net842),
    .Y(_1377_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4068_ (.B1(net876),
    .Y(_1378_),
    .A1(net630),
    .A2(_1369_));
 sg13g2_a21oi_1 _4069_ (.A1(net695),
    .A2(_1377_),
    .Y(_0216_),
    .B1(_1378_));
 sg13g2_a21oi_1 _4070_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .A2(net842),
    .Y(_1379_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4071_ (.B1(net876),
    .Y(_1380_),
    .A1(net592),
    .A2(_1369_));
 sg13g2_a21oi_1 _4072_ (.A1(net685),
    .A2(_1379_),
    .Y(_0217_),
    .B1(_1380_));
 sg13g2_a21oi_1 _4073_ (.A1(net505),
    .A2(net842),
    .Y(_1381_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4074_ (.B1(net876),
    .Y(_1382_),
    .A1(net636),
    .A2(_1369_));
 sg13g2_a21oi_1 _4075_ (.A1(net683),
    .A2(_1381_),
    .Y(_0218_),
    .B1(_1382_));
 sg13g2_a21oi_1 _4076_ (.A1(net454),
    .A2(net848),
    .Y(_1383_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4077_ (.B1(net876),
    .Y(_1384_),
    .A1(net505),
    .A2(_1369_));
 sg13g2_a21oi_1 _4078_ (.A1(net679),
    .A2(_1383_),
    .Y(_0219_),
    .B1(_1384_));
 sg13g2_a21oi_1 _4079_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ),
    .A2(net848),
    .Y(_1385_),
    .B1(_1370_));
 sg13g2_o21ai_1 _4080_ (.B1(net888),
    .Y(_1386_),
    .A1(net454),
    .A2(_1369_));
 sg13g2_a21oi_1 _4081_ (.A1(net681),
    .A2(_1385_),
    .Y(_0220_),
    .B1(_1386_));
 sg13g2_nor2b_1 _4082_ (.A(_1265_),
    .B_N(_1262_),
    .Y(_1387_));
 sg13g2_nand2b_1 _4083_ (.Y(_1388_),
    .B(_1262_),
    .A_N(_1265_));
 sg13g2_nand2_1 _4084_ (.Y(_1389_),
    .A(_1345_),
    .B(_1387_));
 sg13g2_a21oi_2 _4085_ (.B1(net791),
    .Y(_1390_),
    .A2(_1389_),
    .A1(net773));
 sg13g2_a21o_2 _4086_ (.A2(_1389_),
    .A1(net773),
    .B1(net791),
    .X(_1391_));
 sg13g2_a21oi_1 _4087_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ),
    .A2(net850),
    .Y(_1392_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4088_ (.B1(net892),
    .Y(_1393_),
    .A1(net456),
    .A2(_1390_));
 sg13g2_a21oi_1 _4089_ (.A1(net705),
    .A2(_1392_),
    .Y(_0221_),
    .B1(_1393_));
 sg13g2_a21oi_1 _4090_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ),
    .A2(net847),
    .Y(_1394_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4091_ (.B1(net887),
    .Y(_1395_),
    .A1(net490),
    .A2(_1390_));
 sg13g2_a21oi_1 _4092_ (.A1(net709),
    .A2(_1394_),
    .Y(_0222_),
    .B1(_1395_));
 sg13g2_a21oi_1 _4093_ (.A1(net501),
    .A2(net847),
    .Y(_1396_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4094_ (.B1(net887),
    .Y(_1397_),
    .A1(net539),
    .A2(_1390_));
 sg13g2_a21oi_1 _4095_ (.A1(net697),
    .A2(_1396_),
    .Y(_0223_),
    .B1(_1397_));
 sg13g2_a21oi_1 _4096_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ),
    .A2(net847),
    .Y(_1398_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4097_ (.B1(net887),
    .Y(_1399_),
    .A1(net501),
    .A2(_1390_));
 sg13g2_a21oi_1 _4098_ (.A1(net695),
    .A2(_1398_),
    .Y(_0224_),
    .B1(_1399_));
 sg13g2_a21oi_1 _4099_ (.A1(net533),
    .A2(net850),
    .Y(_1400_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4100_ (.B1(net892),
    .Y(_1401_),
    .A1(net600),
    .A2(_1390_));
 sg13g2_a21oi_1 _4101_ (.A1(net685),
    .A2(_1400_),
    .Y(_0225_),
    .B1(_1401_));
 sg13g2_a21oi_1 _4102_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ),
    .A2(net850),
    .Y(_1402_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4103_ (.B1(net892),
    .Y(_1403_),
    .A1(net533),
    .A2(_1390_));
 sg13g2_a21oi_1 _4104_ (.A1(net684),
    .A2(_1402_),
    .Y(_0226_),
    .B1(_1403_));
 sg13g2_a21oi_1 _4105_ (.A1(net506),
    .A2(net847),
    .Y(_1404_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4106_ (.B1(net887),
    .Y(_1405_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ),
    .A2(_1390_));
 sg13g2_a21oi_1 _4107_ (.A1(net679),
    .A2(_1404_),
    .Y(_0227_),
    .B1(_1405_));
 sg13g2_a21oi_1 _4108_ (.A1(net566),
    .A2(net848),
    .Y(_1406_),
    .B1(_1391_));
 sg13g2_o21ai_1 _4109_ (.B1(net887),
    .Y(_1407_),
    .A1(net506),
    .A2(_1390_));
 sg13g2_a21oi_1 _4110_ (.A1(net682),
    .A2(_1406_),
    .Y(_0228_),
    .B1(_1407_));
 sg13g2_nand3_1 _4111_ (.B(_1265_),
    .C(_1345_),
    .A(_1262_),
    .Y(_1408_));
 sg13g2_a21oi_2 _4112_ (.B1(net792),
    .Y(_1409_),
    .A2(_1408_),
    .A1(net774));
 sg13g2_a21o_2 _4113_ (.A2(_1408_),
    .A1(net775),
    .B1(net792),
    .X(_1410_));
 sg13g2_a21oi_1 _4114_ (.A1(net496),
    .A2(net851),
    .Y(_1411_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4115_ (.B1(net891),
    .Y(_1412_),
    .A1(net535),
    .A2(_1409_));
 sg13g2_a21oi_1 _4116_ (.A1(net705),
    .A2(_1411_),
    .Y(_0229_),
    .B1(_1412_));
 sg13g2_a21oi_1 _4117_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ),
    .A2(net849),
    .Y(_1413_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4118_ (.B1(net891),
    .Y(_1414_),
    .A1(net496),
    .A2(_1409_));
 sg13g2_a21oi_1 _4119_ (.A1(net709),
    .A2(_1413_),
    .Y(_0230_),
    .B1(_1414_));
 sg13g2_a21oi_1 _4120_ (.A1(net621),
    .A2(net850),
    .Y(_1415_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4121_ (.B1(net891),
    .Y(_1416_),
    .A1(net635),
    .A2(_1409_));
 sg13g2_a21oi_1 _4122_ (.A1(net697),
    .A2(_1415_),
    .Y(_0231_),
    .B1(_1416_));
 sg13g2_a21oi_1 _4123_ (.A1(net598),
    .A2(net850),
    .Y(_1417_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4124_ (.B1(net891),
    .Y(_1418_),
    .A1(net621),
    .A2(_1409_));
 sg13g2_a21oi_1 _4125_ (.A1(net695),
    .A2(_1417_),
    .Y(_0232_),
    .B1(_1418_));
 sg13g2_a21oi_1 _4126_ (.A1(net560),
    .A2(net850),
    .Y(_1419_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4127_ (.B1(net893),
    .Y(_1420_),
    .A1(net598),
    .A2(_1409_));
 sg13g2_a21oi_1 _4128_ (.A1(net685),
    .A2(_1419_),
    .Y(_0233_),
    .B1(_1420_));
 sg13g2_a21oi_1 _4129_ (.A1(net527),
    .A2(net850),
    .Y(_1421_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4130_ (.B1(net892),
    .Y(_1422_),
    .A1(net560),
    .A2(_1409_));
 sg13g2_a21oi_1 _4131_ (.A1(net683),
    .A2(_1421_),
    .Y(_0234_),
    .B1(_1422_));
 sg13g2_a21oi_1 _4132_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ),
    .A2(net851),
    .Y(_1423_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4133_ (.B1(net892),
    .Y(_1424_),
    .A1(net527),
    .A2(_1409_));
 sg13g2_a21oi_1 _4134_ (.A1(net679),
    .A2(_1423_),
    .Y(_0235_),
    .B1(_1424_));
 sg13g2_a21oi_1 _4135_ (.A1(net456),
    .A2(net850),
    .Y(_1425_),
    .B1(_1410_));
 sg13g2_o21ai_1 _4136_ (.B1(net891),
    .Y(_1426_),
    .A1(net532),
    .A2(_1409_));
 sg13g2_a21oi_1 _4137_ (.A1(net681),
    .A2(_1425_),
    .Y(_0236_),
    .B1(_1426_));
 sg13g2_nand2b_1 _4138_ (.Y(_1427_),
    .B(_1256_),
    .A_N(_1254_));
 sg13g2_inv_1 _4139_ (.Y(_1428_),
    .A(_1427_));
 sg13g2_nand2_1 _4140_ (.Y(_1429_),
    .A(_1344_),
    .B(_1428_));
 sg13g2_a21oi_2 _4141_ (.B1(net792),
    .Y(_1430_),
    .A2(_1429_),
    .A1(net773));
 sg13g2_a21o_2 _4142_ (.A2(_1429_),
    .A1(net773),
    .B1(net792),
    .X(_1431_));
 sg13g2_a21oi_1 _4143_ (.A1(net555),
    .A2(net849),
    .Y(_1432_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4144_ (.B1(net889),
    .Y(_1433_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ),
    .A2(_1430_));
 sg13g2_a21oi_1 _4145_ (.A1(net705),
    .A2(_1432_),
    .Y(_0237_),
    .B1(_1433_));
 sg13g2_a21oi_1 _4146_ (.A1(net525),
    .A2(net849),
    .Y(_1434_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4147_ (.B1(net890),
    .Y(_1435_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ),
    .A2(_1430_));
 sg13g2_a21oi_1 _4148_ (.A1(net709),
    .A2(_1434_),
    .Y(_0238_),
    .B1(_1435_));
 sg13g2_a21oi_1 _4149_ (.A1(net591),
    .A2(net849),
    .Y(_1436_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4150_ (.B1(net889),
    .Y(_1437_),
    .A1(net525),
    .A2(_1430_));
 sg13g2_a21oi_1 _4151_ (.A1(net697),
    .A2(_1436_),
    .Y(_0239_),
    .B1(_1437_));
 sg13g2_a21oi_1 _4152_ (.A1(net503),
    .A2(net849),
    .Y(_1438_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4153_ (.B1(net889),
    .Y(_1439_),
    .A1(net591),
    .A2(_1430_));
 sg13g2_a21oi_1 _4154_ (.A1(net695),
    .A2(_1438_),
    .Y(_0240_),
    .B1(_1439_));
 sg13g2_a21oi_1 _4155_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ),
    .A2(net849),
    .Y(_1440_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4156_ (.B1(net891),
    .Y(_1441_),
    .A1(net503),
    .A2(_1430_));
 sg13g2_a21oi_1 _4157_ (.A1(net685),
    .A2(_1440_),
    .Y(_0241_),
    .B1(_1441_));
 sg13g2_a21oi_1 _4158_ (.A1(net515),
    .A2(net849),
    .Y(_1442_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4159_ (.B1(net891),
    .Y(_1443_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ),
    .A2(_1430_));
 sg13g2_a21oi_1 _4160_ (.A1(net683),
    .A2(_1442_),
    .Y(_0242_),
    .B1(_1443_));
 sg13g2_a21oi_1 _4161_ (.A1(net469),
    .A2(net851),
    .Y(_1444_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4162_ (.B1(net890),
    .Y(_1445_),
    .A1(net515),
    .A2(_1430_));
 sg13g2_a21oi_1 _4163_ (.A1(net679),
    .A2(_1444_),
    .Y(_0243_),
    .B1(_1445_));
 sg13g2_a21oi_1 _4164_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ),
    .A2(net849),
    .Y(_1446_),
    .B1(_1431_));
 sg13g2_o21ai_1 _4165_ (.B1(net891),
    .Y(_1447_),
    .A1(net469),
    .A2(_1430_));
 sg13g2_a21oi_1 _4166_ (.A1(net681),
    .A2(_1446_),
    .Y(_0244_),
    .B1(_1447_));
 sg13g2_nand2_2 _4167_ (.Y(_1448_),
    .A(_1366_),
    .B(_1428_));
 sg13g2_a21oi_2 _4168_ (.B1(net792),
    .Y(_1449_),
    .A2(_1448_),
    .A1(net774));
 sg13g2_a21o_2 _4169_ (.A2(_1448_),
    .A1(net774),
    .B1(net792),
    .X(_1450_));
 sg13g2_a21oi_1 _4170_ (.A1(net529),
    .A2(net844),
    .Y(_1451_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4171_ (.B1(net889),
    .Y(_1452_),
    .A1(net510),
    .A2(_1449_));
 sg13g2_a21oi_1 _4172_ (.A1(net705),
    .A2(_1451_),
    .Y(_0245_),
    .B1(_1452_));
 sg13g2_a21oi_1 _4173_ (.A1(net480),
    .A2(net843),
    .Y(_1453_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4174_ (.B1(net889),
    .Y(_1454_),
    .A1(net529),
    .A2(_1449_));
 sg13g2_a21oi_1 _4175_ (.A1(net709),
    .A2(_1453_),
    .Y(_0246_),
    .B1(_1454_));
 sg13g2_a21oi_1 _4176_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ),
    .A2(net843),
    .Y(_1455_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4177_ (.B1(net884),
    .Y(_1456_),
    .A1(net480),
    .A2(_1449_));
 sg13g2_a21oi_1 _4178_ (.A1(net697),
    .A2(_1455_),
    .Y(_0247_),
    .B1(_1456_));
 sg13g2_a21oi_1 _4179_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ),
    .A2(net843),
    .Y(_1457_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4180_ (.B1(net883),
    .Y(_1458_),
    .A1(net545),
    .A2(_1449_));
 sg13g2_a21oi_1 _4181_ (.A1(net695),
    .A2(_1457_),
    .Y(_0248_),
    .B1(_1458_));
 sg13g2_a21oi_1 _4182_ (.A1(net482),
    .A2(net843),
    .Y(_1459_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4183_ (.B1(net883),
    .Y(_1460_),
    .A1(net604),
    .A2(_1449_));
 sg13g2_a21oi_1 _4184_ (.A1(net685),
    .A2(_1459_),
    .Y(_0249_),
    .B1(_1460_));
 sg13g2_a21oi_1 _4185_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ),
    .A2(net843),
    .Y(_1461_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4186_ (.B1(net884),
    .Y(_1462_),
    .A1(net482),
    .A2(_1449_));
 sg13g2_a21oi_1 _4187_ (.A1(net683),
    .A2(_1461_),
    .Y(_0250_),
    .B1(_1462_));
 sg13g2_a21oi_1 _4188_ (.A1(net475),
    .A2(net843),
    .Y(_1463_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4189_ (.B1(net885),
    .Y(_1464_),
    .A1(net538),
    .A2(_1449_));
 sg13g2_a21oi_1 _4190_ (.A1(net679),
    .A2(_1463_),
    .Y(_0251_),
    .B1(_1464_));
 sg13g2_a21oi_1 _4191_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ),
    .A2(net844),
    .Y(_1465_),
    .B1(_1450_));
 sg13g2_o21ai_1 _4192_ (.B1(net884),
    .Y(_1466_),
    .A1(net475),
    .A2(_1449_));
 sg13g2_a21oi_1 _4193_ (.A1(net681),
    .A2(_1465_),
    .Y(_0252_),
    .B1(_1466_));
 sg13g2_nand2_2 _4194_ (.Y(_1467_),
    .A(_1387_),
    .B(_1428_));
 sg13g2_a21oi_2 _4195_ (.B1(net792),
    .Y(_1468_),
    .A2(_1467_),
    .A1(net774));
 sg13g2_a21o_2 _4196_ (.A2(_1467_),
    .A1(net774),
    .B1(net792),
    .X(_1469_));
 sg13g2_a21oi_1 _4197_ (.A1(net537),
    .A2(net844),
    .Y(_1470_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4198_ (.B1(net889),
    .Y(_1471_),
    .A1(net487),
    .A2(_1468_));
 sg13g2_a21oi_1 _4199_ (.A1(net705),
    .A2(_1470_),
    .Y(_0253_),
    .B1(_1471_));
 sg13g2_a21oi_1 _4200_ (.A1(net541),
    .A2(net844),
    .Y(_1472_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4201_ (.B1(net889),
    .Y(_1473_),
    .A1(net537),
    .A2(_1468_));
 sg13g2_a21oi_1 _4202_ (.A1(net709),
    .A2(_1472_),
    .Y(_0254_),
    .B1(_1473_));
 sg13g2_a21oi_1 _4203_ (.A1(net562),
    .A2(net844),
    .Y(_1474_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4204_ (.B1(net889),
    .Y(_1475_),
    .A1(net541),
    .A2(_1468_));
 sg13g2_a21oi_1 _4205_ (.A1(net697),
    .A2(_1474_),
    .Y(_0255_),
    .B1(_1475_));
 sg13g2_a21oi_1 _4206_ (.A1(net542),
    .A2(net843),
    .Y(_1476_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4207_ (.B1(net884),
    .Y(_1477_),
    .A1(net562),
    .A2(_1468_));
 sg13g2_a21oi_1 _4208_ (.A1(net695),
    .A2(_1476_),
    .Y(_0256_),
    .B1(_1477_));
 sg13g2_a21oi_1 _4209_ (.A1(net478),
    .A2(net843),
    .Y(_1478_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4210_ (.B1(net884),
    .Y(_1479_),
    .A1(net542),
    .A2(_1468_));
 sg13g2_a21oi_1 _4211_ (.A1(net685),
    .A2(_1478_),
    .Y(_0257_),
    .B1(_1479_));
 sg13g2_a21oi_1 _4212_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ),
    .A2(net844),
    .Y(_1480_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4213_ (.B1(net884),
    .Y(_1481_),
    .A1(net478),
    .A2(_1468_));
 sg13g2_a21oi_1 _4214_ (.A1(net683),
    .A2(_1480_),
    .Y(_0258_),
    .B1(_1481_));
 sg13g2_a21oi_1 _4215_ (.A1(net508),
    .A2(net852),
    .Y(_1482_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4216_ (.B1(net884),
    .Y(_1483_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ),
    .A2(_1468_));
 sg13g2_a21oi_1 _4217_ (.A1(net679),
    .A2(_1482_),
    .Y(_0259_),
    .B1(_1483_));
 sg13g2_a21oi_1 _4218_ (.A1(net510),
    .A2(net844),
    .Y(_1484_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4219_ (.B1(net884),
    .Y(_1485_),
    .A1(net508),
    .A2(_1468_));
 sg13g2_a21oi_1 _4220_ (.A1(net681),
    .A2(_1484_),
    .Y(_0260_),
    .B1(_1485_));
 sg13g2_nand3_1 _4221_ (.B(_1265_),
    .C(_1428_),
    .A(_1262_),
    .Y(_1486_));
 sg13g2_a21oi_2 _4222_ (.B1(net791),
    .Y(_1487_),
    .A2(_1486_),
    .A1(net773));
 sg13g2_a21o_2 _4223_ (.A2(_1486_),
    .A1(net773),
    .B1(net791),
    .X(_1488_));
 sg13g2_a21oi_1 _4224_ (.A1(net493),
    .A2(net845),
    .Y(_1489_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4225_ (.B1(net888),
    .Y(_1490_),
    .A1(net540),
    .A2(_1487_));
 sg13g2_a21oi_1 _4226_ (.A1(net705),
    .A2(_1489_),
    .Y(_0261_),
    .B1(_1490_));
 sg13g2_a21oi_1 _4227_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ),
    .A2(net845),
    .Y(_1491_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4228_ (.B1(net888),
    .Y(_1492_),
    .A1(net493),
    .A2(_1487_));
 sg13g2_a21oi_1 _4229_ (.A1(net709),
    .A2(_1491_),
    .Y(_0262_),
    .B1(_1492_));
 sg13g2_a21oi_1 _4230_ (.A1(net370),
    .A2(net845),
    .Y(_1493_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4231_ (.B1(net888),
    .Y(_1494_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ),
    .A2(_1487_));
 sg13g2_a21oi_1 _4232_ (.A1(net697),
    .A2(_1493_),
    .Y(_0263_),
    .B1(_1494_));
 sg13g2_a21oi_1 _4233_ (.A1(net536),
    .A2(net845),
    .Y(_1495_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4234_ (.B1(net888),
    .Y(_1496_),
    .A1(net370),
    .A2(_1487_));
 sg13g2_a21oi_1 _4235_ (.A1(net695),
    .A2(_1495_),
    .Y(_0264_),
    .B1(_1496_));
 sg13g2_a21oi_1 _4236_ (.A1(net512),
    .A2(net845),
    .Y(_1497_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4237_ (.B1(net888),
    .Y(_1498_),
    .A1(net536),
    .A2(_1487_));
 sg13g2_a21oi_1 _4238_ (.A1(net685),
    .A2(_1497_),
    .Y(_0265_),
    .B1(_1498_));
 sg13g2_a21oi_1 _4239_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ),
    .A2(net845),
    .Y(_1499_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4240_ (.B1(net888),
    .Y(_1500_),
    .A1(net512),
    .A2(_1487_));
 sg13g2_a21oi_1 _4241_ (.A1(net683),
    .A2(_1499_),
    .Y(_0266_),
    .B1(_1500_));
 sg13g2_a21oi_1 _4242_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ),
    .A2(net845),
    .Y(_1501_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4243_ (.B1(net881),
    .Y(_1502_),
    .A1(net523),
    .A2(_1487_));
 sg13g2_a21oi_1 _4244_ (.A1(net679),
    .A2(_1501_),
    .Y(_0267_),
    .B1(_1502_));
 sg13g2_a21oi_1 _4245_ (.A1(net487),
    .A2(net845),
    .Y(_1503_),
    .B1(_1488_));
 sg13g2_o21ai_1 _4246_ (.B1(net881),
    .Y(_1504_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ),
    .A2(_1487_));
 sg13g2_a21oi_1 _4247_ (.A1(net681),
    .A2(_1503_),
    .Y(_0268_),
    .B1(_1504_));
 sg13g2_nand2b_2 _4248_ (.Y(_1505_),
    .B(_1254_),
    .A_N(_1256_));
 sg13g2_nand2b_1 _4249_ (.Y(_1506_),
    .B(_1344_),
    .A_N(_1258_));
 sg13g2_nor2_1 _4250_ (.A(_1505_),
    .B(_1506_),
    .Y(_1507_));
 sg13g2_o21ai_1 _4251_ (.B1(net873),
    .Y(_1508_),
    .A1(net440),
    .A2(net721));
 sg13g2_a21oi_1 _4252_ (.A1(net717),
    .A2(net721),
    .Y(_0269_),
    .B1(_1508_));
 sg13g2_o21ai_1 _4253_ (.B1(net879),
    .Y(_1509_),
    .A1(net383),
    .A2(net721));
 sg13g2_a21oi_1 _4254_ (.A1(net715),
    .A2(net722),
    .Y(_0270_),
    .B1(_1509_));
 sg13g2_o21ai_1 _4255_ (.B1(net877),
    .Y(_1510_),
    .A1(net448),
    .A2(net721));
 sg13g2_a21oi_1 _4256_ (.A1(net711),
    .A2(net721),
    .Y(_0271_),
    .B1(_1510_));
 sg13g2_o21ai_1 _4257_ (.B1(net883),
    .Y(_1511_),
    .A1(net390),
    .A2(net722));
 sg13g2_a21oi_1 _4258_ (.A1(net701),
    .A2(net722),
    .Y(_0272_),
    .B1(_1511_));
 sg13g2_o21ai_1 _4259_ (.B1(net879),
    .Y(_1512_),
    .A1(net439),
    .A2(net722));
 sg13g2_a21oi_1 _4260_ (.A1(net703),
    .A2(net722),
    .Y(_0273_),
    .B1(_1512_));
 sg13g2_o21ai_1 _4261_ (.B1(net885),
    .Y(_1513_),
    .A1(net419),
    .A2(net722));
 sg13g2_a21oi_1 _4262_ (.A1(net688),
    .A2(net721),
    .Y(_0274_),
    .B1(_1513_));
 sg13g2_o21ai_1 _4263_ (.B1(net894),
    .Y(_1514_),
    .A1(net380),
    .A2(net723));
 sg13g2_a21oi_1 _4264_ (.A1(net689),
    .A2(net723),
    .Y(_0275_),
    .B1(_1514_));
 sg13g2_o21ai_1 _4265_ (.B1(net873),
    .Y(_1515_),
    .A1(net426),
    .A2(net721));
 sg13g2_a21oi_1 _4266_ (.A1(net691),
    .A2(net721),
    .Y(_0276_),
    .B1(_1515_));
 sg13g2_nor3_1 _4267_ (.A(_1258_),
    .B(_1367_),
    .C(_1505_),
    .Y(_1516_));
 sg13g2_o21ai_1 _4268_ (.B1(net878),
    .Y(_1517_),
    .A1(net376),
    .A2(net737));
 sg13g2_a21oi_1 _4269_ (.A1(net717),
    .A2(net737),
    .Y(_0277_),
    .B1(_1517_));
 sg13g2_o21ai_1 _4270_ (.B1(net881),
    .Y(_1518_),
    .A1(net514),
    .A2(_1516_));
 sg13g2_a21oi_1 _4271_ (.A1(net715),
    .A2(net738),
    .Y(_0278_),
    .B1(_1518_));
 sg13g2_o21ai_1 _4272_ (.B1(net877),
    .Y(_1519_),
    .A1(net471),
    .A2(net737));
 sg13g2_a21oi_1 _4273_ (.A1(net711),
    .A2(net737),
    .Y(_0279_),
    .B1(_1519_));
 sg13g2_o21ai_1 _4274_ (.B1(net878),
    .Y(_1520_),
    .A1(net365),
    .A2(net738));
 sg13g2_a21oi_1 _4275_ (.A1(net700),
    .A2(net738),
    .Y(_0280_),
    .B1(_1520_));
 sg13g2_o21ai_1 _4276_ (.B1(net877),
    .Y(_1521_),
    .A1(net367),
    .A2(net737));
 sg13g2_a21oi_1 _4277_ (.A1(net702),
    .A2(net737),
    .Y(_0281_),
    .B1(_1521_));
 sg13g2_o21ai_1 _4278_ (.B1(net881),
    .Y(_1522_),
    .A1(net405),
    .A2(net738));
 sg13g2_a21oi_1 _4279_ (.A1(net688),
    .A2(net738),
    .Y(_0282_),
    .B1(_1522_));
 sg13g2_o21ai_1 _4280_ (.B1(net881),
    .Y(_1523_),
    .A1(net438),
    .A2(net738));
 sg13g2_a21oi_1 _4281_ (.A1(net690),
    .A2(net738),
    .Y(_0283_),
    .B1(_1523_));
 sg13g2_o21ai_1 _4282_ (.B1(net877),
    .Y(_1524_),
    .A1(net495),
    .A2(net737));
 sg13g2_a21oi_1 _4283_ (.A1(net692),
    .A2(net737),
    .Y(_0284_),
    .B1(_1524_));
 sg13g2_nor3_1 _4284_ (.A(_1258_),
    .B(_1388_),
    .C(_1505_),
    .Y(_1525_));
 sg13g2_o21ai_1 _4285_ (.B1(net885),
    .Y(_1526_),
    .A1(net395),
    .A2(net736));
 sg13g2_a21oi_1 _4286_ (.A1(net718),
    .A2(net736),
    .Y(_0285_),
    .B1(_1526_));
 sg13g2_o21ai_1 _4287_ (.B1(net877),
    .Y(_1527_),
    .A1(net434),
    .A2(net734));
 sg13g2_a21oi_1 _4288_ (.A1(net715),
    .A2(net734),
    .Y(_0286_),
    .B1(_1527_));
 sg13g2_o21ai_1 _4289_ (.B1(net879),
    .Y(_1528_),
    .A1(net378),
    .A2(net734));
 sg13g2_a21oi_1 _4290_ (.A1(net711),
    .A2(net734),
    .Y(_0287_),
    .B1(_1528_));
 sg13g2_o21ai_1 _4291_ (.B1(net882),
    .Y(_1529_),
    .A1(net431),
    .A2(net735));
 sg13g2_a21oi_1 _4292_ (.A1(net701),
    .A2(net735),
    .Y(_0288_),
    .B1(_1529_));
 sg13g2_o21ai_1 _4293_ (.B1(net885),
    .Y(_1530_),
    .A1(net393),
    .A2(net735));
 sg13g2_a21oi_1 _4294_ (.A1(net703),
    .A2(net735),
    .Y(_0289_),
    .B1(_1530_));
 sg13g2_o21ai_1 _4295_ (.B1(net880),
    .Y(_1531_),
    .A1(net428),
    .A2(net734));
 sg13g2_a21oi_1 _4296_ (.A1(net687),
    .A2(net734),
    .Y(_0290_),
    .B1(_1531_));
 sg13g2_o21ai_1 _4297_ (.B1(net890),
    .Y(_1532_),
    .A1(net417),
    .A2(net736));
 sg13g2_a21oi_1 _4298_ (.A1(net689),
    .A2(net736),
    .Y(_0291_),
    .B1(_1532_));
 sg13g2_o21ai_1 _4299_ (.B1(net877),
    .Y(_1533_),
    .A1(net477),
    .A2(net734));
 sg13g2_a21oi_1 _4300_ (.A1(net692),
    .A2(net734),
    .Y(_0292_),
    .B1(_1533_));
 sg13g2_nor3_2 _4301_ (.A(_1258_),
    .B(_1266_),
    .C(_1505_),
    .Y(_1534_));
 sg13g2_o21ai_1 _4302_ (.B1(net881),
    .Y(_1535_),
    .A1(net452),
    .A2(net733));
 sg13g2_a21oi_1 _4303_ (.A1(net717),
    .A2(net733),
    .Y(_0293_),
    .B1(_1535_));
 sg13g2_o21ai_1 _4304_ (.B1(net886),
    .Y(_1536_),
    .A1(net472),
    .A2(net733));
 sg13g2_a21oi_1 _4305_ (.A1(net714),
    .A2(net733),
    .Y(_0294_),
    .B1(_1536_));
 sg13g2_o21ai_1 _4306_ (.B1(net877),
    .Y(_1537_),
    .A1(net492),
    .A2(net732));
 sg13g2_a21oi_1 _4307_ (.A1(net711),
    .A2(net732),
    .Y(_0295_),
    .B1(_1537_));
 sg13g2_o21ai_1 _4308_ (.B1(net878),
    .Y(_1538_),
    .A1(net394),
    .A2(net732));
 sg13g2_a21oi_1 _4309_ (.A1(net700),
    .A2(net732),
    .Y(_0296_),
    .B1(_1538_));
 sg13g2_o21ai_1 _4310_ (.B1(net879),
    .Y(_1539_),
    .A1(net451),
    .A2(net732));
 sg13g2_a21oi_1 _4311_ (.A1(net703),
    .A2(net733),
    .Y(_0297_),
    .B1(_1539_));
 sg13g2_o21ai_1 _4312_ (.B1(net879),
    .Y(_1540_),
    .A1(net406),
    .A2(net733));
 sg13g2_a21oi_1 _4313_ (.A1(net687),
    .A2(net732),
    .Y(_0298_),
    .B1(_1540_));
 sg13g2_o21ai_1 _4314_ (.B1(net885),
    .Y(_1541_),
    .A1(net449),
    .A2(_1534_));
 sg13g2_a21oi_1 _4315_ (.A1(net689),
    .A2(net733),
    .Y(_0299_),
    .B1(_1541_));
 sg13g2_o21ai_1 _4316_ (.B1(net877),
    .Y(_1542_),
    .A1(net464),
    .A2(net732));
 sg13g2_a21oi_1 _4317_ (.A1(net691),
    .A2(net732),
    .Y(_0300_),
    .B1(_1542_));
 sg13g2_nor2_2 _4318_ (.A(_1257_),
    .B(_1506_),
    .Y(_1543_));
 sg13g2_o21ai_1 _4319_ (.B1(net873),
    .Y(_1544_),
    .A1(net460),
    .A2(net719));
 sg13g2_a21oi_1 _4320_ (.A1(net717),
    .A2(net719),
    .Y(_0301_),
    .B1(_1544_));
 sg13g2_o21ai_1 _4321_ (.B1(net878),
    .Y(_1545_),
    .A1(net459),
    .A2(net720));
 sg13g2_a21oi_1 _4322_ (.A1(net714),
    .A2(net720),
    .Y(_0302_),
    .B1(_1545_));
 sg13g2_o21ai_1 _4323_ (.B1(net888),
    .Y(_1546_),
    .A1(net561),
    .A2(net719));
 sg13g2_a21oi_1 _4324_ (.A1(net712),
    .A2(net719),
    .Y(_0303_),
    .B1(_1546_));
 sg13g2_o21ai_1 _4325_ (.B1(net873),
    .Y(_1547_),
    .A1(net427),
    .A2(net719));
 sg13g2_a21oi_1 _4326_ (.A1(net700),
    .A2(net720),
    .Y(_0304_),
    .B1(_1547_));
 sg13g2_o21ai_1 _4327_ (.B1(net873),
    .Y(_1548_),
    .A1(net404),
    .A2(net720));
 sg13g2_a21oi_1 _4328_ (.A1(net702),
    .A2(net720),
    .Y(_0305_),
    .B1(_1548_));
 sg13g2_o21ai_1 _4329_ (.B1(net873),
    .Y(_1549_),
    .A1(net445),
    .A2(net719));
 sg13g2_a21oi_1 _4330_ (.A1(net687),
    .A2(net719),
    .Y(_0306_),
    .B1(_1549_));
 sg13g2_o21ai_1 _4331_ (.B1(net881),
    .Y(_1550_),
    .A1(net409),
    .A2(net719));
 sg13g2_a21oi_1 _4332_ (.A1(net690),
    .A2(_1543_),
    .Y(_0307_),
    .B1(_1550_));
 sg13g2_o21ai_1 _4333_ (.B1(net873),
    .Y(_1551_),
    .A1(net410),
    .A2(net720));
 sg13g2_a21oi_1 _4334_ (.A1(net691),
    .A2(net720),
    .Y(_0308_),
    .B1(_1551_));
 sg13g2_nor3_1 _4335_ (.A(_1257_),
    .B(_1258_),
    .C(_1367_),
    .Y(_1552_));
 sg13g2_o21ai_1 _4336_ (.B1(net883),
    .Y(_1553_),
    .A1(net411),
    .A2(net729));
 sg13g2_a21oi_1 _4337_ (.A1(net717),
    .A2(net729),
    .Y(_0309_),
    .B1(_1553_));
 sg13g2_o21ai_1 _4338_ (.B1(net890),
    .Y(_1554_),
    .A1(net486),
    .A2(net731));
 sg13g2_a21oi_1 _4339_ (.A1(net714),
    .A2(net731),
    .Y(_0310_),
    .B1(_1554_));
 sg13g2_o21ai_1 _4340_ (.B1(net882),
    .Y(_1555_),
    .A1(net391),
    .A2(net730));
 sg13g2_a21oi_1 _4341_ (.A1(net711),
    .A2(net730),
    .Y(_0311_),
    .B1(_1555_));
 sg13g2_o21ai_1 _4342_ (.B1(net882),
    .Y(_1556_),
    .A1(net433),
    .A2(net730));
 sg13g2_a21oi_1 _4343_ (.A1(net700),
    .A2(net730),
    .Y(_0312_),
    .B1(_1556_));
 sg13g2_o21ai_1 _4344_ (.B1(net883),
    .Y(_1557_),
    .A1(net379),
    .A2(net729));
 sg13g2_a21oi_1 _4345_ (.A1(net702),
    .A2(net729),
    .Y(_0313_),
    .B1(_1557_));
 sg13g2_o21ai_1 _4346_ (.B1(net882),
    .Y(_1558_),
    .A1(net377),
    .A2(net729));
 sg13g2_a21oi_1 _4347_ (.A1(net687),
    .A2(net729),
    .Y(_0314_),
    .B1(_1558_));
 sg13g2_o21ai_1 _4348_ (.B1(net885),
    .Y(_1559_),
    .A1(net474),
    .A2(net731));
 sg13g2_a21oi_1 _4349_ (.A1(net689),
    .A2(net731),
    .Y(_0315_),
    .B1(_1559_));
 sg13g2_o21ai_1 _4350_ (.B1(net883),
    .Y(_1560_),
    .A1(net382),
    .A2(net729));
 sg13g2_a21oi_1 _4351_ (.A1(net691),
    .A2(net729),
    .Y(_0316_),
    .B1(_1560_));
 sg13g2_nor3_2 _4352_ (.A(_1257_),
    .B(_1258_),
    .C(_1388_),
    .Y(_1561_));
 sg13g2_o21ai_1 _4353_ (.B1(net892),
    .Y(_1562_),
    .A1(net550),
    .A2(net728));
 sg13g2_a21oi_1 _4354_ (.A1(_1793_),
    .A2(net728),
    .Y(_0317_),
    .B1(_1562_));
 sg13g2_o21ai_1 _4355_ (.B1(net893),
    .Y(_1563_),
    .A1(net381),
    .A2(net728));
 sg13g2_a21oi_1 _4356_ (.A1(net716),
    .A2(net728),
    .Y(_0318_),
    .B1(_1563_));
 sg13g2_o21ai_1 _4357_ (.B1(net882),
    .Y(_1564_),
    .A1(net412),
    .A2(net727));
 sg13g2_a21oi_1 _4358_ (.A1(net711),
    .A2(net727),
    .Y(_0319_),
    .B1(_1564_));
 sg13g2_o21ai_1 _4359_ (.B1(net893),
    .Y(_1565_),
    .A1(net468),
    .A2(net728));
 sg13g2_a21oi_1 _4360_ (.A1(_0542_),
    .A2(net728),
    .Y(_0320_),
    .B1(_1565_));
 sg13g2_o21ai_1 _4361_ (.B1(net879),
    .Y(_1566_),
    .A1(net369),
    .A2(net727));
 sg13g2_a21oi_1 _4362_ (.A1(net702),
    .A2(net727),
    .Y(_0321_),
    .B1(_1566_));
 sg13g2_o21ai_1 _4363_ (.B1(net882),
    .Y(_1567_),
    .A1(net485),
    .A2(net727));
 sg13g2_a21oi_1 _4364_ (.A1(net687),
    .A2(net727),
    .Y(_0322_),
    .B1(_1567_));
 sg13g2_o21ai_1 _4365_ (.B1(net892),
    .Y(_1568_),
    .A1(net465),
    .A2(net728));
 sg13g2_a21oi_1 _4366_ (.A1(_0410_),
    .A2(net728),
    .Y(_0323_),
    .B1(_1568_));
 sg13g2_o21ai_1 _4367_ (.B1(net879),
    .Y(_1569_),
    .A1(net453),
    .A2(net727));
 sg13g2_a21oi_1 _4368_ (.A1(net692),
    .A2(net727),
    .Y(_0324_),
    .B1(_1569_));
 sg13g2_dfrbp_1 _4369_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net79),
    .D(_0027_),
    .Q_N(_2180_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[16] ));
 sg13g2_dfrbp_1 _4370_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net65),
    .D(_0028_),
    .Q_N(_2179_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[17] ));
 sg13g2_dfrbp_1 _4371_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net63),
    .D(_0029_),
    .Q_N(_2178_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[18] ));
 sg13g2_dfrbp_1 _4372_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net61),
    .D(_0030_),
    .Q_N(_2177_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[19] ));
 sg13g2_dfrbp_1 _4373_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net59),
    .D(_0031_),
    .Q_N(_2176_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ));
 sg13g2_dfrbp_1 _4374_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net57),
    .D(_0032_),
    .Q_N(_2175_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ));
 sg13g2_dfrbp_1 _4375_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net55),
    .D(_0033_),
    .Q_N(_2174_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ));
 sg13g2_dfrbp_1 _4376_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net53),
    .D(_0034_),
    .Q_N(_0017_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ));
 sg13g2_dfrbp_1 _4377_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net52),
    .D(net322),
    .Q_N(_2173_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.stop_txn_reg ));
 sg13g2_dfrbp_1 _4378_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net51),
    .D(_0036_),
    .Q_N(_2172_),
    .Q(\cpu_instance.ctrl_instance.state[0] ));
 sg13g2_dfrbp_1 _4379_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net49),
    .D(net661),
    .Q_N(_2171_),
    .Q(\cpu_instance.ctrl_instance.state[1] ));
 sg13g2_dfrbp_1 _4380_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net47),
    .D(net656),
    .Q_N(_2170_),
    .Q(\cpu_instance.ctrl_instance.state[2] ));
 sg13g2_dfrbp_1 _4381_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net45),
    .D(_0039_),
    .Q_N(_2169_),
    .Q(\cpu_instance.ctrl_instance.state[3] ));
 sg13g2_dfrbp_1 _4382_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net43),
    .D(_0040_),
    .Q_N(_2168_),
    .Q(\cpu_instance.mux_instance.sel[0] ));
 sg13g2_dfrbp_1 _4383_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net42),
    .D(_0041_),
    .Q_N(_2167_),
    .Q(\cpu_instance.mux_instance.sel[1] ));
 sg13g2_dfrbp_1 _4384_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net41),
    .D(_0042_),
    .Q_N(_2166_),
    .Q(\cpu_instance.ctrl_instance.use_register_bank_in ));
 sg13g2_dfrbp_1 _4385_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net39),
    .D(_0043_),
    .Q_N(_2165_),
    .Q(\cpu_instance.ctrl_instance.use_register_bank_out_1 ));
 sg13g2_dfrbp_1 _4386_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net37),
    .D(_0044_),
    .Q_N(_2164_),
    .Q(\cpu_instance.alu_instance.op[0] ));
 sg13g2_dfrbp_1 _4387_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net35),
    .D(_0045_),
    .Q_N(_2163_),
    .Q(\cpu_instance.alu_instance.op[1] ));
 sg13g2_dfrbp_1 _4388_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net33),
    .D(_0046_),
    .Q_N(_2162_),
    .Q(\cpu_instance.alu_instance.op[2] ));
 sg13g2_dfrbp_1 _4389_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net31),
    .D(_0047_),
    .Q_N(_2161_),
    .Q(\cpu_instance.alu_instance.op[3] ));
 sg13g2_dfrbp_1 _4390_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net29),
    .D(_0048_),
    .Q_N(_2160_),
    .Q(\cpu_instance.ctrl_instance.flag_carry ));
 sg13g2_dfrbp_1 _4391_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net27),
    .D(_0049_),
    .Q_N(_2159_),
    .Q(\cpu_instance.ctrl_instance.flag_zero ));
 sg13g2_dfrbp_1 _4392_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net25),
    .D(_0050_),
    .Q_N(_0022_),
    .Q(\cpu_instance.reg_op ));
 sg13g2_dfrbp_1 _4393_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net24),
    .D(_0051_),
    .Q_N(_2158_),
    .Q(\cpu_instance.mem_ctrl_op[0] ));
 sg13g2_dfrbp_1 _4394_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net23),
    .D(_0052_),
    .Q_N(_2157_),
    .Q(\cpu_instance.mem_ctrl_op[1] ));
 sg13g2_dfrbp_1 _4395_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net22),
    .D(_0053_),
    .Q_N(_2156_),
    .Q(\cpu_instance.addr_reg_op[0] ));
 sg13g2_dfrbp_1 _4396_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net21),
    .D(_0054_),
    .Q_N(_2155_),
    .Q(\cpu_instance.addr_reg_op[1] ));
 sg13g2_dfrbp_1 _4397_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net20),
    .D(_0055_),
    .Q_N(_0026_),
    .Q(\cpu_instance.addr_reg_op[2] ));
 sg13g2_dfrbp_1 _4398_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net19),
    .D(_0056_),
    .Q_N(_2154_),
    .Q(\cpu_instance.reg_in_sel[0] ));
 sg13g2_dfrbp_1 _4399_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net17),
    .D(_0057_),
    .Q_N(_2153_),
    .Q(\cpu_instance.reg_in_sel[1] ));
 sg13g2_dfrbp_1 _4400_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net15),
    .D(_0058_),
    .Q_N(_2152_),
    .Q(\cpu_instance.reg_1_out_sel[0] ));
 sg13g2_dfrbp_1 _4401_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net13),
    .D(_0059_),
    .Q_N(_2151_),
    .Q(\cpu_instance.reg_1_out_sel[1] ));
 sg13g2_dfrbp_1 _4402_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net309),
    .D(_0060_),
    .Q_N(\cpu_instance.mem_instance.addr[24] ),
    .Q(\cpu_instance.addr_sel ));
 sg13g2_dfrbp_1 _4403_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net308),
    .D(net408),
    .Q_N(_2150_),
    .Q(\cpu_instance.ctrl_instance.jmp_op_addr_sel ));
 sg13g2_dfrbp_1 _4404_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net306),
    .D(_0062_),
    .Q_N(_2149_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][1] ));
 sg13g2_dfrbp_1 _4405_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net304),
    .D(_0063_),
    .Q_N(_2148_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ));
 sg13g2_dfrbp_1 _4406_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net302),
    .D(_0064_),
    .Q_N(_2147_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ));
 sg13g2_dfrbp_1 _4407_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net300),
    .D(_0065_),
    .Q_N(_2146_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ));
 sg13g2_dfrbp_1 _4408_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net298),
    .D(_0066_),
    .Q_N(_2145_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ));
 sg13g2_dfrbp_1 _4409_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net296),
    .D(_0067_),
    .Q_N(_2144_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ));
 sg13g2_dfrbp_1 _4410_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net294),
    .D(_0068_),
    .Q_N(_2143_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][7] ));
 sg13g2_dfrbp_1 _4411_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net292),
    .D(_0069_),
    .Q_N(_2142_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][8] ));
 sg13g2_dfrbp_1 _4412_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net290),
    .D(_0070_),
    .Q_N(_2141_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ));
 sg13g2_dfrbp_1 _4413_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net288),
    .D(_0071_),
    .Q_N(_2140_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ));
 sg13g2_dfrbp_1 _4414_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net286),
    .D(_0072_),
    .Q_N(_2139_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ));
 sg13g2_dfrbp_1 _4415_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net284),
    .D(_0073_),
    .Q_N(_2138_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ));
 sg13g2_dfrbp_1 _4416_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net282),
    .D(_0074_),
    .Q_N(_2137_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ));
 sg13g2_dfrbp_1 _4417_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net280),
    .D(_0075_),
    .Q_N(_2136_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ));
 sg13g2_dfrbp_1 _4418_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net278),
    .D(_0076_),
    .Q_N(_2135_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ));
 sg13g2_dfrbp_1 _4419_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net276),
    .D(_0077_),
    .Q_N(_2134_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ));
 sg13g2_dfrbp_1 _4420_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net275),
    .D(net389),
    .Q_N(_2133_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ));
 sg13g2_dfrbp_1 _4421_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net274),
    .D(_0079_),
    .Q_N(_2132_),
    .Q(\cpu_instance.mem_instance.data_ready ));
 sg13g2_dfrbp_1 _4422_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net273),
    .D(net554),
    .Q_N(_2131_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 _4423_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net271),
    .D(net430),
    .Q_N(_2130_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 _4424_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net269),
    .D(net386),
    .Q_N(_2129_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 _4425_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net267),
    .D(net623),
    .Q_N(_2128_),
    .Q(\cpu_instance.mem_instance.data_req ));
 sg13g2_dfrbp_1 _4426_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net266),
    .D(_0084_),
    .Q_N(_2127_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[0] ));
 sg13g2_dfrbp_1 _4427_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net265),
    .D(_0085_),
    .Q_N(_2126_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[1] ));
 sg13g2_dfrbp_1 _4428_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net264),
    .D(_0086_),
    .Q_N(_2125_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[2] ));
 sg13g2_dfrbp_1 _4429_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net263),
    .D(_0087_),
    .Q_N(_2124_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[3] ));
 sg13g2_dfrbp_1 _4430_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net262),
    .D(_0088_),
    .Q_N(_0016_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ));
 sg13g2_dfrbp_1 _4431_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net260),
    .D(net673),
    .Q_N(_2123_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ));
 sg13g2_dfrbp_1 _4432_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net258),
    .D(_0090_),
    .Q_N(_0023_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ));
 sg13g2_dfrbp_1 _4433_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net256),
    .D(_0091_),
    .Q_N(_0025_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.is_writing ));
 sg13g2_dfrbp_1 _4434_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net254),
    .D(_0092_),
    .Q_N(_2122_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ));
 sg13g2_dfrbp_1 _4435_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net252),
    .D(net628),
    .Q_N(_2121_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ));
 sg13g2_dfrbp_1 _4436_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net250),
    .D(net400),
    .Q_N(_0024_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ));
 sg13g2_dfrbp_1 _4437_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net248),
    .D(net639),
    .Q_N(_2120_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ));
 sg13g2_dfrbp_1 _4438_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net246),
    .D(net462),
    .Q_N(_2119_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[0] ));
 sg13g2_dfrbp_1 _4439_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net245),
    .D(_0097_),
    .Q_N(_2118_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[1] ));
 sg13g2_dfrbp_1 _4440_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net244),
    .D(_0098_),
    .Q_N(_2117_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[2] ));
 sg13g2_dfrbp_1 _4441_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net243),
    .D(_0099_),
    .Q_N(_2116_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[3] ));
 sg13g2_dfrbp_1 _4442_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net242),
    .D(_0100_),
    .Q_N(_2115_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[4] ));
 sg13g2_dfrbp_1 _4443_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net241),
    .D(net447),
    .Q_N(_2114_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[5] ));
 sg13g2_dfrbp_1 _4444_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net240),
    .D(_0102_),
    .Q_N(_2113_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[6] ));
 sg13g2_dfrbp_1 _4445_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net239),
    .D(net519),
    .Q_N(_2112_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[7] ));
 sg13g2_dfrbp_1 _4446_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net238),
    .D(_0104_),
    .Q_N(_2111_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.last_ram_a_sel ));
 sg13g2_dfrbp_1 _4447_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net237),
    .D(_0105_),
    .Q_N(_2110_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.stop_txn ));
 sg13g2_dfrbp_1 _4448_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net236),
    .D(_0106_),
    .Q_N(_2109_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ));
 sg13g2_dfrbp_1 _4449_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net235),
    .D(_0107_),
    .Q_N(_2108_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[1] ));
 sg13g2_dfrbp_1 _4450_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net234),
    .D(_0108_),
    .Q_N(_2107_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[0] ));
 sg13g2_dfrbp_1 _4451_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net233),
    .D(_0109_),
    .Q_N(_2106_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[1] ));
 sg13g2_dfrbp_1 _4452_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net232),
    .D(_0110_),
    .Q_N(_2105_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[2] ));
 sg13g2_dfrbp_1 _4453_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net231),
    .D(_0111_),
    .Q_N(_2104_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[3] ));
 sg13g2_dfrbp_1 _4454_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net230),
    .D(_0112_),
    .Q_N(_2103_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[4] ));
 sg13g2_dfrbp_1 _4455_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net229),
    .D(_0113_),
    .Q_N(_2102_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[5] ));
 sg13g2_dfrbp_1 _4456_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net228),
    .D(_0114_),
    .Q_N(_2101_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[6] ));
 sg13g2_dfrbp_1 _4457_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net227),
    .D(_0115_),
    .Q_N(_2100_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[7] ));
 sg13g2_dfrbp_1 _4458_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net226),
    .D(net343),
    .Q_N(_2099_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[8] ));
 sg13g2_dfrbp_1 _4459_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net225),
    .D(_0117_),
    .Q_N(_2098_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[9] ));
 sg13g2_dfrbp_1 _4460_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net224),
    .D(_0118_),
    .Q_N(_2097_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[10] ));
 sg13g2_dfrbp_1 _4461_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net223),
    .D(_0119_),
    .Q_N(_2096_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[11] ));
 sg13g2_dfrbp_1 _4462_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net222),
    .D(net353),
    .Q_N(_2095_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ));
 sg13g2_dfrbp_1 _4463_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net221),
    .D(_0121_),
    .Q_N(_2094_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[13] ));
 sg13g2_dfrbp_1 _4464_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net220),
    .D(_0122_),
    .Q_N(_2093_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[14] ));
 sg13g2_dfrbp_1 _4465_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net219),
    .D(_0123_),
    .Q_N(_2092_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[15] ));
 sg13g2_dfrbp_1 _4466_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net218),
    .D(net325),
    .Q_N(_0015_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ));
 sg13g2_dfrbp_1 _4467_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net217),
    .D(_0125_),
    .Q_N(_2091_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.start_write ));
 sg13g2_dfrbp_1 _4468_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net216),
    .D(net652),
    .Q_N(_2090_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.start_read ));
 sg13g2_dfrbp_1 _4469_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net215),
    .D(_0127_),
    .Q_N(_0000_),
    .Q(\cpu_instance.ctrl_instance.mem_op_done ));
 sg13g2_dfrbp_1 _4470_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net214),
    .D(_0128_),
    .Q_N(_2089_),
    .Q(\cpu_instance.mem_instance.bus_data_out[0] ));
 sg13g2_dfrbp_1 _4471_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net212),
    .D(_0129_),
    .Q_N(_2088_),
    .Q(\cpu_instance.mem_instance.bus_data_out[1] ));
 sg13g2_dfrbp_1 _4472_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net210),
    .D(_0130_),
    .Q_N(_2087_),
    .Q(\cpu_instance.mem_instance.bus_data_out[2] ));
 sg13g2_dfrbp_1 _4473_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net208),
    .D(net571),
    .Q_N(_2086_),
    .Q(\cpu_instance.mem_instance.bus_data_out[3] ));
 sg13g2_dfrbp_1 _4474_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net206),
    .D(_0132_),
    .Q_N(_2085_),
    .Q(\cpu_instance.mem_instance.bus_data_out[4] ));
 sg13g2_dfrbp_1 _4475_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net204),
    .D(_0133_),
    .Q_N(_2084_),
    .Q(\cpu_instance.mem_instance.bus_data_out[5] ));
 sg13g2_dfrbp_1 _4476_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net202),
    .D(_0134_),
    .Q_N(_2083_),
    .Q(\cpu_instance.mem_instance.bus_data_out[6] ));
 sg13g2_dfrbp_1 _4477_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net200),
    .D(_0135_),
    .Q_N(_2082_),
    .Q(\cpu_instance.mem_instance.bus_data_out[7] ));
 sg13g2_dfrbp_1 _4478_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net198),
    .D(_0136_),
    .Q_N(_2081_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ));
 sg13g2_dfrbp_1 _4479_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net197),
    .D(_0137_),
    .Q_N(_2080_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ));
 sg13g2_dfrbp_1 _4480_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net196),
    .D(_0138_),
    .Q_N(_2079_),
    .Q(\cpu_instance.reg_2_out_sel[0] ));
 sg13g2_dfrbp_1 _4481_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net195),
    .D(_0139_),
    .Q_N(_2078_),
    .Q(\cpu_instance.reg_2_out_sel[1] ));
 sg13g2_dfrbp_1 _4482_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net194),
    .D(_0140_),
    .Q_N(_2077_),
    .Q(\cpu_instance.ctrl_instance.scan_in ));
 sg13g2_dfrbp_1 _4483_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net192),
    .D(_0141_),
    .Q_N(_2076_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[1] ));
 sg13g2_dfrbp_1 _4484_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net190),
    .D(net421),
    .Q_N(_2075_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[2] ));
 sg13g2_dfrbp_1 _4485_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net188),
    .D(_0143_),
    .Q_N(_2074_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[3] ));
 sg13g2_dfrbp_1 _4486_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net186),
    .D(net425),
    .Q_N(_2073_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[4] ));
 sg13g2_dfrbp_1 _4487_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net184),
    .D(_0145_),
    .Q_N(_2072_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[5] ));
 sg13g2_dfrbp_1 _4488_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net182),
    .D(_0146_),
    .Q_N(_2071_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[6] ));
 sg13g2_dfrbp_1 _4489_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net180),
    .D(net373),
    .Q_N(_2070_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[7] ));
 sg13g2_dfrbp_1 _4490_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net178),
    .D(net416),
    .Q_N(_2069_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ));
 sg13g2_dfrbp_1 _4491_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net176),
    .D(_0149_),
    .Q_N(_2068_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ));
 sg13g2_dfrbp_1 _4492_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net174),
    .D(net347),
    .Q_N(_2067_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ));
 sg13g2_dfrbp_1 _4493_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net172),
    .D(_0151_),
    .Q_N(_2066_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ));
 sg13g2_dfrbp_1 _4494_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net170),
    .D(net341),
    .Q_N(_2065_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][4] ));
 sg13g2_dfrbp_1 _4495_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net168),
    .D(_0153_),
    .Q_N(_2064_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ));
 sg13g2_dfrbp_1 _4496_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net166),
    .D(net345),
    .Q_N(_2063_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][6] ));
 sg13g2_dfrbp_1 _4497_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net164),
    .D(_0155_),
    .Q_N(_2062_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ));
 sg13g2_dfrbp_1 _4498_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net162),
    .D(_0156_),
    .Q_N(_2061_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ));
 sg13g2_dfrbp_1 _4499_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net160),
    .D(_0157_),
    .Q_N(_2060_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ));
 sg13g2_dfrbp_1 _4500_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net158),
    .D(net355),
    .Q_N(_2059_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][10] ));
 sg13g2_dfrbp_1 _4501_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net156),
    .D(_0159_),
    .Q_N(_2058_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ));
 sg13g2_dfrbp_1 _4502_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net154),
    .D(net360),
    .Q_N(_2057_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ));
 sg13g2_dfrbp_1 _4503_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net152),
    .D(_0161_),
    .Q_N(_2056_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ));
 sg13g2_dfrbp_1 _4504_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net150),
    .D(_0162_),
    .Q_N(_2055_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ));
 sg13g2_dfrbp_1 _4505_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net148),
    .D(_0163_),
    .Q_N(_2054_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ));
 sg13g2_dfrbp_1 _4506_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net146),
    .D(_0164_),
    .Q_N(_2053_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ));
 sg13g2_dfrbp_1 _4507_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net144),
    .D(_0165_),
    .Q_N(_2052_),
    .Q(\cpu_instance.registers_instance.register_bank[15][0] ));
 sg13g2_dfrbp_1 _4508_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net142),
    .D(_0166_),
    .Q_N(_2051_),
    .Q(\cpu_instance.registers_instance.register_bank[15][1] ));
 sg13g2_dfrbp_1 _4509_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net140),
    .D(_0167_),
    .Q_N(_2050_),
    .Q(\cpu_instance.registers_instance.register_bank[15][2] ));
 sg13g2_dfrbp_1 _4510_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net138),
    .D(_0168_),
    .Q_N(_2049_),
    .Q(\cpu_instance.registers_instance.register_bank[15][3] ));
 sg13g2_dfrbp_1 _4511_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net136),
    .D(_0169_),
    .Q_N(_2048_),
    .Q(\cpu_instance.registers_instance.register_bank[15][4] ));
 sg13g2_dfrbp_1 _4512_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net134),
    .D(_0170_),
    .Q_N(_2047_),
    .Q(\cpu_instance.registers_instance.register_bank[15][5] ));
 sg13g2_dfrbp_1 _4513_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net132),
    .D(_0171_),
    .Q_N(_2046_),
    .Q(\cpu_instance.registers_instance.register_bank[15][6] ));
 sg13g2_dfrbp_1 _4514_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net130),
    .D(_0172_),
    .Q_N(_2045_),
    .Q(\cpu_instance.registers_instance.register_bank[15][7] ));
 sg13g2_dfrbp_1 _4515_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net128),
    .D(net521),
    .Q_N(_0018_),
    .Q(\cpu_instance.registers_instance.registers[0][0] ));
 sg13g2_dfrbp_1 _4516_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net126),
    .D(_0174_),
    .Q_N(_0019_),
    .Q(\cpu_instance.registers_instance.registers[0][1] ));
 sg13g2_dfrbp_1 _4517_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net124),
    .D(_0175_),
    .Q_N(_0005_),
    .Q(\cpu_instance.registers_instance.registers[0][2] ));
 sg13g2_dfrbp_1 _4518_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net122),
    .D(net436),
    .Q_N(_0020_),
    .Q(\cpu_instance.registers_instance.registers[0][3] ));
 sg13g2_dfrbp_1 _4519_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net120),
    .D(_0177_),
    .Q_N(_0003_),
    .Q(\cpu_instance.registers_instance.registers[0][4] ));
 sg13g2_dfrbp_1 _4520_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net118),
    .D(net375),
    .Q_N(_0008_),
    .Q(\cpu_instance.registers_instance.registers[0][5] ));
 sg13g2_dfrbp_1 _4521_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net116),
    .D(_0179_),
    .Q_N(_0009_),
    .Q(\cpu_instance.registers_instance.registers[0][6] ));
 sg13g2_dfrbp_1 _4522_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net114),
    .D(_0180_),
    .Q_N(_0012_),
    .Q(\cpu_instance.registers_instance.registers[0][7] ));
 sg13g2_dfrbp_1 _4523_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net112),
    .D(_0181_),
    .Q_N(_2044_),
    .Q(\cpu_instance.registers_instance.registers[1][0] ));
 sg13g2_dfrbp_1 _4524_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net110),
    .D(_0182_),
    .Q_N(_2043_),
    .Q(\cpu_instance.registers_instance.registers[1][1] ));
 sg13g2_dfrbp_1 _4525_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net108),
    .D(net588),
    .Q_N(_2042_),
    .Q(\cpu_instance.registers_instance.registers[1][2] ));
 sg13g2_dfrbp_1 _4526_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net106),
    .D(_0184_),
    .Q_N(_2041_),
    .Q(\cpu_instance.registers_instance.registers[1][3] ));
 sg13g2_dfrbp_1 _4527_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net104),
    .D(net606),
    .Q_N(_2040_),
    .Q(\cpu_instance.registers_instance.registers[1][4] ));
 sg13g2_dfrbp_1 _4528_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net102),
    .D(net531),
    .Q_N(_2039_),
    .Q(\cpu_instance.registers_instance.registers[1][5] ));
 sg13g2_dfrbp_1 _4529_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net100),
    .D(_0187_),
    .Q_N(_2038_),
    .Q(\cpu_instance.registers_instance.registers[1][6] ));
 sg13g2_dfrbp_1 _4530_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net98),
    .D(_0188_),
    .Q_N(_2037_),
    .Q(\cpu_instance.registers_instance.registers[1][7] ));
 sg13g2_dfrbp_1 _4531_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net96),
    .D(net580),
    .Q_N(_2036_),
    .Q(\cpu_instance.registers_instance.registers[2][0] ));
 sg13g2_dfrbp_1 _4532_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net94),
    .D(_0190_),
    .Q_N(_2035_),
    .Q(\cpu_instance.registers_instance.registers[2][1] ));
 sg13g2_dfrbp_1 _4533_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net92),
    .D(net618),
    .Q_N(_2034_),
    .Q(\cpu_instance.registers_instance.registers[2][2] ));
 sg13g2_dfrbp_1 _4534_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net90),
    .D(_0192_),
    .Q_N(_2033_),
    .Q(\cpu_instance.registers_instance.registers[2][3] ));
 sg13g2_dfrbp_1 _4535_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net88),
    .D(_0193_),
    .Q_N(_2032_),
    .Q(\cpu_instance.registers_instance.registers[2][4] ));
 sg13g2_dfrbp_1 _4536_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net86),
    .D(_0194_),
    .Q_N(_2031_),
    .Q(\cpu_instance.registers_instance.registers[2][5] ));
 sg13g2_dfrbp_1 _4537_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net84),
    .D(net558),
    .Q_N(_2030_),
    .Q(\cpu_instance.registers_instance.registers[2][6] ));
 sg13g2_dfrbp_1 _4538_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net82),
    .D(net319),
    .Q_N(_2029_),
    .Q(\cpu_instance.registers_instance.registers[2][7] ));
 sg13g2_dfrbp_1 _4539_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net80),
    .D(net654),
    .Q_N(_0001_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _4540_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net78),
    .D(_0198_),
    .Q_N(_0002_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _4541_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net76),
    .D(_0199_),
    .Q_N(_2028_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _4542_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net74),
    .D(net584),
    .Q_N(_0021_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _4543_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net72),
    .D(_0201_),
    .Q_N(_2027_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _4544_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net70),
    .D(_0202_),
    .Q_N(_2026_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _4545_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net68),
    .D(net620),
    .Q_N(_0010_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _4546_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net66),
    .D(net632),
    .Q_N(_0013_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _4547_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net62),
    .D(net569),
    .Q_N(_0007_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ));
 sg13g2_dfrbp_1 _4548_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net58),
    .D(_0206_),
    .Q_N(_0006_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ));
 sg13g2_dfrbp_1 _4549_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net54),
    .D(net578),
    .Q_N(_0004_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ));
 sg13g2_dfrbp_1 _4550_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net48),
    .D(net644),
    .Q_N(_2025_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ));
 sg13g2_dfrbp_1 _4551_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net44),
    .D(_0209_),
    .Q_N(_2024_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ));
 sg13g2_dfrbp_1 _4552_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net38),
    .D(_0210_),
    .Q_N(_2023_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ));
 sg13g2_dfrbp_1 _4553_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net34),
    .D(net586),
    .Q_N(_0011_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ));
 sg13g2_dfrbp_1 _4554_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net30),
    .D(net626),
    .Q_N(_0014_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ));
 sg13g2_dfrbp_1 _4555_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net26),
    .D(_0213_),
    .Q_N(_2022_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ));
 sg13g2_dfrbp_1 _4556_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net16),
    .D(net612),
    .Q_N(_2021_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ));
 sg13g2_dfrbp_1 _4557_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net12),
    .D(_0215_),
    .Q_N(_2020_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ));
 sg13g2_dfrbp_1 _4558_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net305),
    .D(_0216_),
    .Q_N(_2019_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ));
 sg13g2_dfrbp_1 _4559_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net301),
    .D(net593),
    .Q_N(_2018_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ));
 sg13g2_dfrbp_1 _4560_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net297),
    .D(_0218_),
    .Q_N(_2017_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ));
 sg13g2_dfrbp_1 _4561_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net293),
    .D(_0219_),
    .Q_N(_2016_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ));
 sg13g2_dfrbp_1 _4562_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net289),
    .D(net455),
    .Q_N(_2015_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ));
 sg13g2_dfrbp_1 _4563_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net285),
    .D(net457),
    .Q_N(_2014_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ));
 sg13g2_dfrbp_1 _4564_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net281),
    .D(net491),
    .Q_N(_2013_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ));
 sg13g2_dfrbp_1 _4565_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net277),
    .D(_0223_),
    .Q_N(_2012_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ));
 sg13g2_dfrbp_1 _4566_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net270),
    .D(net502),
    .Q_N(_2011_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ));
 sg13g2_dfrbp_1 _4567_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net261),
    .D(_0225_),
    .Q_N(_2010_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ));
 sg13g2_dfrbp_1 _4568_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net257),
    .D(net534),
    .Q_N(_2009_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ));
 sg13g2_dfrbp_1 _4569_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net253),
    .D(net507),
    .Q_N(_2008_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ));
 sg13g2_dfrbp_1 _4570_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net249),
    .D(_0228_),
    .Q_N(_2007_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ));
 sg13g2_dfrbp_1 _4571_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net213),
    .D(_0229_),
    .Q_N(_2006_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ));
 sg13g2_dfrbp_1 _4572_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net209),
    .D(net497),
    .Q_N(_2005_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ));
 sg13g2_dfrbp_1 _4573_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net205),
    .D(_0231_),
    .Q_N(_2004_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ));
 sg13g2_dfrbp_1 _4574_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net201),
    .D(_0232_),
    .Q_N(_2003_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ));
 sg13g2_dfrbp_1 _4575_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net193),
    .D(_0233_),
    .Q_N(_2002_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ));
 sg13g2_dfrbp_1 _4576_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net189),
    .D(_0234_),
    .Q_N(_2001_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ));
 sg13g2_dfrbp_1 _4577_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net185),
    .D(net528),
    .Q_N(_2000_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ));
 sg13g2_dfrbp_1 _4578_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net181),
    .D(_0236_),
    .Q_N(_1999_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ));
 sg13g2_dfrbp_1 _4579_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net177),
    .D(net556),
    .Q_N(_1998_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ));
 sg13g2_dfrbp_1 _4580_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net173),
    .D(net526),
    .Q_N(_1997_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ));
 sg13g2_dfrbp_1 _4581_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net169),
    .D(_0239_),
    .Q_N(_1996_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ));
 sg13g2_dfrbp_1 _4582_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net165),
    .D(_0240_),
    .Q_N(_1995_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ));
 sg13g2_dfrbp_1 _4583_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net161),
    .D(net504),
    .Q_N(_1994_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ));
 sg13g2_dfrbp_1 _4584_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net157),
    .D(net516),
    .Q_N(_1993_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ));
 sg13g2_dfrbp_1 _4585_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net153),
    .D(_0243_),
    .Q_N(_1992_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ));
 sg13g2_dfrbp_1 _4586_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net149),
    .D(net470),
    .Q_N(_1991_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ));
 sg13g2_dfrbp_1 _4587_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net145),
    .D(_0245_),
    .Q_N(_1990_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ));
 sg13g2_dfrbp_1 _4588_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net141),
    .D(_0246_),
    .Q_N(_1989_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ));
 sg13g2_dfrbp_1 _4589_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net137),
    .D(net481),
    .Q_N(_1988_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ));
 sg13g2_dfrbp_1 _4590_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net133),
    .D(net546),
    .Q_N(_1987_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ));
 sg13g2_dfrbp_1 _4591_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net129),
    .D(_0249_),
    .Q_N(_1986_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ));
 sg13g2_dfrbp_1 _4592_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net125),
    .D(net483),
    .Q_N(_1985_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ));
 sg13g2_dfrbp_1 _4593_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net121),
    .D(_0251_),
    .Q_N(_1984_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ));
 sg13g2_dfrbp_1 _4594_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net117),
    .D(net476),
    .Q_N(_1983_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ));
 sg13g2_dfrbp_1 _4595_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net113),
    .D(_0253_),
    .Q_N(_1982_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ));
 sg13g2_dfrbp_1 _4596_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net109),
    .D(_0254_),
    .Q_N(_1981_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ));
 sg13g2_dfrbp_1 _4597_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net105),
    .D(_0255_),
    .Q_N(_1980_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ));
 sg13g2_dfrbp_1 _4598_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net101),
    .D(_0256_),
    .Q_N(_1979_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ));
 sg13g2_dfrbp_1 _4599_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net97),
    .D(_0257_),
    .Q_N(_1978_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ));
 sg13g2_dfrbp_1 _4600_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net93),
    .D(net479),
    .Q_N(_1977_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ));
 sg13g2_dfrbp_1 _4601_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net89),
    .D(net509),
    .Q_N(_1976_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ));
 sg13g2_dfrbp_1 _4602_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net85),
    .D(_0260_),
    .Q_N(_1975_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ));
 sg13g2_dfrbp_1 _4603_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net81),
    .D(_0261_),
    .Q_N(_1974_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ));
 sg13g2_dfrbp_1 _4604_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net77),
    .D(net494),
    .Q_N(_1973_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ));
 sg13g2_dfrbp_1 _4605_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net73),
    .D(net371),
    .Q_N(_1972_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ));
 sg13g2_dfrbp_1 _4606_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net69),
    .D(_0264_),
    .Q_N(_1971_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ));
 sg13g2_dfrbp_1 _4607_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net64),
    .D(_0265_),
    .Q_N(_1970_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ));
 sg13g2_dfrbp_1 _4608_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net56),
    .D(net513),
    .Q_N(_1969_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ));
 sg13g2_dfrbp_1 _4609_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net46),
    .D(net524),
    .Q_N(_1968_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ));
 sg13g2_dfrbp_1 _4610_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net36),
    .D(net488),
    .Q_N(_1967_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ));
 sg13g2_dfrbp_1 _4611_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net28),
    .D(_0269_),
    .Q_N(_1966_),
    .Q(\cpu_instance.registers_instance.register_bank[8][0] ));
 sg13g2_dfrbp_1 _4612_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net14),
    .D(_0270_),
    .Q_N(_1965_),
    .Q(\cpu_instance.registers_instance.register_bank[8][1] ));
 sg13g2_dfrbp_1 _4613_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net303),
    .D(_0271_),
    .Q_N(_1964_),
    .Q(\cpu_instance.registers_instance.register_bank[8][2] ));
 sg13g2_dfrbp_1 _4614_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net295),
    .D(_0272_),
    .Q_N(_1963_),
    .Q(\cpu_instance.registers_instance.register_bank[8][3] ));
 sg13g2_dfrbp_1 _4615_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net287),
    .D(_0273_),
    .Q_N(_1962_),
    .Q(\cpu_instance.registers_instance.register_bank[8][4] ));
 sg13g2_dfrbp_1 _4616_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net279),
    .D(_0274_),
    .Q_N(_1961_),
    .Q(\cpu_instance.registers_instance.register_bank[8][5] ));
 sg13g2_dfrbp_1 _4617_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net268),
    .D(_0275_),
    .Q_N(_1960_),
    .Q(\cpu_instance.registers_instance.register_bank[8][6] ));
 sg13g2_dfrbp_1 _4618_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net255),
    .D(_0276_),
    .Q_N(_1959_),
    .Q(\cpu_instance.registers_instance.register_bank[8][7] ));
 sg13g2_dfrbp_1 _4619_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net247),
    .D(_0277_),
    .Q_N(_1958_),
    .Q(\cpu_instance.registers_instance.register_bank[9][0] ));
 sg13g2_dfrbp_1 _4620_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net207),
    .D(_0278_),
    .Q_N(_1957_),
    .Q(\cpu_instance.registers_instance.register_bank[9][1] ));
 sg13g2_dfrbp_1 _4621_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net199),
    .D(_0279_),
    .Q_N(_1956_),
    .Q(\cpu_instance.registers_instance.register_bank[9][2] ));
 sg13g2_dfrbp_1 _4622_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net187),
    .D(_0280_),
    .Q_N(_1955_),
    .Q(\cpu_instance.registers_instance.register_bank[9][3] ));
 sg13g2_dfrbp_1 _4623_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net179),
    .D(_0281_),
    .Q_N(_1954_),
    .Q(\cpu_instance.registers_instance.register_bank[9][4] ));
 sg13g2_dfrbp_1 _4624_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net171),
    .D(_0282_),
    .Q_N(_1953_),
    .Q(\cpu_instance.registers_instance.register_bank[9][5] ));
 sg13g2_dfrbp_1 _4625_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net163),
    .D(_0283_),
    .Q_N(_1952_),
    .Q(\cpu_instance.registers_instance.register_bank[9][6] ));
 sg13g2_dfrbp_1 _4626_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net155),
    .D(_0284_),
    .Q_N(_1951_),
    .Q(\cpu_instance.registers_instance.register_bank[9][7] ));
 sg13g2_dfrbp_1 _4627_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net147),
    .D(_0285_),
    .Q_N(_1950_),
    .Q(\cpu_instance.registers_instance.register_bank[10][0] ));
 sg13g2_dfrbp_1 _4628_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net139),
    .D(_0286_),
    .Q_N(_1949_),
    .Q(\cpu_instance.registers_instance.register_bank[10][1] ));
 sg13g2_dfrbp_1 _4629_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net131),
    .D(_0287_),
    .Q_N(_1948_),
    .Q(\cpu_instance.registers_instance.register_bank[10][2] ));
 sg13g2_dfrbp_1 _4630_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net123),
    .D(_0288_),
    .Q_N(_1947_),
    .Q(\cpu_instance.registers_instance.register_bank[10][3] ));
 sg13g2_dfrbp_1 _4631_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net115),
    .D(_0289_),
    .Q_N(_1946_),
    .Q(\cpu_instance.registers_instance.register_bank[10][4] ));
 sg13g2_dfrbp_1 _4632_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net107),
    .D(_0290_),
    .Q_N(_1945_),
    .Q(\cpu_instance.registers_instance.register_bank[10][5] ));
 sg13g2_dfrbp_1 _4633_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net99),
    .D(_0291_),
    .Q_N(_1944_),
    .Q(\cpu_instance.registers_instance.register_bank[10][6] ));
 sg13g2_dfrbp_1 _4634_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net91),
    .D(_0292_),
    .Q_N(_1943_),
    .Q(\cpu_instance.registers_instance.register_bank[10][7] ));
 sg13g2_dfrbp_1 _4635_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net83),
    .D(_0293_),
    .Q_N(_1942_),
    .Q(\cpu_instance.registers_instance.register_bank[11][0] ));
 sg13g2_dfrbp_1 _4636_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net75),
    .D(_0294_),
    .Q_N(_1941_),
    .Q(\cpu_instance.registers_instance.register_bank[11][1] ));
 sg13g2_dfrbp_1 _4637_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net67),
    .D(_0295_),
    .Q_N(_1940_),
    .Q(\cpu_instance.registers_instance.register_bank[11][2] ));
 sg13g2_dfrbp_1 _4638_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net50),
    .D(_0296_),
    .Q_N(_1939_),
    .Q(\cpu_instance.registers_instance.register_bank[11][3] ));
 sg13g2_dfrbp_1 _4639_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net32),
    .D(_0297_),
    .Q_N(_1938_),
    .Q(\cpu_instance.registers_instance.register_bank[11][4] ));
 sg13g2_dfrbp_1 _4640_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net307),
    .D(_0298_),
    .Q_N(_1937_),
    .Q(\cpu_instance.registers_instance.register_bank[11][5] ));
 sg13g2_dfrbp_1 _4641_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net291),
    .D(_0299_),
    .Q_N(_1936_),
    .Q(\cpu_instance.registers_instance.register_bank[11][6] ));
 sg13g2_dfrbp_1 _4642_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net272),
    .D(_0300_),
    .Q_N(_1935_),
    .Q(\cpu_instance.registers_instance.register_bank[11][7] ));
 sg13g2_dfrbp_1 _4643_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net251),
    .D(_0301_),
    .Q_N(_1934_),
    .Q(\cpu_instance.registers_instance.register_bank[12][0] ));
 sg13g2_dfrbp_1 _4644_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net203),
    .D(_0302_),
    .Q_N(_1933_),
    .Q(\cpu_instance.registers_instance.register_bank[12][1] ));
 sg13g2_dfrbp_1 _4645_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net183),
    .D(_0303_),
    .Q_N(_1932_),
    .Q(\cpu_instance.registers_instance.register_bank[12][2] ));
 sg13g2_dfrbp_1 _4646_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net167),
    .D(_0304_),
    .Q_N(_1931_),
    .Q(\cpu_instance.registers_instance.register_bank[12][3] ));
 sg13g2_dfrbp_1 _4647_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net151),
    .D(_0305_),
    .Q_N(_1930_),
    .Q(\cpu_instance.registers_instance.register_bank[12][4] ));
 sg13g2_dfrbp_1 _4648_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net135),
    .D(_0306_),
    .Q_N(_1929_),
    .Q(\cpu_instance.registers_instance.register_bank[12][5] ));
 sg13g2_dfrbp_1 _4649_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net119),
    .D(_0307_),
    .Q_N(_1928_),
    .Q(\cpu_instance.registers_instance.register_bank[12][6] ));
 sg13g2_dfrbp_1 _4650_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net103),
    .D(_0308_),
    .Q_N(_1927_),
    .Q(\cpu_instance.registers_instance.register_bank[12][7] ));
 sg13g2_dfrbp_1 _4651_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net87),
    .D(_0309_),
    .Q_N(_1926_),
    .Q(\cpu_instance.registers_instance.register_bank[13][0] ));
 sg13g2_dfrbp_1 _4652_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net71),
    .D(_0310_),
    .Q_N(_1925_),
    .Q(\cpu_instance.registers_instance.register_bank[13][1] ));
 sg13g2_dfrbp_1 _4653_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net40),
    .D(_0311_),
    .Q_N(_1924_),
    .Q(\cpu_instance.registers_instance.register_bank[13][2] ));
 sg13g2_dfrbp_1 _4654_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net299),
    .D(_0312_),
    .Q_N(_1923_),
    .Q(\cpu_instance.registers_instance.register_bank[13][3] ));
 sg13g2_dfrbp_1 _4655_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net259),
    .D(_0313_),
    .Q_N(_1922_),
    .Q(\cpu_instance.registers_instance.register_bank[13][4] ));
 sg13g2_dfrbp_1 _4656_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net191),
    .D(_0314_),
    .Q_N(_1921_),
    .Q(\cpu_instance.registers_instance.register_bank[13][5] ));
 sg13g2_dfrbp_1 _4657_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net159),
    .D(_0315_),
    .Q_N(_1920_),
    .Q(\cpu_instance.registers_instance.register_bank[13][6] ));
 sg13g2_dfrbp_1 _4658_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net127),
    .D(_0316_),
    .Q_N(_1919_),
    .Q(\cpu_instance.registers_instance.register_bank[13][7] ));
 sg13g2_dfrbp_1 _4659_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net95),
    .D(net551),
    .Q_N(_1918_),
    .Q(\cpu_instance.registers_instance.register_bank[14][0] ));
 sg13g2_dfrbp_1 _4660_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net60),
    .D(_0318_),
    .Q_N(_1917_),
    .Q(\cpu_instance.registers_instance.register_bank[14][1] ));
 sg13g2_dfrbp_1 _4661_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net283),
    .D(_0319_),
    .Q_N(_1916_),
    .Q(\cpu_instance.registers_instance.register_bank[14][2] ));
 sg13g2_dfrbp_1 _4662_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net175),
    .D(_0320_),
    .Q_N(_1915_),
    .Q(\cpu_instance.registers_instance.register_bank[14][3] ));
 sg13g2_dfrbp_1 _4663_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net111),
    .D(_0321_),
    .Q_N(_1914_),
    .Q(\cpu_instance.registers_instance.register_bank[14][4] ));
 sg13g2_dfrbp_1 _4664_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net18),
    .D(_0322_),
    .Q_N(_1913_),
    .Q(\cpu_instance.registers_instance.register_bank[14][5] ));
 sg13g2_dfrbp_1 _4665_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net143),
    .D(net466),
    .Q_N(_1912_),
    .Q(\cpu_instance.registers_instance.register_bank[14][6] ));
 sg13g2_dfrbp_1 _4666_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net211),
    .D(_0324_),
    .Q_N(_1911_),
    .Q(\cpu_instance.registers_instance.register_bank[14][7] ));
 sg13g2_tiehi _4401__13 (.L_HI(net13));
 sg13g2_tiehi _4612__14 (.L_HI(net14));
 sg13g2_tiehi _4400__15 (.L_HI(net15));
 sg13g2_tiehi _4556__16 (.L_HI(net16));
 sg13g2_tiehi _4399__17 (.L_HI(net17));
 sg13g2_tiehi _4664__18 (.L_HI(net18));
 sg13g2_tiehi _4398__19 (.L_HI(net19));
 sg13g2_tiehi _4397__20 (.L_HI(net20));
 sg13g2_tiehi _4396__21 (.L_HI(net21));
 sg13g2_tiehi _4395__22 (.L_HI(net22));
 sg13g2_tiehi _4394__23 (.L_HI(net23));
 sg13g2_tiehi _4393__24 (.L_HI(net24));
 sg13g2_tiehi _4392__25 (.L_HI(net25));
 sg13g2_tiehi _4555__26 (.L_HI(net26));
 sg13g2_tiehi _4391__27 (.L_HI(net27));
 sg13g2_tiehi _4611__28 (.L_HI(net28));
 sg13g2_tiehi _4390__29 (.L_HI(net29));
 sg13g2_tiehi _4554__30 (.L_HI(net30));
 sg13g2_tiehi _4389__31 (.L_HI(net31));
 sg13g2_tiehi _4639__32 (.L_HI(net32));
 sg13g2_tiehi _4388__33 (.L_HI(net33));
 sg13g2_tiehi _4553__34 (.L_HI(net34));
 sg13g2_tiehi _4387__35 (.L_HI(net35));
 sg13g2_tiehi _4610__36 (.L_HI(net36));
 sg13g2_tiehi _4386__37 (.L_HI(net37));
 sg13g2_tiehi _4552__38 (.L_HI(net38));
 sg13g2_tiehi _4385__39 (.L_HI(net39));
 sg13g2_tiehi _4653__40 (.L_HI(net40));
 sg13g2_tiehi _4384__41 (.L_HI(net41));
 sg13g2_tiehi _4383__42 (.L_HI(net42));
 sg13g2_tiehi _4382__43 (.L_HI(net43));
 sg13g2_tiehi _4551__44 (.L_HI(net44));
 sg13g2_tiehi _4381__45 (.L_HI(net45));
 sg13g2_tiehi _4609__46 (.L_HI(net46));
 sg13g2_tiehi _4380__47 (.L_HI(net47));
 sg13g2_tiehi _4550__48 (.L_HI(net48));
 sg13g2_tiehi _4379__49 (.L_HI(net49));
 sg13g2_tiehi _4638__50 (.L_HI(net50));
 sg13g2_tiehi _4378__51 (.L_HI(net51));
 sg13g2_tiehi _4377__52 (.L_HI(net52));
 sg13g2_tiehi _4376__53 (.L_HI(net53));
 sg13g2_tiehi _4549__54 (.L_HI(net54));
 sg13g2_tiehi _4375__55 (.L_HI(net55));
 sg13g2_tiehi _4608__56 (.L_HI(net56));
 sg13g2_tiehi _4374__57 (.L_HI(net57));
 sg13g2_tiehi _4548__58 (.L_HI(net58));
 sg13g2_tiehi _4373__59 (.L_HI(net59));
 sg13g2_tiehi _4660__60 (.L_HI(net60));
 sg13g2_tiehi _4372__61 (.L_HI(net61));
 sg13g2_tiehi _4547__62 (.L_HI(net62));
 sg13g2_tiehi _4371__63 (.L_HI(net63));
 sg13g2_tiehi _4607__64 (.L_HI(net64));
 sg13g2_tiehi _4370__65 (.L_HI(net65));
 sg13g2_tiehi _4546__66 (.L_HI(net66));
 sg13g2_tiehi _4637__67 (.L_HI(net67));
 sg13g2_tiehi _4545__68 (.L_HI(net68));
 sg13g2_tiehi _4606__69 (.L_HI(net69));
 sg13g2_tiehi _4544__70 (.L_HI(net70));
 sg13g2_tiehi _4652__71 (.L_HI(net71));
 sg13g2_tiehi _4543__72 (.L_HI(net72));
 sg13g2_tiehi _4605__73 (.L_HI(net73));
 sg13g2_tiehi _4542__74 (.L_HI(net74));
 sg13g2_tiehi _4636__75 (.L_HI(net75));
 sg13g2_tiehi _4541__76 (.L_HI(net76));
 sg13g2_tiehi _4604__77 (.L_HI(net77));
 sg13g2_tiehi _4540__78 (.L_HI(net78));
 sg13g2_tiehi _4369__79 (.L_HI(net79));
 sg13g2_tiehi _4539__80 (.L_HI(net80));
 sg13g2_tiehi _4603__81 (.L_HI(net81));
 sg13g2_tiehi _4538__82 (.L_HI(net82));
 sg13g2_tiehi _4635__83 (.L_HI(net83));
 sg13g2_tiehi _4537__84 (.L_HI(net84));
 sg13g2_tiehi _4602__85 (.L_HI(net85));
 sg13g2_tiehi _4536__86 (.L_HI(net86));
 sg13g2_tiehi _4651__87 (.L_HI(net87));
 sg13g2_tiehi _4535__88 (.L_HI(net88));
 sg13g2_tiehi _4601__89 (.L_HI(net89));
 sg13g2_tiehi _4534__90 (.L_HI(net90));
 sg13g2_tiehi _4634__91 (.L_HI(net91));
 sg13g2_tiehi _4533__92 (.L_HI(net92));
 sg13g2_tiehi _4600__93 (.L_HI(net93));
 sg13g2_tiehi _4532__94 (.L_HI(net94));
 sg13g2_tiehi _4659__95 (.L_HI(net95));
 sg13g2_tiehi _4531__96 (.L_HI(net96));
 sg13g2_tiehi _4599__97 (.L_HI(net97));
 sg13g2_tiehi _4530__98 (.L_HI(net98));
 sg13g2_tiehi _4633__99 (.L_HI(net99));
 sg13g2_tiehi _4529__100 (.L_HI(net100));
 sg13g2_tiehi _4598__101 (.L_HI(net101));
 sg13g2_tiehi _4528__102 (.L_HI(net102));
 sg13g2_tiehi _4650__103 (.L_HI(net103));
 sg13g2_tiehi _4527__104 (.L_HI(net104));
 sg13g2_tiehi _4597__105 (.L_HI(net105));
 sg13g2_tiehi _4526__106 (.L_HI(net106));
 sg13g2_tiehi _4632__107 (.L_HI(net107));
 sg13g2_tiehi _4525__108 (.L_HI(net108));
 sg13g2_tiehi _4596__109 (.L_HI(net109));
 sg13g2_tiehi _4524__110 (.L_HI(net110));
 sg13g2_tiehi _4663__111 (.L_HI(net111));
 sg13g2_tiehi _4523__112 (.L_HI(net112));
 sg13g2_tiehi _4595__113 (.L_HI(net113));
 sg13g2_tiehi _4522__114 (.L_HI(net114));
 sg13g2_tiehi _4631__115 (.L_HI(net115));
 sg13g2_tiehi _4521__116 (.L_HI(net116));
 sg13g2_tiehi _4594__117 (.L_HI(net117));
 sg13g2_tiehi _4520__118 (.L_HI(net118));
 sg13g2_tiehi _4649__119 (.L_HI(net119));
 sg13g2_tiehi _4519__120 (.L_HI(net120));
 sg13g2_tiehi _4593__121 (.L_HI(net121));
 sg13g2_tiehi _4518__122 (.L_HI(net122));
 sg13g2_tiehi _4630__123 (.L_HI(net123));
 sg13g2_tiehi _4517__124 (.L_HI(net124));
 sg13g2_tiehi _4592__125 (.L_HI(net125));
 sg13g2_tiehi _4516__126 (.L_HI(net126));
 sg13g2_tiehi _4658__127 (.L_HI(net127));
 sg13g2_tiehi _4515__128 (.L_HI(net128));
 sg13g2_tiehi _4591__129 (.L_HI(net129));
 sg13g2_tiehi _4514__130 (.L_HI(net130));
 sg13g2_tiehi _4629__131 (.L_HI(net131));
 sg13g2_tiehi _4513__132 (.L_HI(net132));
 sg13g2_tiehi _4590__133 (.L_HI(net133));
 sg13g2_tiehi _4512__134 (.L_HI(net134));
 sg13g2_tiehi _4648__135 (.L_HI(net135));
 sg13g2_tiehi _4511__136 (.L_HI(net136));
 sg13g2_tiehi _4589__137 (.L_HI(net137));
 sg13g2_tiehi _4510__138 (.L_HI(net138));
 sg13g2_tiehi _4628__139 (.L_HI(net139));
 sg13g2_tiehi _4509__140 (.L_HI(net140));
 sg13g2_tiehi _4588__141 (.L_HI(net141));
 sg13g2_tiehi _4508__142 (.L_HI(net142));
 sg13g2_tiehi _4665__143 (.L_HI(net143));
 sg13g2_tiehi _4507__144 (.L_HI(net144));
 sg13g2_tiehi _4587__145 (.L_HI(net145));
 sg13g2_tiehi _4506__146 (.L_HI(net146));
 sg13g2_tiehi _4627__147 (.L_HI(net147));
 sg13g2_tiehi _4505__148 (.L_HI(net148));
 sg13g2_tiehi _4586__149 (.L_HI(net149));
 sg13g2_tiehi _4504__150 (.L_HI(net150));
 sg13g2_tiehi _4647__151 (.L_HI(net151));
 sg13g2_tiehi _4503__152 (.L_HI(net152));
 sg13g2_tiehi _4585__153 (.L_HI(net153));
 sg13g2_tiehi _4502__154 (.L_HI(net154));
 sg13g2_tiehi _4626__155 (.L_HI(net155));
 sg13g2_tiehi _4501__156 (.L_HI(net156));
 sg13g2_tiehi _4584__157 (.L_HI(net157));
 sg13g2_tiehi _4500__158 (.L_HI(net158));
 sg13g2_tiehi _4657__159 (.L_HI(net159));
 sg13g2_tiehi _4499__160 (.L_HI(net160));
 sg13g2_tiehi _4583__161 (.L_HI(net161));
 sg13g2_tiehi _4498__162 (.L_HI(net162));
 sg13g2_tiehi _4625__163 (.L_HI(net163));
 sg13g2_tiehi _4497__164 (.L_HI(net164));
 sg13g2_tiehi _4582__165 (.L_HI(net165));
 sg13g2_tiehi _4496__166 (.L_HI(net166));
 sg13g2_tiehi _4646__167 (.L_HI(net167));
 sg13g2_tiehi _4495__168 (.L_HI(net168));
 sg13g2_tiehi _4581__169 (.L_HI(net169));
 sg13g2_tiehi _4494__170 (.L_HI(net170));
 sg13g2_tiehi _4624__171 (.L_HI(net171));
 sg13g2_tiehi _4493__172 (.L_HI(net172));
 sg13g2_tiehi _4580__173 (.L_HI(net173));
 sg13g2_tiehi _4492__174 (.L_HI(net174));
 sg13g2_tiehi _4662__175 (.L_HI(net175));
 sg13g2_tiehi _4491__176 (.L_HI(net176));
 sg13g2_tiehi _4579__177 (.L_HI(net177));
 sg13g2_tiehi _4490__178 (.L_HI(net178));
 sg13g2_tiehi _4623__179 (.L_HI(net179));
 sg13g2_tiehi _4489__180 (.L_HI(net180));
 sg13g2_tiehi _4578__181 (.L_HI(net181));
 sg13g2_tiehi _4488__182 (.L_HI(net182));
 sg13g2_tiehi _4645__183 (.L_HI(net183));
 sg13g2_tiehi _4487__184 (.L_HI(net184));
 sg13g2_tiehi _4577__185 (.L_HI(net185));
 sg13g2_tiehi _4486__186 (.L_HI(net186));
 sg13g2_tiehi _4622__187 (.L_HI(net187));
 sg13g2_tiehi _4485__188 (.L_HI(net188));
 sg13g2_tiehi _4576__189 (.L_HI(net189));
 sg13g2_tiehi _4484__190 (.L_HI(net190));
 sg13g2_tiehi _4656__191 (.L_HI(net191));
 sg13g2_tiehi _4483__192 (.L_HI(net192));
 sg13g2_tiehi _4575__193 (.L_HI(net193));
 sg13g2_tiehi _4482__194 (.L_HI(net194));
 sg13g2_tiehi _4481__195 (.L_HI(net195));
 sg13g2_tiehi _4480__196 (.L_HI(net196));
 sg13g2_tiehi _4479__197 (.L_HI(net197));
 sg13g2_tiehi _4478__198 (.L_HI(net198));
 sg13g2_tiehi _4621__199 (.L_HI(net199));
 sg13g2_tiehi _4477__200 (.L_HI(net200));
 sg13g2_tiehi _4574__201 (.L_HI(net201));
 sg13g2_tiehi _4476__202 (.L_HI(net202));
 sg13g2_tiehi _4644__203 (.L_HI(net203));
 sg13g2_tiehi _4475__204 (.L_HI(net204));
 sg13g2_tiehi _4573__205 (.L_HI(net205));
 sg13g2_tiehi _4474__206 (.L_HI(net206));
 sg13g2_tiehi _4620__207 (.L_HI(net207));
 sg13g2_tiehi _4473__208 (.L_HI(net208));
 sg13g2_tiehi _4572__209 (.L_HI(net209));
 sg13g2_tiehi _4472__210 (.L_HI(net210));
 sg13g2_tiehi _4666__211 (.L_HI(net211));
 sg13g2_tiehi _4471__212 (.L_HI(net212));
 sg13g2_tiehi _4571__213 (.L_HI(net213));
 sg13g2_tiehi _4470__214 (.L_HI(net214));
 sg13g2_tiehi _4469__215 (.L_HI(net215));
 sg13g2_tiehi _4468__216 (.L_HI(net216));
 sg13g2_tiehi _4467__217 (.L_HI(net217));
 sg13g2_tiehi _4466__218 (.L_HI(net218));
 sg13g2_tiehi _4465__219 (.L_HI(net219));
 sg13g2_tiehi _4464__220 (.L_HI(net220));
 sg13g2_tiehi _4463__221 (.L_HI(net221));
 sg13g2_tiehi _4462__222 (.L_HI(net222));
 sg13g2_tiehi _4461__223 (.L_HI(net223));
 sg13g2_tiehi _4460__224 (.L_HI(net224));
 sg13g2_tiehi _4459__225 (.L_HI(net225));
 sg13g2_tiehi _4458__226 (.L_HI(net226));
 sg13g2_tiehi _4457__227 (.L_HI(net227));
 sg13g2_tiehi _4456__228 (.L_HI(net228));
 sg13g2_tiehi _4455__229 (.L_HI(net229));
 sg13g2_tiehi _4454__230 (.L_HI(net230));
 sg13g2_tiehi _4453__231 (.L_HI(net231));
 sg13g2_tiehi _4452__232 (.L_HI(net232));
 sg13g2_tiehi _4451__233 (.L_HI(net233));
 sg13g2_tiehi _4450__234 (.L_HI(net234));
 sg13g2_tiehi _4449__235 (.L_HI(net235));
 sg13g2_tiehi _4448__236 (.L_HI(net236));
 sg13g2_tiehi _4447__237 (.L_HI(net237));
 sg13g2_tiehi _4446__238 (.L_HI(net238));
 sg13g2_tiehi _4445__239 (.L_HI(net239));
 sg13g2_tiehi _4444__240 (.L_HI(net240));
 sg13g2_tiehi _4443__241 (.L_HI(net241));
 sg13g2_tiehi _4442__242 (.L_HI(net242));
 sg13g2_tiehi _4441__243 (.L_HI(net243));
 sg13g2_tiehi _4440__244 (.L_HI(net244));
 sg13g2_tiehi _4439__245 (.L_HI(net245));
 sg13g2_tiehi _4438__246 (.L_HI(net246));
 sg13g2_tiehi _4619__247 (.L_HI(net247));
 sg13g2_tiehi _4437__248 (.L_HI(net248));
 sg13g2_tiehi _4570__249 (.L_HI(net249));
 sg13g2_tiehi _4436__250 (.L_HI(net250));
 sg13g2_tiehi _4643__251 (.L_HI(net251));
 sg13g2_tiehi _4435__252 (.L_HI(net252));
 sg13g2_tiehi _4569__253 (.L_HI(net253));
 sg13g2_tiehi _4434__254 (.L_HI(net254));
 sg13g2_tiehi _4618__255 (.L_HI(net255));
 sg13g2_tiehi _4433__256 (.L_HI(net256));
 sg13g2_tiehi _4568__257 (.L_HI(net257));
 sg13g2_tiehi _4432__258 (.L_HI(net258));
 sg13g2_tiehi _4655__259 (.L_HI(net259));
 sg13g2_tiehi _4431__260 (.L_HI(net260));
 sg13g2_tiehi _4567__261 (.L_HI(net261));
 sg13g2_tiehi _4430__262 (.L_HI(net262));
 sg13g2_tiehi _4429__263 (.L_HI(net263));
 sg13g2_tiehi _4428__264 (.L_HI(net264));
 sg13g2_tiehi _4427__265 (.L_HI(net265));
 sg13g2_tiehi _4426__266 (.L_HI(net266));
 sg13g2_tiehi _4425__267 (.L_HI(net267));
 sg13g2_tiehi _4617__268 (.L_HI(net268));
 sg13g2_tiehi _4424__269 (.L_HI(net269));
 sg13g2_tiehi _4566__270 (.L_HI(net270));
 sg13g2_tiehi _4423__271 (.L_HI(net271));
 sg13g2_tiehi _4642__272 (.L_HI(net272));
 sg13g2_tiehi _4422__273 (.L_HI(net273));
 sg13g2_tiehi _4421__274 (.L_HI(net274));
 sg13g2_tiehi _4420__275 (.L_HI(net275));
 sg13g2_tiehi _4419__276 (.L_HI(net276));
 sg13g2_tiehi _4565__277 (.L_HI(net277));
 sg13g2_tiehi _4418__278 (.L_HI(net278));
 sg13g2_tiehi _4616__279 (.L_HI(net279));
 sg13g2_tiehi _4417__280 (.L_HI(net280));
 sg13g2_tiehi _4564__281 (.L_HI(net281));
 sg13g2_tiehi _4416__282 (.L_HI(net282));
 sg13g2_tiehi _4661__283 (.L_HI(net283));
 sg13g2_tiehi _4415__284 (.L_HI(net284));
 sg13g2_tiehi _4563__285 (.L_HI(net285));
 sg13g2_tiehi _4414__286 (.L_HI(net286));
 sg13g2_tiehi _4615__287 (.L_HI(net287));
 sg13g2_tiehi _4413__288 (.L_HI(net288));
 sg13g2_tiehi _4562__289 (.L_HI(net289));
 sg13g2_tiehi _4412__290 (.L_HI(net290));
 sg13g2_tiehi _4641__291 (.L_HI(net291));
 sg13g2_tiehi _4411__292 (.L_HI(net292));
 sg13g2_tiehi _4561__293 (.L_HI(net293));
 sg13g2_tiehi _4410__294 (.L_HI(net294));
 sg13g2_tiehi _4614__295 (.L_HI(net295));
 sg13g2_tiehi _4409__296 (.L_HI(net296));
 sg13g2_tiehi _4560__297 (.L_HI(net297));
 sg13g2_tiehi _4408__298 (.L_HI(net298));
 sg13g2_tiehi _4654__299 (.L_HI(net299));
 sg13g2_tiehi _4407__300 (.L_HI(net300));
 sg13g2_tiehi _4559__301 (.L_HI(net301));
 sg13g2_tiehi _4406__302 (.L_HI(net302));
 sg13g2_tiehi _4613__303 (.L_HI(net303));
 sg13g2_tiehi _4405__304 (.L_HI(net304));
 sg13g2_tiehi _4558__305 (.L_HI(net305));
 sg13g2_tiehi _4404__306 (.L_HI(net306));
 sg13g2_tiehi _4640__307 (.L_HI(net307));
 sg13g2_tiehi _4403__308 (.L_HI(net308));
 sg13g2_tiehi _4402__309 (.L_HI(net309));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _4965_ (.A(net896),
    .X(uio_oe[0]));
 sg13g2_buf_2 _4966_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_2 _4967_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4968_ (.A(net896),
    .X(uio_oe[3]));
 sg13g2_buf_2 _4969_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4970_ (.A(net896),
    .X(uio_oe[6]));
 sg13g2_buf_1 _4971_ (.A(net896),
    .X(uio_oe[7]));
 sg13g2_buf_2 _4972_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .X(uio_out[0]));
 sg13g2_buf_1 _4973_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .X(uio_out[3]));
 sg13g2_buf_2 _4974_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ),
    .X(uio_out[6]));
 sg13g2_buf_2 _4975_ (.A(\cpu_instance.ctrl_instance.scan_out ),
    .X(uio_out[7]));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_1185_));
 sg13g2_buf_2 fanout680 (.A(_1185_),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(net682));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(_0756_));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(net684));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(_1182_));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(_1179_));
 sg13g2_buf_2 fanout686 (.A(_1179_),
    .X(net686));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net688));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(_0425_));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(net690));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(_0410_));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(net694));
 sg13g2_buf_2 fanout692 (.A(net694),
    .X(net692));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(net694));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(_0397_));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(net696));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(_1176_));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(_1173_));
 sg13g2_buf_2 fanout698 (.A(_1173_),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(_0426_));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(net701));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(_0542_));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(net704));
 sg13g2_buf_2 fanout703 (.A(net704),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_0438_));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(_1168_));
 sg13g2_buf_2 fanout706 (.A(_1168_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_1 fanout708 (.A(_1094_),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_0628_));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(_0628_));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(net713));
 sg13g2_buf_2 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_0512_));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(net716));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(net565));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(net718));
 sg13g2_buf_8 fanout718 (.A(_1793_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_1543_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net723),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_1507_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_0344_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_1899_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_1855_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_1561_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_1561_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_1 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_1552_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(_1534_));
 sg13g2_buf_2 fanout734 (.A(net736),
    .X(net734));
 sg13g2_buf_1 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_1525_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_1516_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(_1267_));
 sg13g2_buf_2 fanout741 (.A(_1191_),
    .X(net741));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(_0659_));
 sg13g2_buf_2 fanout743 (.A(_0659_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_1071_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_0983_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_0667_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_0632_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_1328_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_1314_),
    .X(net751));
 sg13g2_buf_1 fanout752 (.A(_1314_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_1299_),
    .X(net753));
 sg13g2_buf_1 fanout754 (.A(_1299_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_1282_),
    .X(net755));
 sg13g2_buf_4 fanout756 (.X(net756),
    .A(_1052_));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(_1706_));
 sg13g2_buf_1 fanout758 (.A(_1706_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_1654_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_0778_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_1805_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net672),
    .X(net763));
 sg13g2_buf_4 fanout764 (.X(net764),
    .A(_1702_));
 sg13g2_buf_2 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_1673_),
    .X(net766));
 sg13g2_buf_4 fanout767 (.X(net767),
    .A(_1673_));
 sg13g2_buf_2 fanout768 (.A(_1668_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_1652_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_1646_),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(net775));
 sg13g2_buf_2 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(_1276_));
 sg13g2_buf_2 fanout776 (.A(_0892_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_0836_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_0644_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_0639_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_0448_),
    .X(net781));
 sg13g2_buf_4 fanout782 (.X(net782),
    .A(_1694_));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(_1692_));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(_1688_));
 sg13g2_buf_4 fanout785 (.X(net785),
    .A(net786));
 sg13g2_buf_2 fanout786 (.A(_1686_),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(net788));
 sg13g2_buf_2 fanout788 (.A(_1684_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_1667_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_1649_));
 sg13g2_buf_2 fanout791 (.A(_1347_),
    .X(net791));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_1347_));
 sg13g2_buf_2 fanout793 (.A(_0865_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_1727_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_1627_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_1618_));
 sg13g2_buf_2 fanout798 (.A(net799),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_1596_),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(_1592_));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(_1586_));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_1585_));
 sg13g2_buf_2 fanout803 (.A(net622),
    .X(net803));
 sg13g2_buf_1 fanout804 (.A(net622),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_0023_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(net674),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net814),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(net814),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net813),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_1 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(net815));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(net387));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(net667));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(net819));
 sg13g2_buf_2 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(net645),
    .X(net819));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(\cpu_instance.reg_in_sel[1] ));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(net670));
 sg13g2_buf_2 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net824),
    .X(net823));
 sg13g2_buf_1 fanout824 (.A(net830),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(net830),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(net829));
 sg13g2_buf_2 fanout829 (.A(net830),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_1605_),
    .X(net830));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(net832));
 sg13g2_buf_2 fanout832 (.A(_1603_),
    .X(net832));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(net834));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(net835));
 sg13g2_buf_2 fanout835 (.A(_1603_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(net839),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_1 fanout838 (.A(net839),
    .X(net838));
 sg13g2_buf_1 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_1 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(net853));
 sg13g2_buf_2 fanout842 (.A(net853),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net852),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net852),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(net848),
    .X(net846));
 sg13g2_buf_1 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(net852),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net851),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net852),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(ui_in[7]),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net857),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(net856),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(net861),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(net860),
    .X(net858));
 sg13g2_buf_1 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(net871),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net864),
    .X(net862));
 sg13g2_buf_1 fanout863 (.A(net864),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_1 fanout865 (.A(net871),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net871),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(net870),
    .X(net869));
 sg13g2_buf_4 fanout870 (.X(net870),
    .A(net871));
 sg13g2_buf_2 fanout871 (.A(ui_in[7]),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net875),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(net875),
    .X(net873));
 sg13g2_buf_1 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net894),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net894),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net880),
    .X(net877));
 sg13g2_buf_1 fanout878 (.A(net880),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net880),
    .X(net879));
 sg13g2_buf_1 fanout880 (.A(net886),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net886),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(net886),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(net885),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(net886),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(net894),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net893),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net893),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net893),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(net892),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(net893),
    .X(net892));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net894));
 sg13g2_buf_4 fanout894 (.X(net894),
    .A(rst_n));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(net897));
 sg13g2_buf_4 fanout896 (.X(net896),
    .A(net897));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(rst_n));
 sg13g2_buf_2 fanout898 (.A(net903),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net902),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(net902),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net903),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(rst_n),
    .X(net903));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_tiehi _4557__12 (.L_HI(net12));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_3_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_37_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_19_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_20_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[18] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold2 (.A(_1662_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[15] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold4 (.A(_1659_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[17] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold6 (.A(_1661_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[16] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold8 (.A(_1656_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu_instance.registers_instance.registers[1][0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0196_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[14] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.stop_txn ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0035_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[13] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.start_write ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0124_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold17 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold18 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[19] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold19 (.A(_1247_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[3] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[1] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold22 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[2] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[7] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[0] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[0] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[5] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold28 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[2] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[3] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[10] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0152_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[4] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0116_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0154_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0150_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[11] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[1] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0882_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0120_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][10] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0158_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.start_read ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[6] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[9] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0160_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0810_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu_instance.registers_instance.register_bank[9][3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][8] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu_instance.registers_instance.register_bank[9][4] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu_instance.registers_instance.register_bank[15][2] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cpu_instance.registers_instance.register_bank[14][4] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0263_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu_instance.mem_instance.data_qi_mo[7] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0147_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu_instance.registers_instance.registers[0][5] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0178_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu_instance.registers_instance.register_bank[9][0] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cpu_instance.registers_instance.register_bank[13][5] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu_instance.registers_instance.register_bank[10][2] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cpu_instance.registers_instance.register_bank[13][4] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu_instance.registers_instance.register_bank[8][6] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cpu_instance.registers_instance.register_bank[14][1] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu_instance.registers_instance.register_bank[13][7] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu_instance.registers_instance.register_bank[8][1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[2] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0941_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0082_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu_instance.addr_sel ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[1] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0078_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cpu_instance.registers_instance.register_bank[8][3] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu_instance.registers_instance.register_bank[13][2] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu_instance.registers_instance.register_bank[15][0] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu_instance.registers_instance.register_bank[10][4] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cpu_instance.registers_instance.register_bank[11][3] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu_instance.registers_instance.register_bank[10][0] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu_instance.mem_instance.data_qi_mo[6] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][1] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0660_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0094_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0864_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cpu_instance.registers_instance.register_bank[15][6] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu_instance.registers_instance.register_bank[12][4] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cpu_instance.registers_instance.register_bank[9][5] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu_instance.registers_instance.register_bank[11][5] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu_instance.ctrl_instance.jmp_op_addr_sel ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0061_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cpu_instance.registers_instance.register_bank[12][6] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu_instance.registers_instance.register_bank[12][7] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu_instance.registers_instance.register_bank[13][0] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu_instance.registers_instance.register_bank[14][2] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu_instance.registers_instance.register_bank[15][3] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu_instance.registers_instance.register_bank[15][4] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0148_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu_instance.registers_instance.register_bank[10][6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu_instance.registers_instance.registers[0][7] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu_instance.registers_instance.register_bank[8][5] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu_instance.mem_instance.data_qi_mo[2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0142_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][7] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu_instance.mem_instance.data_qi_mo[4] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0144_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu_instance.registers_instance.register_bank[8][7] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu_instance.registers_instance.register_bank[12][3] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cpu_instance.registers_instance.register_bank[10][5] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[1] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0081_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu_instance.registers_instance.register_bank[10][3] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu_instance.mem_instance.data_qi_mo[1] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu_instance.registers_instance.register_bank[13][3] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cpu_instance.registers_instance.register_bank[10][1] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu_instance.registers_instance.registers[0][3] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0176_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu_instance.registers_instance.register_bank[15][7] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cpu_instance.registers_instance.register_bank[9][6] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold130 (.A(\cpu_instance.registers_instance.register_bank[8][4] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cpu_instance.registers_instance.register_bank[8][0] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0733_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu_instance.mem_instance.data_qi_mo[5] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu_instance.addr_reg_op[2] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cpu_instance.registers_instance.register_bank[12][5] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cpu_instance.mem_instance.data_qo_mi[5] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0101_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cpu_instance.registers_instance.register_bank[8][2] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu_instance.registers_instance.register_bank[11][6] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu_instance.mem_instance.data_qi_mo[3] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu_instance.registers_instance.register_bank[11][4] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cpu_instance.registers_instance.register_bank[11][0] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu_instance.registers_instance.register_bank[14][7] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0220_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0221_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu_instance.registers_instance.register_bank[15][1] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu_instance.registers_instance.register_bank[12][1] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu_instance.registers_instance.register_bank[12][0] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu_instance.mem_instance.data_qo_mi[0] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0096_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu_instance.registers_instance.register_bank[15][5] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu_instance.registers_instance.register_bank[11][7] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu_instance.registers_instance.register_bank[14][6] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0323_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cpu_instance.registers_instance.register_bank[14][3] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0244_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu_instance.registers_instance.register_bank[9][2] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu_instance.registers_instance.register_bank[11][1] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu_instance.registers_instance.registers[0][4] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cpu_instance.registers_instance.register_bank[13][6] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0252_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cpu_instance.registers_instance.register_bank[10][7] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0258_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0247_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0250_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cpu_instance.mem_instance.data_qo_mi[4] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cpu_instance.registers_instance.register_bank[14][5] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cpu_instance.registers_instance.register_bank[13][1] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0268_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cpu_instance.mem_instance.bus_data_out[7] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold181 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0222_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold183 (.A(\cpu_instance.registers_instance.register_bank[11][2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold184 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0262_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cpu_instance.registers_instance.register_bank[9][7] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold187 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0230_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cpu_instance.registers_instance.registers[0][6] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cpu_instance.ctrl_instance.scan_in ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0224_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold194 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0241_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0227_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0259_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold202 (.A(\cpu_instance.mem_instance.data_qo_mi[2] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold203 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0266_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold205 (.A(\cpu_instance.registers_instance.register_bank[9][1] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0242_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold208 (.A(\cpu_instance.mem_instance.data_qo_mi[1] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold209 (.A(\cpu_instance.mem_instance.data_qo_mi[7] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0103_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold211 (.A(\cpu_instance.registers_instance.registers[0][0] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0173_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold213 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold214 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0267_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold216 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0238_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold218 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0235_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cpu_instance.registers_instance.registers[1][6] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0186_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold223 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold224 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0226_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold226 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold228 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold230 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold231 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold232 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold233 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold234 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold235 (.A(_1242_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold236 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0248_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold239 (.A(\cpu_instance.mem_instance.data_qo_mi[6] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold240 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold241 (.A(\cpu_instance.registers_instance.register_bank[14][0] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0317_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold243 (.A(\cpu_instance.registers_instance.registers[0][2] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold244 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0080_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold246 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0237_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold248 (.A(\cpu_instance.registers_instance.registers[2][6] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0195_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cpu_instance.registers_instance.registers[1][7] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold251 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold252 (.A(\cpu_instance.registers_instance.register_bank[12][2] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold253 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold254 (.A(\cpu_instance.mem_instance.bus_data_out[6] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold255 (.A(\cpu_instance.mem_instance.bus_data_out[1] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0525_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold257 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold258 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold259 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0205_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold261 (.A(\cpu_instance.mem_instance.bus_data_out[4] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0131_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold263 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0696_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold265 (.A(\cpu_instance.registers_instance.registers[2][5] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cpu_instance.mem_instance.bus_data_out[5] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold267 (.A(\cpu_instance.mem_instance.data_req ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0207_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold270 (.A(\cpu_instance.registers_instance.registers[2][1] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0189_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cpu_instance.mem_ctrl_op[1] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0585_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold274 (.A(uo_out[3]),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0200_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold276 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0211_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold278 (.A(\cpu_instance.registers_instance.registers[1][3] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0183_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold280 (.A(\cpu_instance.ctrl_instance.state[0] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0589_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold282 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold283 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0217_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold285 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold286 (.A(\cpu_instance.mux_instance.sel[1] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0493_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold288 (.A(\cpu_instance.mem_instance.bus_data_out[2] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold289 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold290 (.A(\cpu_instance.mem_instance.data_qo_mi[3] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold291 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold292 (.A(\cpu_instance.registers_instance.registers[2][4] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold293 (.A(\cpu_instance.registers_instance.registers[1][1] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold294 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold295 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold296 (.A(\cpu_instance.registers_instance.registers[1][5] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0185_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold298 (.A(\cpu_instance.reg_2_out_sel[1] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold299 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold300 (.A(uo_out[2]),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold301 (.A(\cpu_instance.mem_instance.bus_data_out[3] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold302 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0214_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold304 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold305 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold306 (.A(\cpu_instance.ctrl_instance.flag_carry ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0572_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold308 (.A(\cpu_instance.registers_instance.registers[2][3] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0191_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold310 (.A(uo_out[6]),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0203_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold312 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold313 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.is_writing ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0083_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold315 (.A(\cpu_instance.registers_instance.registers[0][1] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold316 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0212_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold318 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0093_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold320 (.A(\cpu_instance.registers_instance.registers[2][2] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold321 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold322 (.A(uo_out[7]),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0204_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold324 (.A(uo_out[5]),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold325 (.A(\cpu_instance.ctrl_instance.flag_zero ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold326 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold327 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold328 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold329 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0095_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold331 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold332 (.A(\cpu_instance.registers_instance.registers[1][4] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold333 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold334 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0208_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold336 (.A(\cpu_instance.reg_1_out_sel[0] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold337 (.A(\cpu_instance.registers_instance.registers[1][2] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold338 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold339 (.A(uo_out[4]),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold340 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold341 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold342 (.A(\cpu_instance.ctrl_instance.mem_op_done ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0126_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold344 (.A(uo_out[1]),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0197_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold346 (.A(\cpu_instance.ctrl_instance.state[2] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0038_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold348 (.A(\cpu_instance.addr_reg_op[1] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold349 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold350 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold351 (.A(\cpu_instance.ctrl_instance.state[1] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0037_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold353 (.A(\cpu_instance.mem_ctrl_op[0] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold354 (.A(\cpu_instance.alu_instance.op[0] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold355 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold356 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold357 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold358 (.A(\cpu_instance.reg_1_out_sel[1] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold359 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold360 (.A(\cpu_instance.mem_instance.bus_data_out[0] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold361 (.A(\cpu_instance.reg_in_sel[0] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold362 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.stop_txn_reg ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold363 (.A(_1805_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0089_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold365 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold366 (.A(\cpu_instance.ctrl_instance.use_register_bank_in ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0551_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold368 (.A(\cpu_instance.alu_instance.op[1] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold369 (.A(\cpu_instance.alu_instance.op[2] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold370 (.A(\cpu_instance.addr_reg_op[0] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold371 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.stop_txn ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold372 (.A(\cpu_instance.alu_instance.op[3] ),
    .X(net906));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_4 FILLER_0_287 ();
 sg13g2_fill_1 FILLER_0_291 ();
 sg13g2_fill_2 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_4 FILLER_0_309 ();
 sg13g2_fill_2 FILLER_0_313 ();
 sg13g2_fill_1 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_fill_2 FILLER_1_280 ();
 sg13g2_fill_2 FILLER_1_328 ();
 sg13g2_fill_1 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_4 FILLER_2_196 ();
 sg13g2_fill_1 FILLER_2_200 ();
 sg13g2_fill_1 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_251 ();
 sg13g2_fill_1 FILLER_2_278 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_fill_2 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_128 ();
 sg13g2_decap_8 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_decap_8 FILLER_3_176 ();
 sg13g2_decap_8 FILLER_3_183 ();
 sg13g2_decap_8 FILLER_3_190 ();
 sg13g2_decap_4 FILLER_3_197 ();
 sg13g2_fill_1 FILLER_3_201 ();
 sg13g2_decap_4 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_250 ();
 sg13g2_fill_2 FILLER_3_296 ();
 sg13g2_fill_1 FILLER_3_312 ();
 sg13g2_fill_2 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_fill_1 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_68 ();
 sg13g2_decap_8 FILLER_4_75 ();
 sg13g2_decap_8 FILLER_4_82 ();
 sg13g2_decap_8 FILLER_4_89 ();
 sg13g2_decap_8 FILLER_4_96 ();
 sg13g2_decap_4 FILLER_4_103 ();
 sg13g2_decap_8 FILLER_4_167 ();
 sg13g2_decap_8 FILLER_4_174 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_1 FILLER_4_191 ();
 sg13g2_decap_8 FILLER_4_197 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_4 FILLER_4_211 ();
 sg13g2_decap_4 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_239 ();
 sg13g2_fill_2 FILLER_4_245 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_320 ();
 sg13g2_fill_1 FILLER_4_322 ();
 sg13g2_fill_1 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_4 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_83 ();
 sg13g2_decap_4 FILLER_5_90 ();
 sg13g2_fill_2 FILLER_5_94 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_4 FILLER_5_147 ();
 sg13g2_fill_1 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_decap_8 FILLER_5_163 ();
 sg13g2_fill_2 FILLER_5_170 ();
 sg13g2_fill_1 FILLER_5_172 ();
 sg13g2_fill_2 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_decap_4 FILLER_5_239 ();
 sg13g2_fill_1 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_4 FILLER_6_113 ();
 sg13g2_fill_2 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_128 ();
 sg13g2_decap_4 FILLER_6_138 ();
 sg13g2_fill_1 FILLER_6_155 ();
 sg13g2_decap_4 FILLER_6_182 ();
 sg13g2_fill_2 FILLER_6_195 ();
 sg13g2_fill_1 FILLER_6_216 ();
 sg13g2_fill_2 FILLER_6_292 ();
 sg13g2_fill_1 FILLER_6_294 ();
 sg13g2_fill_2 FILLER_6_354 ();
 sg13g2_fill_1 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_44 ();
 sg13g2_fill_2 FILLER_7_64 ();
 sg13g2_fill_2 FILLER_7_92 ();
 sg13g2_decap_4 FILLER_7_112 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_fill_2 FILLER_7_270 ();
 sg13g2_fill_1 FILLER_7_272 ();
 sg13g2_decap_4 FILLER_7_316 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_fill_1 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_4 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_25 ();
 sg13g2_fill_1 FILLER_8_52 ();
 sg13g2_fill_1 FILLER_8_57 ();
 sg13g2_fill_2 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_65 ();
 sg13g2_decap_4 FILLER_8_71 ();
 sg13g2_fill_2 FILLER_8_75 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_95 ();
 sg13g2_fill_1 FILLER_8_115 ();
 sg13g2_fill_2 FILLER_8_130 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_fill_2 FILLER_8_181 ();
 sg13g2_fill_1 FILLER_8_183 ();
 sg13g2_fill_2 FILLER_8_244 ();
 sg13g2_fill_1 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_262 ();
 sg13g2_fill_2 FILLER_8_269 ();
 sg13g2_decap_4 FILLER_8_277 ();
 sg13g2_fill_1 FILLER_8_281 ();
 sg13g2_fill_1 FILLER_8_291 ();
 sg13g2_decap_4 FILLER_8_315 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_351 ();
 sg13g2_fill_1 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_36 ();
 sg13g2_fill_1 FILLER_9_41 ();
 sg13g2_fill_2 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_97 ();
 sg13g2_fill_1 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_131 ();
 sg13g2_decap_8 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_195 ();
 sg13g2_fill_2 FILLER_9_206 ();
 sg13g2_fill_1 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_279 ();
 sg13g2_fill_2 FILLER_9_286 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_fill_1 FILLER_9_335 ();
 sg13g2_fill_2 FILLER_9_366 ();
 sg13g2_fill_1 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_65 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_164 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_decap_8 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_195 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_decap_4 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_242 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_254 ();
 sg13g2_fill_2 FILLER_10_260 ();
 sg13g2_fill_1 FILLER_10_262 ();
 sg13g2_decap_4 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_313 ();
 sg13g2_fill_1 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_fill_2 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_47 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_fill_2 FILLER_11_134 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_fill_2 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_fill_2 FILLER_11_219 ();
 sg13g2_fill_1 FILLER_11_221 ();
 sg13g2_decap_4 FILLER_11_228 ();
 sg13g2_fill_1 FILLER_11_232 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_4 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_fill_2 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_fill_2 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_1 FILLER_11_330 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_fill_2 FILLER_11_353 ();
 sg13g2_fill_1 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_4 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_57 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_fill_1 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_fill_2 FILLER_12_142 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_fill_2 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_decap_4 FILLER_12_260 ();
 sg13g2_fill_1 FILLER_12_278 ();
 sg13g2_decap_4 FILLER_12_338 ();
 sg13g2_fill_2 FILLER_12_342 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_33 ();
 sg13g2_fill_1 FILLER_13_69 ();
 sg13g2_decap_4 FILLER_13_108 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_2 FILLER_13_132 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_178 ();
 sg13g2_fill_2 FILLER_13_188 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_277 ();
 sg13g2_fill_2 FILLER_13_283 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_339 ();
 sg13g2_fill_1 FILLER_13_341 ();
 sg13g2_fill_2 FILLER_13_373 ();
 sg13g2_fill_1 FILLER_13_375 ();
 sg13g2_fill_2 FILLER_13_385 ();
 sg13g2_fill_1 FILLER_13_387 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_fill_2 FILLER_14_60 ();
 sg13g2_fill_2 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_106 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_114 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_140 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_164 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_2 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_205 ();
 sg13g2_decap_4 FILLER_14_211 ();
 sg13g2_decap_8 FILLER_14_281 ();
 sg13g2_fill_2 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_290 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_fill_2 FILLER_14_316 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_fill_2 FILLER_14_371 ();
 sg13g2_decap_4 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_fill_2 FILLER_15_26 ();
 sg13g2_fill_2 FILLER_15_37 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_fill_1 FILLER_15_48 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_decap_8 FILLER_15_64 ();
 sg13g2_fill_2 FILLER_15_71 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_2 FILLER_15_87 ();
 sg13g2_fill_2 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_fill_2 FILLER_15_233 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_1 FILLER_15_316 ();
 sg13g2_fill_1 FILLER_15_322 ();
 sg13g2_decap_4 FILLER_15_333 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_24 ();
 sg13g2_decap_8 FILLER_16_50 ();
 sg13g2_decap_8 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_69 ();
 sg13g2_fill_2 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_113 ();
 sg13g2_decap_4 FILLER_16_128 ();
 sg13g2_fill_2 FILLER_16_132 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_decap_4 FILLER_16_195 ();
 sg13g2_fill_2 FILLER_16_199 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_217 ();
 sg13g2_fill_2 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_245 ();
 sg13g2_fill_2 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_315 ();
 sg13g2_fill_1 FILLER_16_357 ();
 sg13g2_fill_2 FILLER_16_363 ();
 sg13g2_fill_2 FILLER_16_380 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_20 ();
 sg13g2_fill_2 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_fill_1 FILLER_17_104 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_decap_8 FILLER_17_227 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_4 FILLER_17_241 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_decap_4 FILLER_17_336 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_26 ();
 sg13g2_decap_4 FILLER_18_37 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_99 ();
 sg13g2_fill_1 FILLER_18_101 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_decap_8 FILLER_18_128 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_4 FILLER_18_157 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_fill_2 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_decap_4 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_246 ();
 sg13g2_decap_4 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_4 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_348 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_26 ();
 sg13g2_decap_8 FILLER_19_45 ();
 sg13g2_decap_8 FILLER_19_57 ();
 sg13g2_decap_8 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_71 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_decap_4 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_decap_4 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_186 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_264 ();
 sg13g2_decap_4 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_375 ();
 sg13g2_fill_1 FILLER_19_381 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_19 ();
 sg13g2_fill_1 FILLER_20_26 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_43 ();
 sg13g2_fill_2 FILLER_20_54 ();
 sg13g2_decap_8 FILLER_20_61 ();
 sg13g2_decap_8 FILLER_20_68 ();
 sg13g2_decap_8 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_82 ();
 sg13g2_decap_8 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_decap_4 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_130 ();
 sg13g2_fill_2 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_213 ();
 sg13g2_decap_4 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_311 ();
 sg13g2_decap_4 FILLER_20_319 ();
 sg13g2_fill_1 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_fill_2 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_15 ();
 sg13g2_fill_1 FILLER_21_22 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_69 ();
 sg13g2_decap_8 FILLER_21_79 ();
 sg13g2_decap_8 FILLER_21_86 ();
 sg13g2_fill_1 FILLER_21_93 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_4 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_154 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_decap_4 FILLER_21_273 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_1 FILLER_22_40 ();
 sg13g2_decap_4 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_2 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_decap_4 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_121 ();
 sg13g2_fill_2 FILLER_22_145 ();
 sg13g2_fill_1 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_170 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_decap_4 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_decap_4 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_decap_4 FILLER_22_390 ();
 sg13g2_fill_2 FILLER_22_394 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_fill_2 FILLER_23_52 ();
 sg13g2_fill_2 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_102 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_132 ();
 sg13g2_fill_2 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_decap_4 FILLER_23_308 ();
 sg13g2_decap_4 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_32 ();
 sg13g2_fill_2 FILLER_24_36 ();
 sg13g2_decap_8 FILLER_24_52 ();
 sg13g2_decap_4 FILLER_24_59 ();
 sg13g2_decap_4 FILLER_24_68 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_150 ();
 sg13g2_decap_4 FILLER_24_157 ();
 sg13g2_decap_8 FILLER_24_169 ();
 sg13g2_decap_8 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_decap_4 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_decap_4 FILLER_24_356 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_18 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_76 ();
 sg13g2_decap_8 FILLER_25_87 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_decap_4 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_decap_4 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_262 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_313 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_fill_2 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_16 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_2 FILLER_26_40 ();
 sg13g2_fill_2 FILLER_26_57 ();
 sg13g2_fill_2 FILLER_26_65 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_90 ();
 sg13g2_fill_2 FILLER_26_97 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_decap_4 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_decap_4 FILLER_26_149 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_decap_4 FILLER_26_280 ();
 sg13g2_decap_4 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_fill_1 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_11 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_114 ();
 sg13g2_decap_4 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_decap_4 FILLER_27_292 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_4 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_decap_4 FILLER_28_101 ();
 sg13g2_decap_4 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_120 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_decap_4 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_199 ();
 sg13g2_decap_8 FILLER_28_243 ();
 sg13g2_decap_4 FILLER_28_250 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_decap_4 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_decap_8 FILLER_28_337 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_fill_1 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_395 ();
 sg13g2_fill_1 FILLER_28_397 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_40 ();
 sg13g2_decap_4 FILLER_29_50 ();
 sg13g2_fill_1 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_4 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_223 ();
 sg13g2_decap_4 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_fill_2 FILLER_29_365 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_26 ();
 sg13g2_decap_8 FILLER_30_34 ();
 sg13g2_decap_8 FILLER_30_41 ();
 sg13g2_decap_8 FILLER_30_48 ();
 sg13g2_decap_8 FILLER_30_55 ();
 sg13g2_decap_4 FILLER_30_62 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_76 ();
 sg13g2_decap_8 FILLER_30_83 ();
 sg13g2_decap_4 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_94 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_decap_4 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_decap_8 FILLER_31_47 ();
 sg13g2_decap_8 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_68 ();
 sg13g2_decap_8 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_93 ();
 sg13g2_decap_8 FILLER_31_97 ();
 sg13g2_decap_8 FILLER_31_104 ();
 sg13g2_decap_8 FILLER_31_111 ();
 sg13g2_decap_4 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_134 ();
 sg13g2_decap_8 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_155 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_4 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_273 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_1 FILLER_32_29 ();
 sg13g2_fill_1 FILLER_32_43 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_113 ();
 sg13g2_fill_2 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_145 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_261 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_338 ();
 sg13g2_decap_8 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_356 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_fill_1 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_38 ();
 sg13g2_decap_4 FILLER_33_45 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_93 ();
 sg13g2_decap_4 FILLER_33_100 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_decap_4 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_decap_4 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_decap_4 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_2 FILLER_34_72 ();
 sg13g2_fill_2 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_92 ();
 sg13g2_fill_1 FILLER_34_94 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_156 ();
 sg13g2_decap_4 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_201 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_332 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_fill_1 FILLER_34_369 ();
 sg13g2_decap_4 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_27 ();
 sg13g2_fill_1 FILLER_35_46 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_decap_8 FILLER_35_103 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_134 ();
 sg13g2_decap_4 FILLER_35_141 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_227 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_287 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_36_26 ();
 sg13g2_fill_1 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_59 ();
 sg13g2_fill_2 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_89 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_decap_8 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_decap_4 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_4 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_363 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_24 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_110 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_222 ();
 sg13g2_decap_4 FILLER_37_229 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_decap_4 FILLER_37_263 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_293 ();
 sg13g2_fill_2 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_4 FILLER_37_360 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_371 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_25 ();
 sg13g2_decap_4 FILLER_38_31 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_40 ();
 sg13g2_fill_1 FILLER_38_67 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_131 ();
 sg13g2_decap_4 FILLER_38_146 ();
 sg13g2_decap_4 FILLER_38_171 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_184 ();
 sg13g2_decap_4 FILLER_38_191 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_258 ();
 sg13g2_decap_4 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_decap_4 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_fill_2 FILLER_39_32 ();
 sg13g2_decap_8 FILLER_39_40 ();
 sg13g2_decap_8 FILLER_39_47 ();
 sg13g2_fill_1 FILLER_39_54 ();
 sg13g2_decap_8 FILLER_39_128 ();
 sg13g2_decap_4 FILLER_39_135 ();
 sg13g2_fill_2 FILLER_39_139 ();
 sg13g2_decap_8 FILLER_39_151 ();
 sg13g2_decap_8 FILLER_39_158 ();
 sg13g2_fill_2 FILLER_39_165 ();
 sg13g2_decap_8 FILLER_39_177 ();
 sg13g2_decap_8 FILLER_39_184 ();
 sg13g2_decap_8 FILLER_39_191 ();
 sg13g2_decap_8 FILLER_39_198 ();
 sg13g2_decap_8 FILLER_39_205 ();
 sg13g2_decap_4 FILLER_39_212 ();
 sg13g2_fill_1 FILLER_39_220 ();
 sg13g2_fill_2 FILLER_39_280 ();
 sg13g2_fill_2 FILLER_39_296 ();
 sg13g2_decap_8 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_314 ();
 sg13g2_decap_8 FILLER_39_321 ();
 sg13g2_decap_4 FILLER_39_333 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_364 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_55 ();
 sg13g2_decap_8 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_69 ();
 sg13g2_decap_8 FILLER_40_75 ();
 sg13g2_decap_8 FILLER_40_82 ();
 sg13g2_fill_2 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_decap_4 FILLER_40_109 ();
 sg13g2_fill_2 FILLER_40_113 ();
 sg13g2_decap_8 FILLER_40_123 ();
 sg13g2_decap_8 FILLER_40_130 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_decap_4 FILLER_40_144 ();
 sg13g2_fill_2 FILLER_40_148 ();
 sg13g2_fill_2 FILLER_40_176 ();
 sg13g2_decap_8 FILLER_40_181 ();
 sg13g2_fill_1 FILLER_40_196 ();
 sg13g2_decap_4 FILLER_40_241 ();
 sg13g2_decap_4 FILLER_40_276 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_fill_2 FILLER_40_319 ();
 sg13g2_fill_1 FILLER_40_327 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_fill_1 FILLER_40_387 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_4 ();
 sg13g2_fill_2 FILLER_41_27 ();
 sg13g2_fill_2 FILLER_41_64 ();
 sg13g2_fill_1 FILLER_41_80 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_fill_1 FILLER_41_89 ();
 sg13g2_decap_4 FILLER_41_99 ();
 sg13g2_fill_1 FILLER_41_103 ();
 sg13g2_fill_1 FILLER_41_134 ();
 sg13g2_fill_2 FILLER_41_140 ();
 sg13g2_fill_2 FILLER_41_153 ();
 sg13g2_fill_1 FILLER_41_155 ();
 sg13g2_fill_1 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_176 ();
 sg13g2_decap_4 FILLER_41_187 ();
 sg13g2_fill_2 FILLER_41_191 ();
 sg13g2_fill_2 FILLER_41_262 ();
 sg13g2_decap_8 FILLER_41_298 ();
 sg13g2_decap_4 FILLER_41_305 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_decap_4 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_360 ();
 sg13g2_decap_8 FILLER_41_367 ();
 sg13g2_decap_8 FILLER_42_97 ();
 sg13g2_fill_1 FILLER_42_104 ();
 sg13g2_fill_2 FILLER_42_163 ();
 sg13g2_fill_1 FILLER_42_165 ();
 sg13g2_fill_2 FILLER_42_176 ();
 sg13g2_fill_1 FILLER_42_178 ();
 sg13g2_fill_1 FILLER_42_188 ();
 sg13g2_fill_2 FILLER_42_197 ();
 sg13g2_fill_1 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_246 ();
 sg13g2_decap_8 FILLER_42_253 ();
 sg13g2_fill_2 FILLER_42_260 ();
 sg13g2_decap_4 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_270 ();
 sg13g2_fill_1 FILLER_42_321 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_fill_2 FILLER_42_362 ();
 sg13g2_decap_4 FILLER_42_374 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_15 ();
 sg13g2_fill_1 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_86 ();
 sg13g2_fill_1 FILLER_43_93 ();
 sg13g2_decap_8 FILLER_43_102 ();
 sg13g2_decap_8 FILLER_43_109 ();
 sg13g2_fill_2 FILLER_43_120 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_fill_2 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_157 ();
 sg13g2_fill_2 FILLER_43_199 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_decap_4 FILLER_43_217 ();
 sg13g2_fill_2 FILLER_43_221 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_239 ();
 sg13g2_fill_1 FILLER_43_272 ();
 sg13g2_fill_2 FILLER_43_297 ();
 sg13g2_fill_1 FILLER_43_299 ();
 sg13g2_decap_8 FILLER_43_318 ();
 sg13g2_fill_2 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_341 ();
 sg13g2_fill_2 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_80 ();
 sg13g2_fill_1 FILLER_44_82 ();
 sg13g2_decap_8 FILLER_44_115 ();
 sg13g2_decap_4 FILLER_44_122 ();
 sg13g2_fill_2 FILLER_44_135 ();
 sg13g2_fill_1 FILLER_44_157 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_fill_1 FILLER_44_174 ();
 sg13g2_decap_4 FILLER_44_195 ();
 sg13g2_fill_2 FILLER_44_199 ();
 sg13g2_decap_8 FILLER_44_209 ();
 sg13g2_fill_2 FILLER_44_216 ();
 sg13g2_decap_4 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_267 ();
 sg13g2_decap_8 FILLER_44_297 ();
 sg13g2_decap_4 FILLER_44_304 ();
 sg13g2_fill_2 FILLER_44_321 ();
 sg13g2_fill_1 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_381 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_11 ();
 sg13g2_decap_4 FILLER_45_19 ();
 sg13g2_fill_1 FILLER_45_23 ();
 sg13g2_decap_4 FILLER_45_62 ();
 sg13g2_decap_8 FILLER_45_71 ();
 sg13g2_decap_8 FILLER_45_78 ();
 sg13g2_decap_8 FILLER_45_85 ();
 sg13g2_fill_2 FILLER_45_92 ();
 sg13g2_fill_2 FILLER_45_98 ();
 sg13g2_fill_1 FILLER_45_100 ();
 sg13g2_decap_8 FILLER_45_149 ();
 sg13g2_decap_8 FILLER_45_156 ();
 sg13g2_decap_8 FILLER_45_163 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_decap_8 FILLER_45_177 ();
 sg13g2_decap_8 FILLER_45_184 ();
 sg13g2_decap_4 FILLER_45_191 ();
 sg13g2_fill_1 FILLER_45_195 ();
 sg13g2_decap_4 FILLER_45_204 ();
 sg13g2_fill_1 FILLER_45_208 ();
 sg13g2_fill_2 FILLER_45_333 ();
 sg13g2_decap_8 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_346 ();
 sg13g2_fill_1 FILLER_45_348 ();
 sg13g2_fill_1 FILLER_45_363 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_15 ();
 sg13g2_decap_4 FILLER_46_22 ();
 sg13g2_fill_2 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_52 ();
 sg13g2_decap_8 FILLER_46_59 ();
 sg13g2_decap_8 FILLER_46_66 ();
 sg13g2_decap_4 FILLER_46_77 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_decap_8 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_144 ();
 sg13g2_decap_8 FILLER_46_151 ();
 sg13g2_decap_4 FILLER_46_158 ();
 sg13g2_fill_2 FILLER_46_162 ();
 sg13g2_fill_2 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_181 ();
 sg13g2_decap_4 FILLER_46_188 ();
 sg13g2_fill_2 FILLER_46_205 ();
 sg13g2_decap_4 FILLER_46_248 ();
 sg13g2_fill_2 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_258 ();
 sg13g2_decap_4 FILLER_46_265 ();
 sg13g2_fill_2 FILLER_46_269 ();
 sg13g2_fill_2 FILLER_46_297 ();
 sg13g2_fill_1 FILLER_46_299 ();
 sg13g2_fill_2 FILLER_46_316 ();
 sg13g2_fill_1 FILLER_46_318 ();
 sg13g2_decap_8 FILLER_46_339 ();
 sg13g2_decap_4 FILLER_46_346 ();
 sg13g2_fill_1 FILLER_46_350 ();
 sg13g2_fill_2 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_393 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_fill_1 FILLER_47_26 ();
 sg13g2_decap_8 FILLER_47_41 ();
 sg13g2_decap_8 FILLER_47_48 ();
 sg13g2_decap_8 FILLER_47_55 ();
 sg13g2_fill_1 FILLER_47_62 ();
 sg13g2_fill_1 FILLER_47_110 ();
 sg13g2_decap_4 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_119 ();
 sg13g2_fill_1 FILLER_47_125 ();
 sg13g2_decap_8 FILLER_47_136 ();
 sg13g2_fill_1 FILLER_47_143 ();
 sg13g2_fill_2 FILLER_47_148 ();
 sg13g2_fill_1 FILLER_47_150 ();
 sg13g2_fill_2 FILLER_47_167 ();
 sg13g2_decap_8 FILLER_47_205 ();
 sg13g2_fill_1 FILLER_47_221 ();
 sg13g2_fill_1 FILLER_47_227 ();
 sg13g2_fill_1 FILLER_47_242 ();
 sg13g2_decap_8 FILLER_47_269 ();
 sg13g2_decap_4 FILLER_47_276 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_286 ();
 sg13g2_decap_8 FILLER_47_293 ();
 sg13g2_decap_4 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_327 ();
 sg13g2_decap_8 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_356 ();
 sg13g2_fill_1 FILLER_47_363 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_77 ();
 sg13g2_fill_1 FILLER_48_79 ();
 sg13g2_fill_2 FILLER_48_106 ();
 sg13g2_decap_8 FILLER_48_117 ();
 sg13g2_decap_4 FILLER_48_134 ();
 sg13g2_fill_2 FILLER_48_143 ();
 sg13g2_fill_1 FILLER_48_150 ();
 sg13g2_fill_2 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_decap_4 FILLER_48_181 ();
 sg13g2_decap_8 FILLER_48_220 ();
 sg13g2_fill_2 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_fill_2 FILLER_48_294 ();
 sg13g2_fill_1 FILLER_48_296 ();
 sg13g2_decap_8 FILLER_48_304 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_48_316 ();
 sg13g2_decap_4 FILLER_48_323 ();
 sg13g2_fill_1 FILLER_48_327 ();
 sg13g2_decap_8 FILLER_48_332 ();
 sg13g2_decap_8 FILLER_48_349 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_48_370 ();
 sg13g2_decap_8 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_48_384 ();
 sg13g2_fill_1 FILLER_48_391 ();
 sg13g2_decap_8 FILLER_48_396 ();
 sg13g2_decap_4 FILLER_48_403 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_fill_2 FILLER_49_26 ();
 sg13g2_fill_1 FILLER_49_55 ();
 sg13g2_fill_1 FILLER_49_78 ();
 sg13g2_fill_1 FILLER_49_90 ();
 sg13g2_decap_8 FILLER_49_164 ();
 sg13g2_decap_8 FILLER_49_171 ();
 sg13g2_decap_8 FILLER_49_178 ();
 sg13g2_decap_8 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_192 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_216 ();
 sg13g2_fill_1 FILLER_49_218 ();
 sg13g2_decap_4 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_299 ();
 sg13g2_fill_2 FILLER_49_320 ();
 sg13g2_decap_4 FILLER_49_361 ();
 sg13g2_fill_2 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_fill_2 FILLER_49_379 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_fill_1 FILLER_50_32 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_decap_4 FILLER_50_67 ();
 sg13g2_fill_2 FILLER_50_71 ();
 sg13g2_fill_2 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_79 ();
 sg13g2_decap_8 FILLER_50_88 ();
 sg13g2_decap_8 FILLER_50_95 ();
 sg13g2_decap_4 FILLER_50_102 ();
 sg13g2_fill_2 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_134 ();
 sg13g2_decap_8 FILLER_50_165 ();
 sg13g2_fill_1 FILLER_50_172 ();
 sg13g2_decap_4 FILLER_50_177 ();
 sg13g2_fill_1 FILLER_50_181 ();
 sg13g2_decap_8 FILLER_50_191 ();
 sg13g2_decap_8 FILLER_50_198 ();
 sg13g2_decap_8 FILLER_50_205 ();
 sg13g2_fill_2 FILLER_50_212 ();
 sg13g2_decap_4 FILLER_50_218 ();
 sg13g2_fill_2 FILLER_50_222 ();
 sg13g2_fill_1 FILLER_50_229 ();
 sg13g2_decap_4 FILLER_50_238 ();
 sg13g2_fill_1 FILLER_50_242 ();
 sg13g2_decap_4 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_252 ();
 sg13g2_fill_2 FILLER_50_262 ();
 sg13g2_fill_1 FILLER_50_264 ();
 sg13g2_decap_8 FILLER_50_325 ();
 sg13g2_decap_4 FILLER_50_332 ();
 sg13g2_fill_1 FILLER_50_341 ();
 sg13g2_fill_2 FILLER_50_347 ();
 sg13g2_fill_2 FILLER_50_380 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_52 ();
 sg13g2_decap_8 FILLER_51_60 ();
 sg13g2_decap_8 FILLER_51_72 ();
 sg13g2_decap_8 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_86 ();
 sg13g2_decap_8 FILLER_51_96 ();
 sg13g2_decap_4 FILLER_51_103 ();
 sg13g2_decap_4 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_115 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_1 FILLER_51_184 ();
 sg13g2_fill_1 FILLER_51_230 ();
 sg13g2_decap_8 FILLER_51_244 ();
 sg13g2_decap_8 FILLER_51_251 ();
 sg13g2_decap_4 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_fill_1 FILLER_51_291 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_fill_2 FILLER_51_335 ();
 sg13g2_fill_1 FILLER_51_374 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_11 ();
 sg13g2_decap_4 FILLER_52_17 ();
 sg13g2_fill_1 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_36 ();
 sg13g2_decap_4 FILLER_52_55 ();
 sg13g2_fill_2 FILLER_52_59 ();
 sg13g2_decap_8 FILLER_52_69 ();
 sg13g2_decap_4 FILLER_52_76 ();
 sg13g2_fill_2 FILLER_52_80 ();
 sg13g2_fill_1 FILLER_52_95 ();
 sg13g2_fill_1 FILLER_52_127 ();
 sg13g2_fill_2 FILLER_52_133 ();
 sg13g2_fill_2 FILLER_52_149 ();
 sg13g2_fill_2 FILLER_52_156 ();
 sg13g2_fill_2 FILLER_52_162 ();
 sg13g2_fill_2 FILLER_52_182 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_decap_4 FILLER_52_217 ();
 sg13g2_fill_1 FILLER_52_221 ();
 sg13g2_decap_8 FILLER_52_230 ();
 sg13g2_decap_8 FILLER_52_257 ();
 sg13g2_decap_8 FILLER_52_264 ();
 sg13g2_decap_8 FILLER_52_271 ();
 sg13g2_fill_2 FILLER_52_278 ();
 sg13g2_fill_2 FILLER_52_306 ();
 sg13g2_fill_1 FILLER_52_327 ();
 sg13g2_decap_8 FILLER_52_346 ();
 sg13g2_fill_1 FILLER_52_353 ();
 sg13g2_fill_1 FILLER_52_368 ();
 sg13g2_fill_2 FILLER_52_380 ();
 sg13g2_decap_8 FILLER_52_397 ();
 sg13g2_decap_4 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_21 ();
 sg13g2_fill_1 FILLER_53_23 ();
 sg13g2_decap_4 FILLER_53_29 ();
 sg13g2_fill_2 FILLER_53_52 ();
 sg13g2_fill_1 FILLER_53_74 ();
 sg13g2_fill_1 FILLER_53_101 ();
 sg13g2_fill_2 FILLER_53_141 ();
 sg13g2_fill_1 FILLER_53_143 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_fill_1 FILLER_53_175 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_211 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_231 ();
 sg13g2_decap_8 FILLER_53_275 ();
 sg13g2_decap_4 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_286 ();
 sg13g2_fill_2 FILLER_53_292 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_decap_8 FILLER_53_332 ();
 sg13g2_decap_4 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_343 ();
 sg13g2_fill_1 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_384 ();
 sg13g2_fill_1 FILLER_53_390 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_fill_1 FILLER_54_26 ();
 sg13g2_fill_2 FILLER_54_100 ();
 sg13g2_fill_1 FILLER_54_107 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_152 ();
 sg13g2_fill_2 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_181 ();
 sg13g2_fill_2 FILLER_54_209 ();
 sg13g2_fill_2 FILLER_54_233 ();
 sg13g2_fill_1 FILLER_54_235 ();
 sg13g2_fill_2 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_253 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_294 ();
 sg13g2_decap_4 FILLER_54_301 ();
 sg13g2_fill_2 FILLER_54_305 ();
 sg13g2_decap_8 FILLER_54_312 ();
 sg13g2_decap_8 FILLER_54_319 ();
 sg13g2_decap_4 FILLER_54_333 ();
 sg13g2_decap_4 FILLER_54_364 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_decap_4 FILLER_54_374 ();
 sg13g2_fill_1 FILLER_54_378 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_4 FILLER_55_26 ();
 sg13g2_fill_2 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_71 ();
 sg13g2_fill_2 FILLER_55_78 ();
 sg13g2_fill_2 FILLER_55_114 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_144 ();
 sg13g2_fill_1 FILLER_55_157 ();
 sg13g2_decap_8 FILLER_55_171 ();
 sg13g2_decap_4 FILLER_55_178 ();
 sg13g2_fill_1 FILLER_55_193 ();
 sg13g2_decap_8 FILLER_55_199 ();
 sg13g2_fill_2 FILLER_55_206 ();
 sg13g2_fill_1 FILLER_55_208 ();
 sg13g2_decap_8 FILLER_55_218 ();
 sg13g2_decap_4 FILLER_55_225 ();
 sg13g2_fill_1 FILLER_55_292 ();
 sg13g2_decap_8 FILLER_55_297 ();
 sg13g2_decap_8 FILLER_55_304 ();
 sg13g2_decap_8 FILLER_55_311 ();
 sg13g2_decap_8 FILLER_55_318 ();
 sg13g2_fill_2 FILLER_55_325 ();
 sg13g2_fill_2 FILLER_55_333 ();
 sg13g2_decap_8 FILLER_55_339 ();
 sg13g2_decap_8 FILLER_55_346 ();
 sg13g2_decap_8 FILLER_55_353 ();
 sg13g2_fill_2 FILLER_55_384 ();
 sg13g2_decap_4 FILLER_55_391 ();
 sg13g2_fill_1 FILLER_55_395 ();
 sg13g2_decap_4 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_4 ();
 sg13g2_fill_2 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_48 ();
 sg13g2_decap_8 FILLER_56_55 ();
 sg13g2_decap_8 FILLER_56_62 ();
 sg13g2_decap_8 FILLER_56_69 ();
 sg13g2_decap_8 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_83 ();
 sg13g2_decap_8 FILLER_56_107 ();
 sg13g2_decap_8 FILLER_56_114 ();
 sg13g2_fill_1 FILLER_56_138 ();
 sg13g2_decap_4 FILLER_56_162 ();
 sg13g2_fill_2 FILLER_56_166 ();
 sg13g2_decap_8 FILLER_56_172 ();
 sg13g2_decap_8 FILLER_56_179 ();
 sg13g2_fill_1 FILLER_56_186 ();
 sg13g2_decap_8 FILLER_56_191 ();
 sg13g2_decap_8 FILLER_56_198 ();
 sg13g2_decap_4 FILLER_56_205 ();
 sg13g2_decap_4 FILLER_56_235 ();
 sg13g2_fill_2 FILLER_56_239 ();
 sg13g2_decap_4 FILLER_56_246 ();
 sg13g2_decap_8 FILLER_56_276 ();
 sg13g2_fill_1 FILLER_56_309 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_fill_2 FILLER_56_338 ();
 sg13g2_fill_1 FILLER_56_340 ();
 sg13g2_fill_1 FILLER_56_354 ();
 sg13g2_decap_4 FILLER_56_364 ();
 sg13g2_fill_2 FILLER_56_368 ();
 sg13g2_decap_8 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_fill_1 FILLER_56_387 ();
 sg13g2_fill_2 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_15 ();
 sg13g2_fill_2 FILLER_57_19 ();
 sg13g2_decap_8 FILLER_57_36 ();
 sg13g2_fill_1 FILLER_57_43 ();
 sg13g2_decap_8 FILLER_57_59 ();
 sg13g2_decap_4 FILLER_57_66 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_fill_2 FILLER_57_102 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_126 ();
 sg13g2_fill_1 FILLER_57_128 ();
 sg13g2_decap_4 FILLER_57_133 ();
 sg13g2_fill_2 FILLER_57_137 ();
 sg13g2_fill_1 FILLER_57_145 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_decap_4 FILLER_57_189 ();
 sg13g2_decap_4 FILLER_57_203 ();
 sg13g2_fill_2 FILLER_57_216 ();
 sg13g2_fill_1 FILLER_57_218 ();
 sg13g2_decap_4 FILLER_57_242 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_fill_2 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_fill_2 FILLER_57_322 ();
 sg13g2_fill_1 FILLER_57_324 ();
 sg13g2_decap_4 FILLER_57_371 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_decap_4 FILLER_57_385 ();
 sg13g2_fill_2 FILLER_57_389 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_11 ();
 sg13g2_fill_2 FILLER_58_28 ();
 sg13g2_fill_1 FILLER_58_60 ();
 sg13g2_fill_1 FILLER_58_152 ();
 sg13g2_fill_1 FILLER_58_168 ();
 sg13g2_fill_1 FILLER_58_196 ();
 sg13g2_fill_1 FILLER_58_231 ();
 sg13g2_decap_4 FILLER_58_240 ();
 sg13g2_fill_2 FILLER_58_244 ();
 sg13g2_decap_8 FILLER_58_274 ();
 sg13g2_decap_4 FILLER_58_281 ();
 sg13g2_fill_1 FILLER_58_285 ();
 sg13g2_decap_8 FILLER_58_314 ();
 sg13g2_decap_8 FILLER_58_321 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_59_31 ();
 sg13g2_fill_1 FILLER_59_33 ();
 sg13g2_fill_2 FILLER_59_63 ();
 sg13g2_fill_1 FILLER_59_91 ();
 sg13g2_decap_4 FILLER_59_120 ();
 sg13g2_decap_4 FILLER_59_128 ();
 sg13g2_fill_1 FILLER_59_132 ();
 sg13g2_decap_4 FILLER_59_150 ();
 sg13g2_fill_2 FILLER_59_154 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_decap_8 FILLER_59_228 ();
 sg13g2_fill_2 FILLER_59_243 ();
 sg13g2_fill_1 FILLER_59_245 ();
 sg13g2_fill_1 FILLER_59_257 ();
 sg13g2_fill_2 FILLER_59_326 ();
 sg13g2_fill_1 FILLER_59_328 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_fill_1 FILLER_59_350 ();
 sg13g2_decap_8 FILLER_59_355 ();
 sg13g2_decap_4 FILLER_59_362 ();
 sg13g2_fill_1 FILLER_59_366 ();
 sg13g2_decap_4 FILLER_59_376 ();
 sg13g2_decap_4 FILLER_59_384 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_23 ();
 sg13g2_decap_4 FILLER_60_30 ();
 sg13g2_fill_2 FILLER_60_34 ();
 sg13g2_fill_2 FILLER_60_55 ();
 sg13g2_fill_1 FILLER_60_62 ();
 sg13g2_fill_1 FILLER_60_72 ();
 sg13g2_fill_1 FILLER_60_86 ();
 sg13g2_fill_1 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_115 ();
 sg13g2_decap_8 FILLER_60_122 ();
 sg13g2_decap_8 FILLER_60_129 ();
 sg13g2_decap_8 FILLER_60_141 ();
 sg13g2_fill_1 FILLER_60_148 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_4 FILLER_60_161 ();
 sg13g2_decap_4 FILLER_60_173 ();
 sg13g2_fill_2 FILLER_60_177 ();
 sg13g2_fill_2 FILLER_60_188 ();
 sg13g2_fill_1 FILLER_60_190 ();
 sg13g2_fill_2 FILLER_60_208 ();
 sg13g2_decap_8 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_225 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_253 ();
 sg13g2_fill_1 FILLER_60_275 ();
 sg13g2_fill_1 FILLER_60_292 ();
 sg13g2_decap_8 FILLER_60_314 ();
 sg13g2_decap_8 FILLER_60_321 ();
 sg13g2_decap_8 FILLER_60_328 ();
 sg13g2_fill_1 FILLER_60_335 ();
 sg13g2_decap_8 FILLER_60_340 ();
 sg13g2_decap_8 FILLER_60_347 ();
 sg13g2_fill_1 FILLER_60_354 ();
 sg13g2_fill_1 FILLER_60_367 ();
 sg13g2_decap_4 FILLER_60_385 ();
 sg13g2_fill_1 FILLER_60_389 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_14 ();
 sg13g2_fill_2 FILLER_61_18 ();
 sg13g2_decap_8 FILLER_61_24 ();
 sg13g2_decap_8 FILLER_61_40 ();
 sg13g2_fill_1 FILLER_61_47 ();
 sg13g2_fill_2 FILLER_61_54 ();
 sg13g2_fill_1 FILLER_61_56 ();
 sg13g2_decap_4 FILLER_61_83 ();
 sg13g2_decap_4 FILLER_61_91 ();
 sg13g2_decap_4 FILLER_61_118 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_142 ();
 sg13g2_decap_8 FILLER_61_148 ();
 sg13g2_decap_8 FILLER_61_155 ();
 sg13g2_decap_8 FILLER_61_162 ();
 sg13g2_decap_4 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_fill_2 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_220 ();
 sg13g2_fill_1 FILLER_61_255 ();
 sg13g2_fill_2 FILLER_61_275 ();
 sg13g2_fill_1 FILLER_61_277 ();
 sg13g2_fill_2 FILLER_61_292 ();
 sg13g2_decap_4 FILLER_61_306 ();
 sg13g2_fill_2 FILLER_61_310 ();
 sg13g2_decap_4 FILLER_61_347 ();
 sg13g2_fill_1 FILLER_61_351 ();
 sg13g2_fill_1 FILLER_61_365 ();
 sg13g2_decap_4 FILLER_61_372 ();
 sg13g2_fill_2 FILLER_61_376 ();
 sg13g2_fill_2 FILLER_61_388 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_17 ();
 sg13g2_fill_1 FILLER_62_19 ();
 sg13g2_fill_1 FILLER_62_40 ();
 sg13g2_fill_1 FILLER_62_47 ();
 sg13g2_fill_1 FILLER_62_88 ();
 sg13g2_fill_2 FILLER_62_97 ();
 sg13g2_fill_2 FILLER_62_158 ();
 sg13g2_fill_2 FILLER_62_174 ();
 sg13g2_fill_1 FILLER_62_176 ();
 sg13g2_fill_2 FILLER_62_182 ();
 sg13g2_fill_2 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_195 ();
 sg13g2_fill_1 FILLER_62_205 ();
 sg13g2_fill_2 FILLER_62_243 ();
 sg13g2_fill_2 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_302 ();
 sg13g2_fill_1 FILLER_62_304 ();
 sg13g2_fill_1 FILLER_62_321 ();
 sg13g2_decap_8 FILLER_62_326 ();
 sg13g2_decap_8 FILLER_62_333 ();
 sg13g2_decap_8 FILLER_62_340 ();
 sg13g2_fill_1 FILLER_62_347 ();
 sg13g2_decap_4 FILLER_62_374 ();
 sg13g2_fill_1 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_384 ();
 sg13g2_decap_4 FILLER_62_404 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_17 ();
 sg13g2_decap_4 FILLER_63_54 ();
 sg13g2_fill_1 FILLER_63_58 ();
 sg13g2_fill_1 FILLER_63_80 ();
 sg13g2_fill_2 FILLER_63_100 ();
 sg13g2_fill_1 FILLER_63_124 ();
 sg13g2_fill_1 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_227 ();
 sg13g2_fill_1 FILLER_63_229 ();
 sg13g2_decap_8 FILLER_63_251 ();
 sg13g2_decap_8 FILLER_63_258 ();
 sg13g2_decap_4 FILLER_63_265 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_decap_8 FILLER_63_325 ();
 sg13g2_decap_8 FILLER_63_332 ();
 sg13g2_fill_2 FILLER_63_339 ();
 sg13g2_fill_1 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_352 ();
 sg13g2_fill_2 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_360 ();
 sg13g2_fill_2 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_fill_1 FILLER_64_32 ();
 sg13g2_fill_2 FILLER_64_43 ();
 sg13g2_decap_4 FILLER_64_51 ();
 sg13g2_decap_8 FILLER_64_65 ();
 sg13g2_fill_1 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_103 ();
 sg13g2_fill_2 FILLER_64_121 ();
 sg13g2_fill_2 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_167 ();
 sg13g2_fill_1 FILLER_64_174 ();
 sg13g2_decap_8 FILLER_64_213 ();
 sg13g2_decap_4 FILLER_64_225 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_16 ();
 sg13g2_decap_8 FILLER_65_40 ();
 sg13g2_fill_2 FILLER_65_47 ();
 sg13g2_fill_1 FILLER_65_49 ();
 sg13g2_fill_1 FILLER_65_68 ();
 sg13g2_decap_8 FILLER_65_78 ();
 sg13g2_fill_2 FILLER_65_85 ();
 sg13g2_fill_1 FILLER_65_87 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_fill_2 FILLER_65_119 ();
 sg13g2_fill_2 FILLER_65_126 ();
 sg13g2_fill_1 FILLER_65_128 ();
 sg13g2_decap_8 FILLER_65_152 ();
 sg13g2_decap_8 FILLER_65_159 ();
 sg13g2_decap_8 FILLER_65_166 ();
 sg13g2_decap_8 FILLER_65_173 ();
 sg13g2_decap_8 FILLER_65_180 ();
 sg13g2_decap_8 FILLER_65_187 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_fill_2 FILLER_65_245 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_decap_8 FILLER_65_261 ();
 sg13g2_fill_2 FILLER_65_268 ();
 sg13g2_decap_4 FILLER_65_275 ();
 sg13g2_fill_2 FILLER_65_279 ();
 sg13g2_decap_4 FILLER_65_285 ();
 sg13g2_fill_2 FILLER_65_289 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_fill_1 FILLER_65_306 ();
 sg13g2_fill_2 FILLER_65_312 ();
 sg13g2_fill_1 FILLER_65_314 ();
 sg13g2_decap_4 FILLER_65_336 ();
 sg13g2_fill_2 FILLER_65_350 ();
 sg13g2_fill_1 FILLER_65_352 ();
 sg13g2_decap_4 FILLER_65_372 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_11 ();
 sg13g2_decap_8 FILLER_66_16 ();
 sg13g2_fill_2 FILLER_66_23 ();
 sg13g2_fill_1 FILLER_66_25 ();
 sg13g2_decap_8 FILLER_66_34 ();
 sg13g2_decap_8 FILLER_66_41 ();
 sg13g2_decap_4 FILLER_66_48 ();
 sg13g2_decap_4 FILLER_66_82 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_decap_4 FILLER_66_107 ();
 sg13g2_fill_1 FILLER_66_111 ();
 sg13g2_decap_4 FILLER_66_116 ();
 sg13g2_fill_1 FILLER_66_137 ();
 sg13g2_decap_8 FILLER_66_181 ();
 sg13g2_decap_8 FILLER_66_188 ();
 sg13g2_decap_8 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_202 ();
 sg13g2_fill_2 FILLER_66_210 ();
 sg13g2_fill_1 FILLER_66_238 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_decap_8 FILLER_66_264 ();
 sg13g2_fill_2 FILLER_66_271 ();
 sg13g2_fill_1 FILLER_66_273 ();
 sg13g2_decap_4 FILLER_66_279 ();
 sg13g2_fill_1 FILLER_66_283 ();
 sg13g2_decap_8 FILLER_66_293 ();
 sg13g2_fill_1 FILLER_66_326 ();
 sg13g2_decap_8 FILLER_66_332 ();
 sg13g2_decap_8 FILLER_66_339 ();
 sg13g2_decap_8 FILLER_66_346 ();
 sg13g2_decap_8 FILLER_66_353 ();
 sg13g2_decap_4 FILLER_66_360 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_decap_4 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_398 ();
 sg13g2_decap_4 FILLER_66_405 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_25 ();
 sg13g2_fill_2 FILLER_67_31 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_decap_8 FILLER_67_68 ();
 sg13g2_fill_2 FILLER_67_75 ();
 sg13g2_decap_4 FILLER_67_111 ();
 sg13g2_fill_1 FILLER_67_115 ();
 sg13g2_fill_2 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_123 ();
 sg13g2_fill_2 FILLER_67_128 ();
 sg13g2_decap_4 FILLER_67_135 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_fill_2 FILLER_67_196 ();
 sg13g2_fill_1 FILLER_67_198 ();
 sg13g2_decap_4 FILLER_67_205 ();
 sg13g2_decap_8 FILLER_67_213 ();
 sg13g2_fill_2 FILLER_67_220 ();
 sg13g2_fill_1 FILLER_67_231 ();
 sg13g2_fill_1 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_341 ();
 sg13g2_decap_8 FILLER_67_348 ();
 sg13g2_decap_8 FILLER_67_355 ();
 sg13g2_decap_8 FILLER_67_362 ();
 sg13g2_decap_8 FILLER_67_369 ();
 sg13g2_decap_8 FILLER_67_376 ();
 sg13g2_decap_8 FILLER_67_383 ();
 sg13g2_decap_8 FILLER_67_390 ();
 sg13g2_decap_8 FILLER_67_397 ();
 sg13g2_decap_4 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_68_48 ();
 sg13g2_fill_1 FILLER_68_50 ();
 sg13g2_fill_2 FILLER_68_94 ();
 sg13g2_decap_8 FILLER_68_100 ();
 sg13g2_decap_4 FILLER_68_114 ();
 sg13g2_fill_2 FILLER_68_126 ();
 sg13g2_fill_2 FILLER_68_144 ();
 sg13g2_decap_4 FILLER_68_173 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_221 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_decap_4 FILLER_68_234 ();
 sg13g2_fill_2 FILLER_68_238 ();
 sg13g2_decap_4 FILLER_68_248 ();
 sg13g2_fill_2 FILLER_68_264 ();
 sg13g2_fill_2 FILLER_68_278 ();
 sg13g2_decap_4 FILLER_68_294 ();
 sg13g2_fill_1 FILLER_68_298 ();
 sg13g2_decap_4 FILLER_68_309 ();
 sg13g2_fill_2 FILLER_68_353 ();
 sg13g2_fill_1 FILLER_68_355 ();
 sg13g2_decap_8 FILLER_68_360 ();
 sg13g2_fill_2 FILLER_68_367 ();
 sg13g2_decap_8 FILLER_68_374 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_2 ();
 sg13g2_decap_8 FILLER_69_67 ();
 sg13g2_decap_4 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_78 ();
 sg13g2_fill_2 FILLER_69_83 ();
 sg13g2_decap_8 FILLER_69_89 ();
 sg13g2_fill_2 FILLER_69_131 ();
 sg13g2_fill_1 FILLER_69_138 ();
 sg13g2_fill_2 FILLER_69_207 ();
 sg13g2_fill_1 FILLER_69_209 ();
 sg13g2_fill_2 FILLER_69_214 ();
 sg13g2_fill_1 FILLER_69_216 ();
 sg13g2_fill_2 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_228 ();
 sg13g2_fill_1 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_242 ();
 sg13g2_fill_2 FILLER_69_262 ();
 sg13g2_decap_4 FILLER_69_292 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_fill_1 FILLER_69_319 ();
 sg13g2_fill_2 FILLER_69_363 ();
 sg13g2_fill_1 FILLER_69_365 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_9 ();
 sg13g2_fill_1 FILLER_70_22 ();
 sg13g2_fill_1 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_39 ();
 sg13g2_fill_1 FILLER_70_46 ();
 sg13g2_fill_2 FILLER_70_51 ();
 sg13g2_fill_1 FILLER_70_89 ();
 sg13g2_fill_2 FILLER_70_95 ();
 sg13g2_fill_1 FILLER_70_97 ();
 sg13g2_decap_8 FILLER_70_103 ();
 sg13g2_decap_4 FILLER_70_110 ();
 sg13g2_fill_1 FILLER_70_114 ();
 sg13g2_fill_2 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_fill_1 FILLER_70_164 ();
 sg13g2_fill_2 FILLER_70_180 ();
 sg13g2_fill_1 FILLER_70_182 ();
 sg13g2_decap_4 FILLER_70_200 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_decap_8 FILLER_70_258 ();
 sg13g2_decap_4 FILLER_70_265 ();
 sg13g2_fill_1 FILLER_70_269 ();
 sg13g2_decap_8 FILLER_70_291 ();
 sg13g2_decap_8 FILLER_70_298 ();
 sg13g2_decap_4 FILLER_70_305 ();
 sg13g2_fill_1 FILLER_70_309 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_decap_4 FILLER_70_343 ();
 sg13g2_fill_2 FILLER_70_369 ();
 sg13g2_fill_2 FILLER_70_376 ();
 sg13g2_fill_1 FILLER_70_378 ();
 sg13g2_fill_2 FILLER_70_388 ();
 sg13g2_fill_1 FILLER_70_390 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_4 ();
 sg13g2_fill_1 FILLER_71_23 ();
 sg13g2_fill_2 FILLER_71_33 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_fill_1 FILLER_71_53 ();
 sg13g2_fill_2 FILLER_71_113 ();
 sg13g2_fill_1 FILLER_71_115 ();
 sg13g2_fill_2 FILLER_71_142 ();
 sg13g2_fill_2 FILLER_71_148 ();
 sg13g2_decap_8 FILLER_71_157 ();
 sg13g2_decap_4 FILLER_71_164 ();
 sg13g2_fill_1 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_178 ();
 sg13g2_decap_8 FILLER_71_185 ();
 sg13g2_fill_2 FILLER_71_192 ();
 sg13g2_fill_2 FILLER_71_225 ();
 sg13g2_fill_1 FILLER_71_227 ();
 sg13g2_decap_4 FILLER_71_237 ();
 sg13g2_decap_8 FILLER_71_271 ();
 sg13g2_fill_2 FILLER_71_278 ();
 sg13g2_decap_4 FILLER_71_307 ();
 sg13g2_fill_2 FILLER_71_311 ();
 sg13g2_fill_2 FILLER_71_322 ();
 sg13g2_fill_1 FILLER_71_324 ();
 sg13g2_fill_2 FILLER_71_351 ();
 sg13g2_fill_2 FILLER_71_387 ();
 sg13g2_decap_4 FILLER_71_393 ();
 sg13g2_fill_1 FILLER_71_397 ();
 sg13g2_decap_4 FILLER_72_45 ();
 sg13g2_fill_2 FILLER_72_97 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_fill_2 FILLER_72_115 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_fill_2 FILLER_72_138 ();
 sg13g2_fill_1 FILLER_72_140 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_4 FILLER_72_214 ();
 sg13g2_fill_1 FILLER_72_218 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_fill_2 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_fill_2 FILLER_72_267 ();
 sg13g2_fill_1 FILLER_72_269 ();
 sg13g2_decap_4 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_decap_8 FILLER_72_319 ();
 sg13g2_fill_2 FILLER_72_326 ();
 sg13g2_fill_1 FILLER_72_328 ();
 sg13g2_fill_1 FILLER_72_338 ();
 sg13g2_fill_2 FILLER_72_347 ();
 sg13g2_fill_1 FILLER_72_368 ();
 sg13g2_decap_4 FILLER_72_374 ();
 sg13g2_decap_4 FILLER_72_404 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_15 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_decap_4 FILLER_73_59 ();
 sg13g2_fill_2 FILLER_73_100 ();
 sg13g2_fill_1 FILLER_73_102 ();
 sg13g2_fill_2 FILLER_73_169 ();
 sg13g2_fill_1 FILLER_73_197 ();
 sg13g2_decap_8 FILLER_73_212 ();
 sg13g2_fill_1 FILLER_73_219 ();
 sg13g2_fill_1 FILLER_73_241 ();
 sg13g2_decap_4 FILLER_73_290 ();
 sg13g2_fill_2 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_299 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_fill_2 FILLER_73_329 ();
 sg13g2_fill_1 FILLER_73_331 ();
 sg13g2_decap_8 FILLER_73_337 ();
 sg13g2_fill_2 FILLER_73_344 ();
 sg13g2_fill_1 FILLER_73_346 ();
 sg13g2_fill_2 FILLER_73_362 ();
 sg13g2_fill_1 FILLER_73_364 ();
 sg13g2_decap_4 FILLER_74_40 ();
 sg13g2_fill_2 FILLER_74_48 ();
 sg13g2_fill_1 FILLER_74_50 ();
 sg13g2_fill_2 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_58 ();
 sg13g2_fill_2 FILLER_74_64 ();
 sg13g2_fill_1 FILLER_74_66 ();
 sg13g2_fill_1 FILLER_74_91 ();
 sg13g2_fill_2 FILLER_74_128 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_decap_4 FILLER_74_172 ();
 sg13g2_decap_8 FILLER_74_186 ();
 sg13g2_fill_2 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_263 ();
 sg13g2_decap_8 FILLER_74_268 ();
 sg13g2_fill_2 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_277 ();
 sg13g2_decap_4 FILLER_74_290 ();
 sg13g2_decap_8 FILLER_74_333 ();
 sg13g2_fill_2 FILLER_74_340 ();
 sg13g2_fill_1 FILLER_74_342 ();
 sg13g2_decap_8 FILLER_74_349 ();
 sg13g2_fill_2 FILLER_74_356 ();
 sg13g2_fill_1 FILLER_74_358 ();
 sg13g2_fill_1 FILLER_74_374 ();
 sg13g2_fill_2 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_15 ();
 sg13g2_decap_8 FILLER_75_40 ();
 sg13g2_decap_4 FILLER_75_47 ();
 sg13g2_decap_4 FILLER_75_56 ();
 sg13g2_decap_4 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_78 ();
 sg13g2_decap_8 FILLER_75_85 ();
 sg13g2_fill_2 FILLER_75_92 ();
 sg13g2_fill_1 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_108 ();
 sg13g2_fill_1 FILLER_75_127 ();
 sg13g2_fill_2 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_172 ();
 sg13g2_fill_2 FILLER_75_185 ();
 sg13g2_decap_8 FILLER_75_192 ();
 sg13g2_decap_4 FILLER_75_204 ();
 sg13g2_fill_1 FILLER_75_208 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_decap_8 FILLER_75_220 ();
 sg13g2_decap_4 FILLER_75_227 ();
 sg13g2_fill_1 FILLER_75_236 ();
 sg13g2_fill_2 FILLER_75_251 ();
 sg13g2_fill_1 FILLER_75_253 ();
 sg13g2_fill_2 FILLER_75_317 ();
 sg13g2_fill_2 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_342 ();
 sg13g2_fill_2 FILLER_75_366 ();
 sg13g2_fill_1 FILLER_75_368 ();
 sg13g2_decap_4 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_12 ();
 sg13g2_fill_2 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_99 ();
 sg13g2_fill_1 FILLER_76_106 ();
 sg13g2_fill_2 FILLER_76_122 ();
 sg13g2_fill_1 FILLER_76_145 ();
 sg13g2_fill_1 FILLER_76_172 ();
 sg13g2_decap_8 FILLER_76_186 ();
 sg13g2_decap_8 FILLER_76_202 ();
 sg13g2_fill_2 FILLER_76_209 ();
 sg13g2_fill_1 FILLER_76_211 ();
 sg13g2_fill_1 FILLER_76_217 ();
 sg13g2_fill_2 FILLER_76_232 ();
 sg13g2_fill_2 FILLER_76_269 ();
 sg13g2_fill_2 FILLER_76_314 ();
 sg13g2_fill_1 FILLER_76_316 ();
 sg13g2_fill_1 FILLER_76_346 ();
 sg13g2_fill_2 FILLER_76_396 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_4 FILLER_77_7 ();
 sg13g2_fill_1 FILLER_77_57 ();
 sg13g2_fill_2 FILLER_77_64 ();
 sg13g2_decap_8 FILLER_77_102 ();
 sg13g2_fill_2 FILLER_77_109 ();
 sg13g2_fill_1 FILLER_77_111 ();
 sg13g2_fill_2 FILLER_77_207 ();
 sg13g2_fill_2 FILLER_77_240 ();
 sg13g2_fill_1 FILLER_77_242 ();
 sg13g2_fill_2 FILLER_77_281 ();
 sg13g2_fill_1 FILLER_77_283 ();
 sg13g2_fill_2 FILLER_77_301 ();
 sg13g2_fill_1 FILLER_77_373 ();
 sg13g2_fill_2 FILLER_78_26 ();
 sg13g2_fill_1 FILLER_78_67 ();
 sg13g2_fill_2 FILLER_78_182 ();
 sg13g2_fill_2 FILLER_78_250 ();
 sg13g2_fill_1 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_325 ();
 sg13g2_fill_1 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_15 ();
 sg13g2_fill_2 FILLER_79_22 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_fill_2 FILLER_79_35 ();
 sg13g2_fill_1 FILLER_79_51 ();
 sg13g2_fill_2 FILLER_79_67 ();
 sg13g2_fill_1 FILLER_79_69 ();
 sg13g2_decap_4 FILLER_79_106 ();
 sg13g2_fill_2 FILLER_79_110 ();
 sg13g2_fill_1 FILLER_79_129 ();
 sg13g2_fill_1 FILLER_79_139 ();
 sg13g2_fill_1 FILLER_79_160 ();
 sg13g2_decap_4 FILLER_79_174 ();
 sg13g2_decap_8 FILLER_79_204 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_238 ();
 sg13g2_fill_1 FILLER_79_274 ();
 sg13g2_fill_2 FILLER_79_306 ();
 sg13g2_fill_2 FILLER_79_334 ();
 sg13g2_fill_1 FILLER_79_336 ();
 sg13g2_fill_2 FILLER_79_356 ();
 sg13g2_fill_1 FILLER_79_358 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_4 FILLER_80_42 ();
 sg13g2_decap_4 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_decap_8 FILLER_80_110 ();
 sg13g2_fill_1 FILLER_80_117 ();
 sg13g2_decap_8 FILLER_80_125 ();
 sg13g2_decap_8 FILLER_80_132 ();
 sg13g2_decap_8 FILLER_80_139 ();
 sg13g2_decap_8 FILLER_80_146 ();
 sg13g2_fill_1 FILLER_80_153 ();
 sg13g2_decap_4 FILLER_80_158 ();
 sg13g2_decap_8 FILLER_80_166 ();
 sg13g2_decap_8 FILLER_80_173 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_4 FILLER_80_215 ();
 sg13g2_fill_1 FILLER_80_219 ();
 sg13g2_decap_8 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_fill_1 FILLER_80_249 ();
 sg13g2_decap_4 FILLER_80_254 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_fill_2 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_fill_2 FILLER_80_277 ();
 sg13g2_fill_2 FILLER_80_289 ();
 sg13g2_fill_1 FILLER_80_291 ();
 sg13g2_decap_8 FILLER_80_310 ();
 sg13g2_fill_2 FILLER_80_317 ();
 sg13g2_fill_1 FILLER_80_327 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_1 FILLER_80_374 ();
 sg13g2_fill_2 FILLER_80_407 ();
endmodule
