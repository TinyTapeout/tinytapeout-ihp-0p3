module tt_um_calonso88_spi_test (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire \config_regs[0] ;
 wire \config_regs[100] ;
 wire \config_regs[101] ;
 wire \config_regs[102] ;
 wire \config_regs[103] ;
 wire \config_regs[104] ;
 wire \config_regs[105] ;
 wire \config_regs[106] ;
 wire \config_regs[107] ;
 wire \config_regs[108] ;
 wire \config_regs[109] ;
 wire \config_regs[10] ;
 wire \config_regs[110] ;
 wire \config_regs[111] ;
 wire \config_regs[112] ;
 wire \config_regs[113] ;
 wire \config_regs[114] ;
 wire \config_regs[115] ;
 wire \config_regs[116] ;
 wire \config_regs[117] ;
 wire \config_regs[118] ;
 wire \config_regs[119] ;
 wire \config_regs[11] ;
 wire \config_regs[120] ;
 wire \config_regs[121] ;
 wire \config_regs[122] ;
 wire \config_regs[123] ;
 wire \config_regs[124] ;
 wire \config_regs[125] ;
 wire \config_regs[126] ;
 wire \config_regs[127] ;
 wire \config_regs[12] ;
 wire \config_regs[13] ;
 wire \config_regs[14] ;
 wire \config_regs[15] ;
 wire \config_regs[16] ;
 wire \config_regs[17] ;
 wire \config_regs[18] ;
 wire \config_regs[19] ;
 wire \config_regs[1] ;
 wire \config_regs[20] ;
 wire \config_regs[21] ;
 wire \config_regs[22] ;
 wire \config_regs[23] ;
 wire \config_regs[24] ;
 wire \config_regs[25] ;
 wire \config_regs[26] ;
 wire \config_regs[27] ;
 wire \config_regs[28] ;
 wire \config_regs[29] ;
 wire \config_regs[2] ;
 wire \config_regs[30] ;
 wire \config_regs[31] ;
 wire \config_regs[32] ;
 wire \config_regs[33] ;
 wire \config_regs[34] ;
 wire \config_regs[35] ;
 wire \config_regs[36] ;
 wire \config_regs[37] ;
 wire \config_regs[38] ;
 wire \config_regs[39] ;
 wire \config_regs[3] ;
 wire \config_regs[40] ;
 wire \config_regs[41] ;
 wire \config_regs[42] ;
 wire \config_regs[43] ;
 wire \config_regs[44] ;
 wire \config_regs[45] ;
 wire \config_regs[46] ;
 wire \config_regs[47] ;
 wire \config_regs[48] ;
 wire \config_regs[49] ;
 wire \config_regs[4] ;
 wire \config_regs[50] ;
 wire \config_regs[51] ;
 wire \config_regs[52] ;
 wire \config_regs[53] ;
 wire \config_regs[54] ;
 wire \config_regs[55] ;
 wire \config_regs[56] ;
 wire \config_regs[57] ;
 wire \config_regs[58] ;
 wire \config_regs[59] ;
 wire \config_regs[5] ;
 wire \config_regs[60] ;
 wire \config_regs[61] ;
 wire \config_regs[62] ;
 wire \config_regs[63] ;
 wire \config_regs[64] ;
 wire \config_regs[65] ;
 wire \config_regs[66] ;
 wire \config_regs[67] ;
 wire \config_regs[68] ;
 wire \config_regs[69] ;
 wire \config_regs[6] ;
 wire \config_regs[70] ;
 wire \config_regs[71] ;
 wire \config_regs[72] ;
 wire \config_regs[73] ;
 wire \config_regs[74] ;
 wire \config_regs[75] ;
 wire \config_regs[76] ;
 wire \config_regs[77] ;
 wire \config_regs[78] ;
 wire \config_regs[79] ;
 wire \config_regs[7] ;
 wire \config_regs[80] ;
 wire \config_regs[81] ;
 wire \config_regs[82] ;
 wire \config_regs[83] ;
 wire \config_regs[84] ;
 wire \config_regs[85] ;
 wire \config_regs[86] ;
 wire \config_regs[87] ;
 wire \config_regs[88] ;
 wire \config_regs[89] ;
 wire \config_regs[8] ;
 wire \config_regs[90] ;
 wire \config_regs[91] ;
 wire \config_regs[92] ;
 wire \config_regs[93] ;
 wire \config_regs[94] ;
 wire \config_regs[95] ;
 wire \config_regs[96] ;
 wire \config_regs[97] ;
 wire \config_regs[98] ;
 wire \config_regs[99] ;
 wire \config_regs[9] ;
 wire cpha_sync;
 wire cpol_sync;
 wire spi_clk_sync;
 wire spi_cs_n_sync;
 wire spi_miso;
 wire spi_mosi_sync;
 wire \spi_wrapper_i.reg_addr[0] ;
 wire \spi_wrapper_i.reg_addr[1] ;
 wire \spi_wrapper_i.reg_addr[2] ;
 wire \spi_wrapper_i.reg_addr[3] ;
 wire \spi_wrapper_i.reg_addr[4] ;
 wire \spi_wrapper_i.reg_data_o[0] ;
 wire \spi_wrapper_i.reg_data_o[1] ;
 wire \spi_wrapper_i.reg_data_o[2] ;
 wire \spi_wrapper_i.reg_data_o[3] ;
 wire \spi_wrapper_i.reg_data_o[4] ;
 wire \spi_wrapper_i.reg_data_o[5] ;
 wire \spi_wrapper_i.reg_data_o[6] ;
 wire \spi_wrapper_i.reg_data_o[7] ;
 wire \spi_wrapper_i.reg_data_o_vld ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.buffer_counter[3] ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.reg_rw ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[7] ;
 wire \spi_wrapper_i.spi_reg_inst.state[0] ;
 wire \spi_wrapper_i.spi_reg_inst.state[1] ;
 wire \spi_wrapper_i.spi_reg_inst.state[2] ;
 wire \spi_wrapper_i.spi_reg_inst.state[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[6] ;
 wire \synchronizer_spi_clk_inst.data_sync[1] ;
 wire \synchronizer_spi_cs_n_inst.data_sync[1] ;
 wire \synchronizer_spi_mode_cpha.data_sync[1] ;
 wire \synchronizer_spi_mode_cpol.data_sync[1] ;
 wire \synchronizer_spi_mosi_inst.data_sync[1] ;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;

 sg13g2_inv_1 _0576_ (.Y(_0196_),
    .A(net349));
 sg13g2_inv_1 _0577_ (.Y(_0197_),
    .A(net47));
 sg13g2_inv_1 _0578_ (.Y(_0198_),
    .A(net21));
 sg13g2_inv_1 _0579_ (.Y(_0199_),
    .A(net31));
 sg13g2_inv_2 _0580_ (.Y(_0200_),
    .A(net302));
 sg13g2_nor3_2 _0581_ (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ),
    .B(\spi_wrapper_i.spi_reg_inst.buffer_counter[0] ),
    .C(\spi_wrapper_i.spi_reg_inst.buffer_counter[2] ),
    .Y(_0201_));
 sg13g2_and2_2 _0582_ (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ),
    .B(_0201_),
    .X(_0202_));
 sg13g2_nor2b_1 _0583_ (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .B_N(spi_cs_n_sync),
    .Y(_0203_));
 sg13g2_o21ai_1 _0584_ (.B1(_0203_),
    .Y(_0204_),
    .A1(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .A2(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_or2_1 _0585_ (.X(_0205_),
    .B(_0204_),
    .A(_0202_));
 sg13g2_nor2b_2 _0586_ (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ),
    .B_N(_0201_),
    .Y(_0206_));
 sg13g2_o21ai_1 _0587_ (.B1(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .Y(_0207_),
    .A1(_0201_),
    .A2(_0203_));
 sg13g2_o21ai_1 _0588_ (.B1(_0205_),
    .Y(_0208_),
    .A1(_0206_),
    .A2(_0207_));
 sg13g2_nand2_1 _0589_ (.Y(_0209_),
    .A(net334),
    .B(_0202_));
 sg13g2_nand3_1 _0590_ (.B(net177),
    .C(_0202_),
    .A(net334),
    .Y(_0210_));
 sg13g2_nor2b_1 _0591_ (.A(spi_cs_n_sync),
    .B_N(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .Y(_0211_));
 sg13g2_inv_1 _0592_ (.Y(_0212_),
    .A(_0211_));
 sg13g2_nand2_1 _0593_ (.Y(_0213_),
    .A(net335),
    .B(_0211_));
 sg13g2_a22oi_1 _0594_ (.Y(_0214_),
    .B1(_0213_),
    .B2(net21),
    .A2(_0208_),
    .A1(net334));
 sg13g2_and2_1 _0595_ (.A(net261),
    .B(_0214_),
    .X(_0020_));
 sg13g2_nand3_1 _0596_ (.B(net224),
    .C(_0202_),
    .A(net334),
    .Y(_0215_));
 sg13g2_o21ai_1 _0597_ (.B1(net260),
    .Y(_0001_),
    .A1(net334),
    .A2(_0197_));
 sg13g2_o21ai_1 _0598_ (.B1(net334),
    .Y(_0216_),
    .A1(_0202_),
    .A2(_0203_));
 sg13g2_nand2_1 _0599_ (.Y(_0217_),
    .A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .B(_0216_));
 sg13g2_o21ai_1 _0600_ (.B1(_0217_),
    .Y(_0002_),
    .A1(_0198_),
    .A2(_0213_));
 sg13g2_nand2_1 _0601_ (.Y(_0218_),
    .A(net177),
    .B(_0216_));
 sg13g2_nand2_1 _0602_ (.Y(_0219_),
    .A(net334),
    .B(net47));
 sg13g2_o21ai_1 _0603_ (.B1(_0218_),
    .Y(_0003_),
    .A1(_0199_),
    .A2(_0219_));
 sg13g2_and2_1 _0604_ (.A(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_0206_),
    .X(_0220_));
 sg13g2_nand2_2 _0605_ (.Y(_0221_),
    .A(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_0206_));
 sg13g2_a21oi_1 _0606_ (.A1(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .A2(_0216_),
    .Y(_0222_),
    .B1(_0220_));
 sg13g2_o21ai_1 _0607_ (.B1(_0222_),
    .Y(_0000_),
    .A1(net31),
    .A2(_0219_));
 sg13g2_xnor2_1 _0608_ (.Y(_0223_),
    .A(cpha_sync),
    .B(cpol_sync));
 sg13g2_nand3b_1 _0609_ (.B(uio_oe[3]),
    .C(spi_clk_sync),
    .Y(_0224_),
    .A_N(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_nand2_1 _0610_ (.Y(_0225_),
    .A(_0223_),
    .B(_0224_));
 sg13g2_nand3b_1 _0611_ (.B(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .C(uio_oe[3]),
    .Y(_0226_),
    .A_N(spi_clk_sync));
 sg13g2_nand2b_1 _0612_ (.Y(_0227_),
    .B(_0226_),
    .A_N(_0223_));
 sg13g2_nand3_1 _0613_ (.B(_0225_),
    .C(_0227_),
    .A(net336),
    .Y(_0228_));
 sg13g2_nor2_2 _0614_ (.A(_0196_),
    .B(net257),
    .Y(_0229_));
 sg13g2_or2_1 _0615_ (.X(_0230_),
    .B(net256),
    .A(_0202_));
 sg13g2_a21oi_1 _0616_ (.A1(_0196_),
    .A2(_0230_),
    .Y(_0021_),
    .B1(_0229_));
 sg13g2_xor2_1 _0617_ (.B(_0229_),
    .A(net342),
    .X(_0022_));
 sg13g2_a21oi_1 _0618_ (.A1(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ),
    .A2(_0229_),
    .Y(_0231_),
    .B1(net248));
 sg13g2_and2_1 _0619_ (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ),
    .B(net248),
    .X(_0232_));
 sg13g2_a21oi_1 _0620_ (.A1(_0229_),
    .A2(_0232_),
    .Y(_0023_),
    .B1(net249));
 sg13g2_nand3_1 _0621_ (.B(_0209_),
    .C(net256),
    .A(net348),
    .Y(_0233_));
 sg13g2_nand2_1 _0622_ (.Y(_0234_),
    .A(net349),
    .B(_0232_));
 sg13g2_xor2_1 _0623_ (.B(_0234_),
    .A(net348),
    .X(_0235_));
 sg13g2_o21ai_1 _0624_ (.B1(_0233_),
    .Y(_0024_),
    .A1(_0230_),
    .A2(_0235_));
 sg13g2_nor2_1 _0625_ (.A(net203),
    .B(net260),
    .Y(_0236_));
 sg13g2_a21oi_1 _0626_ (.A1(_0199_),
    .A2(net260),
    .Y(_0025_),
    .B1(_0236_));
 sg13g2_mux2_1 _0627_ (.A0(net245),
    .A1(net350),
    .S(net260),
    .X(_0026_));
 sg13g2_mux2_1 _0628_ (.A0(net229),
    .A1(net339),
    .S(_0215_),
    .X(_0027_));
 sg13g2_mux2_1 _0629_ (.A0(net172),
    .A1(net207),
    .S(net260),
    .X(_0028_));
 sg13g2_mux2_1 _0630_ (.A0(net344),
    .A1(net346),
    .S(net260),
    .X(_0029_));
 sg13g2_nor2_1 _0631_ (.A(net225),
    .B(net260),
    .Y(_0237_));
 sg13g2_a21oi_1 _0632_ (.A1(_0200_),
    .A2(net260),
    .Y(_0030_),
    .B1(_0237_));
 sg13g2_nand2b_1 _0633_ (.Y(_0238_),
    .B(net37),
    .A_N(net334));
 sg13g2_o21ai_1 _0634_ (.B1(_0238_),
    .Y(_0031_),
    .A1(_0199_),
    .A2(net261));
 sg13g2_mux2_1 _0635_ (.A0(net245),
    .A1(net300),
    .S(net261),
    .X(_0032_));
 sg13g2_mux2_1 _0636_ (.A0(net229),
    .A1(net299),
    .S(_0210_),
    .X(_0033_));
 sg13g2_mux2_1 _0637_ (.A0(net172),
    .A1(net296),
    .S(net261),
    .X(_0034_));
 sg13g2_mux2_1 _0638_ (.A0(net344),
    .A1(net294),
    .S(_0210_),
    .X(_0035_));
 sg13g2_mux2_1 _0639_ (.A0(net225),
    .A1(net292),
    .S(net261),
    .X(_0036_));
 sg13g2_mux2_1 _0640_ (.A0(net189),
    .A1(net290),
    .S(net261),
    .X(_0037_));
 sg13g2_mux2_1 _0641_ (.A0(net192),
    .A1(net288),
    .S(net261),
    .X(_0038_));
 sg13g2_mux2_1 _0642_ (.A0(net203),
    .A1(net285),
    .S(net261),
    .X(_0039_));
 sg13g2_mux2_1 _0643_ (.A0(_0224_),
    .A1(_0226_),
    .S(_0223_),
    .X(_0239_));
 sg13g2_nand2_1 _0644_ (.Y(_0240_),
    .A(_0221_),
    .B(_0239_));
 sg13g2_o21ai_1 _0645_ (.B1(net336),
    .Y(_0241_),
    .A1(_0211_),
    .A2(_0240_));
 sg13g2_nand2_1 _0646_ (.Y(_0242_),
    .A(net27),
    .B(_0241_));
 sg13g2_nor2b_2 _0647_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B_N(\spi_wrapper_i.reg_addr[3] ),
    .Y(_0243_));
 sg13g2_nor2b_2 _0648_ (.A(\spi_wrapper_i.reg_addr[1] ),
    .B_N(\spi_wrapper_i.reg_addr[0] ),
    .Y(_0244_));
 sg13g2_and2_1 _0649_ (.A(_0243_),
    .B(_0244_),
    .X(_0245_));
 sg13g2_nor2_2 _0650_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(\spi_wrapper_i.reg_addr[3] ),
    .Y(_0246_));
 sg13g2_nor2b_2 _0651_ (.A(\spi_wrapper_i.reg_addr[0] ),
    .B_N(\spi_wrapper_i.reg_addr[1] ),
    .Y(_0247_));
 sg13g2_and2_2 _0652_ (.A(_0246_),
    .B(_0247_),
    .X(_0248_));
 sg13g2_a22oi_1 _0653_ (.Y(_0249_),
    .B1(_0248_),
    .B2(\config_regs[16] ),
    .A2(_0245_),
    .A1(\config_regs[72] ));
 sg13g2_and2_1 _0654_ (.A(\spi_wrapper_i.reg_addr[2] ),
    .B(\spi_wrapper_i.reg_addr[3] ),
    .X(_0250_));
 sg13g2_and2_1 _0655_ (.A(_0244_),
    .B(_0250_),
    .X(_0251_));
 sg13g2_nor2b_2 _0656_ (.A(\spi_wrapper_i.reg_addr[3] ),
    .B_N(\spi_wrapper_i.reg_addr[2] ),
    .Y(_0252_));
 sg13g2_and2_1 _0657_ (.A(\spi_wrapper_i.reg_addr[1] ),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .X(_0253_));
 sg13g2_and2_1 _0658_ (.A(_0252_),
    .B(_0253_),
    .X(_0254_));
 sg13g2_a22oi_1 _0659_ (.Y(_0255_),
    .B1(net277),
    .B2(\config_regs[56] ),
    .A2(_0251_),
    .A1(\config_regs[104] ));
 sg13g2_and2_1 _0660_ (.A(_0247_),
    .B(_0250_),
    .X(_0256_));
 sg13g2_and2_1 _0661_ (.A(_0243_),
    .B(_0247_),
    .X(_0257_));
 sg13g2_a22oi_1 _0662_ (.Y(_0258_),
    .B1(net275),
    .B2(\config_regs[80] ),
    .A2(net276),
    .A1(\config_regs[112] ));
 sg13g2_and2_1 _0663_ (.A(_0246_),
    .B(_0253_),
    .X(_0259_));
 sg13g2_and2_1 _0664_ (.A(_0243_),
    .B(_0253_),
    .X(_0260_));
 sg13g2_a22oi_1 _0665_ (.Y(_0261_),
    .B1(_0260_),
    .B2(\config_regs[88] ),
    .A2(net274),
    .A1(\config_regs[24] ));
 sg13g2_nand4_1 _0666_ (.B(_0255_),
    .C(_0258_),
    .A(_0249_),
    .Y(_0262_),
    .D(_0261_));
 sg13g2_and2_1 _0667_ (.A(_0244_),
    .B(_0246_),
    .X(_0263_));
 sg13g2_nand2_1 _0668_ (.Y(_0264_),
    .A(\config_regs[8] ),
    .B(net271));
 sg13g2_nor2_2 _0669_ (.A(\spi_wrapper_i.reg_addr[1] ),
    .B(\spi_wrapper_i.reg_addr[0] ),
    .Y(_0265_));
 sg13g2_and2_1 _0670_ (.A(_0243_),
    .B(_0265_),
    .X(_0266_));
 sg13g2_and2_1 _0671_ (.A(_0250_),
    .B(_0265_),
    .X(_0267_));
 sg13g2_a22oi_1 _0672_ (.Y(_0268_),
    .B1(net269),
    .B2(\config_regs[96] ),
    .A2(net270),
    .A1(\config_regs[64] ));
 sg13g2_and2_1 _0673_ (.A(_0250_),
    .B(_0253_),
    .X(_0269_));
 sg13g2_and2_1 _0674_ (.A(_0244_),
    .B(_0252_),
    .X(_0270_));
 sg13g2_a22oi_1 _0675_ (.Y(_0271_),
    .B1(net267),
    .B2(\config_regs[40] ),
    .A2(net268),
    .A1(\config_regs[120] ));
 sg13g2_nand2b_1 _0676_ (.Y(_0272_),
    .B(_0252_),
    .A_N(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_and2_1 _0677_ (.A(_0247_),
    .B(_0252_),
    .X(_0273_));
 sg13g2_and2_1 _0678_ (.A(_0252_),
    .B(_0265_),
    .X(_0274_));
 sg13g2_a22oi_1 _0679_ (.Y(_0275_),
    .B1(net264),
    .B2(\config_regs[32] ),
    .A2(net266),
    .A1(\config_regs[48] ));
 sg13g2_nand4_1 _0680_ (.B(_0268_),
    .C(_0271_),
    .A(_0264_),
    .Y(_0276_),
    .D(_0275_));
 sg13g2_and2_1 _0681_ (.A(_0246_),
    .B(_0265_),
    .X(_0277_));
 sg13g2_nand2_1 _0682_ (.Y(_0278_),
    .A(_0246_),
    .B(_0265_));
 sg13g2_o21ai_1 _0683_ (.B1(_0200_),
    .Y(_0279_),
    .A1(_0004_),
    .A2(_0278_));
 sg13g2_nor3_2 _0684_ (.A(_0262_),
    .B(_0276_),
    .C(_0279_),
    .Y(_0280_));
 sg13g2_nand3b_1 _0685_ (.B(_0272_),
    .C(net302),
    .Y(_0281_),
    .A_N(net273));
 sg13g2_nand4_1 _0686_ (.B(_0212_),
    .C(_0220_),
    .A(net336),
    .Y(_0282_),
    .D(_0281_));
 sg13g2_o21ai_1 _0687_ (.B1(_0242_),
    .Y(_0040_),
    .A1(_0280_),
    .A2(_0282_));
 sg13g2_nand2_1 _0688_ (.Y(_0283_),
    .A(net302),
    .B(_0278_));
 sg13g2_nor4_1 _0689_ (.A(net280),
    .B(net278),
    .C(net264),
    .D(_0283_),
    .Y(_0284_));
 sg13g2_nand2_1 _0690_ (.Y(_0285_),
    .A(_0006_),
    .B(net263));
 sg13g2_a22oi_1 _0691_ (.Y(_0286_),
    .B1(net271),
    .B2(\config_regs[9] ),
    .A2(net280),
    .A1(\config_regs[17] ));
 sg13g2_a22oi_1 _0692_ (.Y(_0287_),
    .B1(_0269_),
    .B2(\config_regs[121] ),
    .A2(_0256_),
    .A1(\config_regs[113] ));
 sg13g2_a21oi_1 _0693_ (.A1(\config_regs[33] ),
    .A2(net265),
    .Y(_0288_),
    .B1(net263));
 sg13g2_a22oi_1 _0694_ (.Y(_0289_),
    .B1(_0266_),
    .B2(\config_regs[65] ),
    .A2(net274),
    .A1(\config_regs[25] ));
 sg13g2_a22oi_1 _0695_ (.Y(_0290_),
    .B1(net266),
    .B2(\config_regs[49] ),
    .A2(_0267_),
    .A1(\config_regs[97] ));
 sg13g2_nand4_1 _0696_ (.B(_0288_),
    .C(_0289_),
    .A(_0286_),
    .Y(_0291_),
    .D(_0290_));
 sg13g2_a22oi_1 _0697_ (.Y(_0292_),
    .B1(net277),
    .B2(\config_regs[57] ),
    .A2(net279),
    .A1(\config_regs[105] ));
 sg13g2_a22oi_1 _0698_ (.Y(_0293_),
    .B1(net272),
    .B2(\config_regs[89] ),
    .A2(net281),
    .A1(\config_regs[73] ));
 sg13g2_a22oi_1 _0699_ (.Y(_0294_),
    .B1(net267),
    .B2(\config_regs[41] ),
    .A2(net275),
    .A1(\config_regs[81] ));
 sg13g2_nand4_1 _0700_ (.B(_0292_),
    .C(_0293_),
    .A(_0287_),
    .Y(_0295_),
    .D(_0294_));
 sg13g2_o21ai_1 _0701_ (.B1(_0285_),
    .Y(_0296_),
    .A1(_0291_),
    .A2(_0295_));
 sg13g2_a21oi_1 _0702_ (.A1(_0200_),
    .A2(_0296_),
    .Y(_0297_),
    .B1(_0284_));
 sg13g2_nand3_1 _0703_ (.B(_0212_),
    .C(_0240_),
    .A(net336),
    .Y(_0298_));
 sg13g2_a21oi_1 _0704_ (.A1(_0005_),
    .A2(net258),
    .Y(_0299_),
    .B1(_0298_));
 sg13g2_o21ai_1 _0705_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net258),
    .A2(_0297_));
 sg13g2_nand2_1 _0706_ (.Y(_0301_),
    .A(net23),
    .B(_0241_));
 sg13g2_nand2_1 _0707_ (.Y(_0041_),
    .A(_0300_),
    .B(_0301_));
 sg13g2_nand2_1 _0708_ (.Y(_0302_),
    .A(_0008_),
    .B(net263));
 sg13g2_a21oi_1 _0709_ (.A1(\config_regs[74] ),
    .A2(net281),
    .Y(_0303_),
    .B1(net263));
 sg13g2_a22oi_1 _0710_ (.Y(_0304_),
    .B1(net266),
    .B2(\config_regs[50] ),
    .A2(net267),
    .A1(\config_regs[42] ));
 sg13g2_a22oi_1 _0711_ (.Y(_0305_),
    .B1(net268),
    .B2(\config_regs[122] ),
    .A2(_0263_),
    .A1(\config_regs[10] ));
 sg13g2_a22oi_1 _0712_ (.Y(_0306_),
    .B1(net269),
    .B2(\config_regs[98] ),
    .A2(net272),
    .A1(\config_regs[90] ));
 sg13g2_nand4_1 _0713_ (.B(_0304_),
    .C(_0305_),
    .A(_0303_),
    .Y(_0307_),
    .D(_0306_));
 sg13g2_a22oi_1 _0714_ (.Y(_0308_),
    .B1(net270),
    .B2(\config_regs[66] ),
    .A2(net278),
    .A1(\config_regs[58] ));
 sg13g2_a22oi_1 _0715_ (.Y(_0309_),
    .B1(net276),
    .B2(\config_regs[114] ),
    .A2(net279),
    .A1(\config_regs[106] ));
 sg13g2_a22oi_1 _0716_ (.Y(_0310_),
    .B1(net265),
    .B2(\config_regs[34] ),
    .A2(net274),
    .A1(\config_regs[26] ));
 sg13g2_a22oi_1 _0717_ (.Y(_0311_),
    .B1(net275),
    .B2(\config_regs[82] ),
    .A2(_0248_),
    .A1(\config_regs[18] ));
 sg13g2_nand4_1 _0718_ (.B(_0309_),
    .C(_0310_),
    .A(_0308_),
    .Y(_0312_),
    .D(_0311_));
 sg13g2_o21ai_1 _0719_ (.B1(_0302_),
    .Y(_0313_),
    .A1(_0307_),
    .A2(_0312_));
 sg13g2_nand2_1 _0720_ (.Y(_0314_),
    .A(_0200_),
    .B(_0313_));
 sg13g2_a21oi_1 _0721_ (.A1(_0281_),
    .A2(_0314_),
    .Y(_0315_),
    .B1(net258));
 sg13g2_a21o_1 _0722_ (.A2(net259),
    .A1(_0007_),
    .B1(_0298_),
    .X(_0316_));
 sg13g2_nand2_1 _0723_ (.Y(_0317_),
    .A(net33),
    .B(_0241_));
 sg13g2_o21ai_1 _0724_ (.B1(_0317_),
    .Y(_0042_),
    .A1(_0315_),
    .A2(_0316_));
 sg13g2_nand2_1 _0725_ (.Y(_0318_),
    .A(_0010_),
    .B(net263));
 sg13g2_a22oi_1 _0726_ (.Y(_0319_),
    .B1(net269),
    .B2(\config_regs[99] ),
    .A2(net279),
    .A1(\config_regs[107] ));
 sg13g2_a22oi_1 _0727_ (.Y(_0320_),
    .B1(net271),
    .B2(\config_regs[11] ),
    .A2(net280),
    .A1(\config_regs[19] ));
 sg13g2_a21oi_1 _0728_ (.A1(\config_regs[35] ),
    .A2(net264),
    .Y(_0321_),
    .B1(net262));
 sg13g2_a22oi_1 _0729_ (.Y(_0322_),
    .B1(net270),
    .B2(\config_regs[67] ),
    .A2(net273),
    .A1(\config_regs[27] ));
 sg13g2_a22oi_1 _0730_ (.Y(_0323_),
    .B1(net266),
    .B2(\config_regs[51] ),
    .A2(net276),
    .A1(\config_regs[115] ));
 sg13g2_nand4_1 _0731_ (.B(_0321_),
    .C(_0322_),
    .A(_0320_),
    .Y(_0324_),
    .D(_0323_));
 sg13g2_a22oi_1 _0732_ (.Y(_0325_),
    .B1(net268),
    .B2(\config_regs[123] ),
    .A2(net277),
    .A1(\config_regs[59] ));
 sg13g2_a22oi_1 _0733_ (.Y(_0326_),
    .B1(net267),
    .B2(\config_regs[43] ),
    .A2(net275),
    .A1(\config_regs[83] ));
 sg13g2_a22oi_1 _0734_ (.Y(_0327_),
    .B1(net272),
    .B2(\config_regs[91] ),
    .A2(net281),
    .A1(\config_regs[75] ));
 sg13g2_nand4_1 _0735_ (.B(_0325_),
    .C(_0326_),
    .A(_0319_),
    .Y(_0328_),
    .D(_0327_));
 sg13g2_o21ai_1 _0736_ (.B1(_0318_),
    .Y(_0329_),
    .A1(_0324_),
    .A2(_0328_));
 sg13g2_a21oi_1 _0737_ (.A1(_0200_),
    .A2(_0329_),
    .Y(_0330_),
    .B1(_0284_));
 sg13g2_a21oi_1 _0738_ (.A1(_0009_),
    .A2(net259),
    .Y(_0331_),
    .B1(_0298_));
 sg13g2_o21ai_1 _0739_ (.B1(_0331_),
    .Y(_0332_),
    .A1(net258),
    .A2(_0330_));
 sg13g2_nand2_1 _0740_ (.Y(_0333_),
    .A(net29),
    .B(_0241_));
 sg13g2_nand2_1 _0741_ (.Y(_0043_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_a22oi_1 _0742_ (.Y(_0334_),
    .B1(net270),
    .B2(\config_regs[68] ),
    .A2(net279),
    .A1(\config_regs[108] ));
 sg13g2_a21oi_1 _0743_ (.A1(\config_regs[44] ),
    .A2(net267),
    .Y(_0335_),
    .B1(net262));
 sg13g2_a22oi_1 _0744_ (.Y(_0336_),
    .B1(net266),
    .B2(\config_regs[52] ),
    .A2(net271),
    .A1(\config_regs[12] ));
 sg13g2_a22oi_1 _0745_ (.Y(_0337_),
    .B1(net269),
    .B2(\config_regs[100] ),
    .A2(net280),
    .A1(\config_regs[20] ));
 sg13g2_nand4_1 _0746_ (.B(_0335_),
    .C(_0336_),
    .A(_0334_),
    .Y(_0338_),
    .D(_0337_));
 sg13g2_a22oi_1 _0747_ (.Y(_0339_),
    .B1(net264),
    .B2(\config_regs[36] ),
    .A2(net276),
    .A1(\config_regs[116] ));
 sg13g2_a22oi_1 _0748_ (.Y(_0340_),
    .B1(net275),
    .B2(\config_regs[84] ),
    .A2(net277),
    .A1(\config_regs[60] ));
 sg13g2_a22oi_1 _0749_ (.Y(_0341_),
    .B1(net272),
    .B2(\config_regs[92] ),
    .A2(net274),
    .A1(\config_regs[28] ));
 sg13g2_a22oi_1 _0750_ (.Y(_0342_),
    .B1(net268),
    .B2(\config_regs[124] ),
    .A2(net281),
    .A1(\config_regs[76] ));
 sg13g2_nand4_1 _0751_ (.B(_0340_),
    .C(_0341_),
    .A(_0339_),
    .Y(_0343_),
    .D(_0342_));
 sg13g2_a21oi_1 _0752_ (.A1(_0012_),
    .A2(net262),
    .Y(_0344_),
    .B1(\spi_wrapper_i.reg_addr[4] ));
 sg13g2_o21ai_1 _0753_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0338_),
    .A2(_0343_));
 sg13g2_or4_1 _0754_ (.A(net278),
    .B(net273),
    .C(net271),
    .D(net264),
    .X(_0346_));
 sg13g2_a21oi_1 _0755_ (.A1(net302),
    .A2(_0346_),
    .Y(_0347_),
    .B1(net258));
 sg13g2_a221oi_1 _0756_ (.B2(_0347_),
    .C1(_0298_),
    .B1(_0345_),
    .A1(_0011_),
    .Y(_0348_),
    .A2(net259));
 sg13g2_a21o_1 _0757_ (.A2(_0241_),
    .A1(net51),
    .B1(_0348_),
    .X(_0044_));
 sg13g2_a22oi_1 _0758_ (.Y(_0349_),
    .B1(net264),
    .B2(\config_regs[37] ),
    .A2(net272),
    .A1(\config_regs[93] ));
 sg13g2_a22oi_1 _0759_ (.Y(_0350_),
    .B1(net271),
    .B2(\config_regs[13] ),
    .A2(net273),
    .A1(\config_regs[29] ));
 sg13g2_a22oi_1 _0760_ (.Y(_0351_),
    .B1(net276),
    .B2(\config_regs[117] ),
    .A2(net279),
    .A1(\config_regs[109] ));
 sg13g2_a21oi_1 _0761_ (.A1(\config_regs[53] ),
    .A2(_0273_),
    .Y(_0352_),
    .B1(net262));
 sg13g2_a22oi_1 _0762_ (.Y(_0353_),
    .B1(net267),
    .B2(\config_regs[45] ),
    .A2(net269),
    .A1(\config_regs[101] ));
 sg13g2_nand4_1 _0763_ (.B(_0351_),
    .C(_0352_),
    .A(_0350_),
    .Y(_0354_),
    .D(_0353_));
 sg13g2_a22oi_1 _0764_ (.Y(_0355_),
    .B1(net270),
    .B2(\config_regs[69] ),
    .A2(net278),
    .A1(\config_regs[61] ));
 sg13g2_a22oi_1 _0765_ (.Y(_0356_),
    .B1(net268),
    .B2(\config_regs[125] ),
    .A2(net281),
    .A1(\config_regs[77] ));
 sg13g2_a22oi_1 _0766_ (.Y(_0357_),
    .B1(_0257_),
    .B2(\config_regs[85] ),
    .A2(net280),
    .A1(\config_regs[21] ));
 sg13g2_nand4_1 _0767_ (.B(_0355_),
    .C(_0356_),
    .A(_0349_),
    .Y(_0358_),
    .D(_0357_));
 sg13g2_a21oi_1 _0768_ (.A1(_0014_),
    .A2(net262),
    .Y(_0359_),
    .B1(net302));
 sg13g2_o21ai_1 _0769_ (.B1(_0359_),
    .Y(_0360_),
    .A1(_0354_),
    .A2(_0358_));
 sg13g2_nand2b_1 _0770_ (.Y(_0361_),
    .B(_0272_),
    .A_N(net280));
 sg13g2_a21oi_1 _0771_ (.A1(net302),
    .A2(_0361_),
    .Y(_0362_),
    .B1(_0221_));
 sg13g2_a221oi_1 _0772_ (.B2(_0362_),
    .C1(_0298_),
    .B1(_0360_),
    .A1(_0013_),
    .Y(_0363_),
    .A2(net258));
 sg13g2_a21o_1 _0773_ (.A2(_0241_),
    .A1(net93),
    .B1(_0363_),
    .X(_0045_));
 sg13g2_nand2_1 _0774_ (.Y(_0364_),
    .A(_0016_),
    .B(net262));
 sg13g2_a22oi_1 _0775_ (.Y(_0365_),
    .B1(net269),
    .B2(\config_regs[102] ),
    .A2(net279),
    .A1(\config_regs[110] ));
 sg13g2_a22oi_1 _0776_ (.Y(_0366_),
    .B1(net273),
    .B2(\config_regs[30] ),
    .A2(net280),
    .A1(\config_regs[22] ));
 sg13g2_a21oi_1 _0777_ (.A1(\config_regs[86] ),
    .A2(net275),
    .Y(_0367_),
    .B1(net263));
 sg13g2_a22oi_1 _0778_ (.Y(_0368_),
    .B1(net268),
    .B2(\config_regs[126] ),
    .A2(net281),
    .A1(\config_regs[78] ));
 sg13g2_nand4_1 _0779_ (.B(_0366_),
    .C(_0367_),
    .A(_0365_),
    .Y(_0369_),
    .D(_0368_));
 sg13g2_a22oi_1 _0780_ (.Y(_0370_),
    .B1(net270),
    .B2(\config_regs[70] ),
    .A2(net277),
    .A1(\config_regs[62] ));
 sg13g2_a22oi_1 _0781_ (.Y(_0371_),
    .B1(_0263_),
    .B2(\config_regs[14] ),
    .A2(net276),
    .A1(\config_regs[118] ));
 sg13g2_a22oi_1 _0782_ (.Y(_0372_),
    .B1(net266),
    .B2(\config_regs[54] ),
    .A2(net267),
    .A1(\config_regs[46] ));
 sg13g2_a22oi_1 _0783_ (.Y(_0373_),
    .B1(net264),
    .B2(\config_regs[38] ),
    .A2(net272),
    .A1(\config_regs[94] ));
 sg13g2_nand4_1 _0784_ (.B(_0371_),
    .C(_0372_),
    .A(_0370_),
    .Y(_0374_),
    .D(_0373_));
 sg13g2_o21ai_1 _0785_ (.B1(_0364_),
    .Y(_0375_),
    .A1(_0369_),
    .A2(_0374_));
 sg13g2_nor4_1 _0786_ (.A(net277),
    .B(net273),
    .C(net264),
    .D(_0283_),
    .Y(_0376_));
 sg13g2_a21oi_1 _0787_ (.A1(_0200_),
    .A2(_0375_),
    .Y(_0377_),
    .B1(_0376_));
 sg13g2_a21oi_1 _0788_ (.A1(_0015_),
    .A2(net258),
    .Y(_0378_),
    .B1(_0298_));
 sg13g2_o21ai_1 _0789_ (.B1(_0378_),
    .Y(_0379_),
    .A1(net258),
    .A2(_0377_));
 sg13g2_nand2_1 _0790_ (.Y(_0380_),
    .A(net25),
    .B(_0241_));
 sg13g2_nand2_1 _0791_ (.Y(_0046_),
    .A(_0379_),
    .B(_0380_));
 sg13g2_a22oi_1 _0792_ (.Y(_0381_),
    .B1(net269),
    .B2(\config_regs[103] ),
    .A2(net279),
    .A1(\config_regs[111] ));
 sg13g2_a22oi_1 _0793_ (.Y(_0382_),
    .B1(net266),
    .B2(\config_regs[55] ),
    .A2(net271),
    .A1(\config_regs[15] ));
 sg13g2_a22oi_1 _0794_ (.Y(_0383_),
    .B1(net268),
    .B2(\config_regs[127] ),
    .A2(net276),
    .A1(\config_regs[119] ));
 sg13g2_a22oi_1 _0795_ (.Y(_0384_),
    .B1(net277),
    .B2(\config_regs[63] ),
    .A2(_0248_),
    .A1(\config_regs[23] ));
 sg13g2_a21oi_1 _0796_ (.A1(\config_regs[39] ),
    .A2(net265),
    .Y(_0385_),
    .B1(net263));
 sg13g2_a22oi_1 _0797_ (.Y(_0386_),
    .B1(net270),
    .B2(\config_regs[71] ),
    .A2(net275),
    .A1(\config_regs[87] ));
 sg13g2_and4_1 _0798_ (.A(_0382_),
    .B(_0384_),
    .C(_0385_),
    .D(_0386_),
    .X(_0387_));
 sg13g2_a22oi_1 _0799_ (.Y(_0388_),
    .B1(net273),
    .B2(\config_regs[31] ),
    .A2(net281),
    .A1(\config_regs[79] ));
 sg13g2_a22oi_1 _0800_ (.Y(_0389_),
    .B1(_0270_),
    .B2(\config_regs[47] ),
    .A2(net272),
    .A1(\config_regs[95] ));
 sg13g2_and4_1 _0801_ (.A(_0381_),
    .B(_0383_),
    .C(_0388_),
    .D(_0389_),
    .X(_0390_));
 sg13g2_a22oi_1 _0802_ (.Y(_0391_),
    .B1(_0387_),
    .B2(_0390_),
    .A2(net262),
    .A1(_0018_));
 sg13g2_o21ai_1 _0803_ (.B1(net302),
    .Y(_0392_),
    .A1(\spi_wrapper_i.reg_addr[0] ),
    .A2(\spi_wrapper_i.reg_addr[3] ));
 sg13g2_o21ai_1 _0804_ (.B1(_0392_),
    .Y(_0393_),
    .A1(net302),
    .A2(_0391_));
 sg13g2_a21o_1 _0805_ (.A2(net259),
    .A1(_0017_),
    .B1(_0298_),
    .X(_0394_));
 sg13g2_a21oi_1 _0806_ (.A1(_0220_),
    .A2(_0393_),
    .Y(_0395_),
    .B1(_0394_));
 sg13g2_a21o_1 _0807_ (.A2(_0241_),
    .A1(net158),
    .B1(_0395_),
    .X(_0047_));
 sg13g2_and2_1 _0808_ (.A(net335),
    .B(\spi_wrapper_i.reg_data_o_vld ),
    .X(_0396_));
 sg13g2_and2_2 _0809_ (.A(net268),
    .B(net282),
    .X(_0397_));
 sg13g2_mux2_1 _0810_ (.A0(net46),
    .A1(net300),
    .S(_0397_),
    .X(_0048_));
 sg13g2_mux2_1 _0811_ (.A0(net77),
    .A1(net297),
    .S(_0397_),
    .X(_0049_));
 sg13g2_mux2_1 _0812_ (.A0(net142),
    .A1(net296),
    .S(_0397_),
    .X(_0050_));
 sg13g2_mux2_1 _0813_ (.A0(net64),
    .A1(net293),
    .S(_0397_),
    .X(_0051_));
 sg13g2_mux2_1 _0814_ (.A0(net112),
    .A1(net291),
    .S(_0397_),
    .X(_0052_));
 sg13g2_mux2_1 _0815_ (.A0(net154),
    .A1(net289),
    .S(_0397_),
    .X(_0053_));
 sg13g2_mux2_1 _0816_ (.A0(net147),
    .A1(net286),
    .S(_0397_),
    .X(_0054_));
 sg13g2_mux2_1 _0817_ (.A0(net176),
    .A1(net284),
    .S(_0397_),
    .X(_0055_));
 sg13g2_mux2_1 _0818_ (.A0(net38),
    .A1(net49),
    .S(net336),
    .X(_0056_));
 sg13g2_mux2_1 _0819_ (.A0(net38),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .S(net257),
    .X(_0057_));
 sg13g2_mux2_1 _0820_ (.A0(net245),
    .A1(net229),
    .S(net257),
    .X(_0058_));
 sg13g2_mux2_1 _0821_ (.A0(net229),
    .A1(net172),
    .S(net256),
    .X(_0059_));
 sg13g2_mux2_1 _0822_ (.A0(net172),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .S(net256),
    .X(_0060_));
 sg13g2_mux2_1 _0823_ (.A0(net344),
    .A1(net225),
    .S(net256),
    .X(_0061_));
 sg13g2_mux2_1 _0824_ (.A0(net225),
    .A1(net189),
    .S(net256),
    .X(_0062_));
 sg13g2_mux2_1 _0825_ (.A0(net189),
    .A1(net192),
    .S(net256),
    .X(_0063_));
 sg13g2_mux2_1 _0826_ (.A0(net192),
    .A1(net203),
    .S(net256),
    .X(_0064_));
 sg13g2_mux2_1 _0827_ (.A0(net180),
    .A1(spi_cs_n_sync),
    .S(net335),
    .X(_0065_));
 sg13g2_and2_2 _0828_ (.A(net281),
    .B(net282),
    .X(_0398_));
 sg13g2_mux2_1 _0829_ (.A0(net40),
    .A1(\spi_wrapper_i.reg_data_o[0] ),
    .S(_0398_),
    .X(_0066_));
 sg13g2_mux2_1 _0830_ (.A0(net157),
    .A1(net297),
    .S(_0398_),
    .X(_0067_));
 sg13g2_mux2_1 _0831_ (.A0(net123),
    .A1(net295),
    .S(_0398_),
    .X(_0068_));
 sg13g2_mux2_1 _0832_ (.A0(net148),
    .A1(net294),
    .S(_0398_),
    .X(_0069_));
 sg13g2_mux2_1 _0833_ (.A0(net101),
    .A1(net291),
    .S(_0398_),
    .X(_0070_));
 sg13g2_mux2_1 _0834_ (.A0(net126),
    .A1(net289),
    .S(_0398_),
    .X(_0071_));
 sg13g2_mux2_1 _0835_ (.A0(net53),
    .A1(net287),
    .S(_0398_),
    .X(_0072_));
 sg13g2_mux2_1 _0836_ (.A0(net92),
    .A1(net284),
    .S(_0398_),
    .X(_0073_));
 sg13g2_and2_2 _0837_ (.A(net269),
    .B(net283),
    .X(_0399_));
 sg13g2_mux2_1 _0838_ (.A0(net109),
    .A1(net300),
    .S(_0399_),
    .X(_0074_));
 sg13g2_mux2_1 _0839_ (.A0(net70),
    .A1(net299),
    .S(_0399_),
    .X(_0075_));
 sg13g2_mux2_1 _0840_ (.A0(net238),
    .A1(net296),
    .S(_0399_),
    .X(_0076_));
 sg13g2_mux2_1 _0841_ (.A0(net87),
    .A1(net293),
    .S(_0399_),
    .X(_0077_));
 sg13g2_mux2_1 _0842_ (.A0(net191),
    .A1(net292),
    .S(_0399_),
    .X(_0078_));
 sg13g2_mux2_1 _0843_ (.A0(net134),
    .A1(net290),
    .S(_0399_),
    .X(_0079_));
 sg13g2_mux2_1 _0844_ (.A0(net121),
    .A1(net288),
    .S(_0399_),
    .X(_0080_));
 sg13g2_mux2_1 _0845_ (.A0(net155),
    .A1(net285),
    .S(_0399_),
    .X(_0081_));
 sg13g2_nand2_2 _0846_ (.Y(_0400_),
    .A(net270),
    .B(net283));
 sg13g2_mux2_1 _0847_ (.A0(net300),
    .A1(net210),
    .S(_0400_),
    .X(_0082_));
 sg13g2_mux2_1 _0848_ (.A0(net298),
    .A1(net235),
    .S(_0400_),
    .X(_0083_));
 sg13g2_mux2_1 _0849_ (.A0(net295),
    .A1(net221),
    .S(_0400_),
    .X(_0084_));
 sg13g2_mux2_1 _0850_ (.A0(net294),
    .A1(net347),
    .S(_0400_),
    .X(_0085_));
 sg13g2_mux2_1 _0851_ (.A0(\spi_wrapper_i.reg_data_o[4] ),
    .A1(net239),
    .S(_0400_),
    .X(_0086_));
 sg13g2_mux2_1 _0852_ (.A0(\spi_wrapper_i.reg_data_o[5] ),
    .A1(net231),
    .S(_0400_),
    .X(_0087_));
 sg13g2_mux2_1 _0853_ (.A0(net287),
    .A1(net216),
    .S(_0400_),
    .X(_0088_));
 sg13g2_mux2_1 _0854_ (.A0(\spi_wrapper_i.reg_data_o[7] ),
    .A1(net251),
    .S(_0400_),
    .X(_0089_));
 sg13g2_and2_2 _0855_ (.A(net277),
    .B(net282),
    .X(_0401_));
 sg13g2_mux2_1 _0856_ (.A0(net149),
    .A1(net301),
    .S(_0401_),
    .X(_0090_));
 sg13g2_mux2_1 _0857_ (.A0(net104),
    .A1(net297),
    .S(_0401_),
    .X(_0091_));
 sg13g2_mux2_1 _0858_ (.A0(net67),
    .A1(\spi_wrapper_i.reg_data_o[2] ),
    .S(_0401_),
    .X(_0092_));
 sg13g2_mux2_1 _0859_ (.A0(net103),
    .A1(net293),
    .S(_0401_),
    .X(_0093_));
 sg13g2_mux2_1 _0860_ (.A0(net74),
    .A1(net291),
    .S(_0401_),
    .X(_0094_));
 sg13g2_mux2_1 _0861_ (.A0(net78),
    .A1(net289),
    .S(_0401_),
    .X(_0095_));
 sg13g2_mux2_1 _0862_ (.A0(net97),
    .A1(net287),
    .S(_0401_),
    .X(_0096_));
 sg13g2_mux2_1 _0863_ (.A0(net85),
    .A1(net284),
    .S(_0401_),
    .X(_0097_));
 sg13g2_and2_2 _0864_ (.A(net266),
    .B(net283),
    .X(_0402_));
 sg13g2_mux2_1 _0865_ (.A0(net166),
    .A1(net300),
    .S(_0402_),
    .X(_0098_));
 sg13g2_mux2_1 _0866_ (.A0(net164),
    .A1(net299),
    .S(_0402_),
    .X(_0099_));
 sg13g2_mux2_1 _0867_ (.A0(net83),
    .A1(net296),
    .S(_0402_),
    .X(_0100_));
 sg13g2_mux2_1 _0868_ (.A0(net167),
    .A1(net293),
    .S(_0402_),
    .X(_0101_));
 sg13g2_mux2_1 _0869_ (.A0(net169),
    .A1(net292),
    .S(_0402_),
    .X(_0102_));
 sg13g2_mux2_1 _0870_ (.A0(net254),
    .A1(net290),
    .S(_0402_),
    .X(_0103_));
 sg13g2_mux2_1 _0871_ (.A0(net130),
    .A1(net288),
    .S(_0402_),
    .X(_0104_));
 sg13g2_mux2_1 _0872_ (.A0(net152),
    .A1(net285),
    .S(_0402_),
    .X(_0105_));
 sg13g2_and2_2 _0873_ (.A(net279),
    .B(net282),
    .X(_0403_));
 sg13g2_mux2_1 _0874_ (.A0(net42),
    .A1(net301),
    .S(_0403_),
    .X(_0106_));
 sg13g2_mux2_1 _0875_ (.A0(net69),
    .A1(net297),
    .S(_0403_),
    .X(_0107_));
 sg13g2_mux2_1 _0876_ (.A0(net151),
    .A1(net295),
    .S(_0403_),
    .X(_0108_));
 sg13g2_mux2_1 _0877_ (.A0(net95),
    .A1(net293),
    .S(_0403_),
    .X(_0109_));
 sg13g2_mux2_1 _0878_ (.A0(net145),
    .A1(net292),
    .S(_0403_),
    .X(_0110_));
 sg13g2_mux2_1 _0879_ (.A0(net58),
    .A1(net290),
    .S(_0403_),
    .X(_0111_));
 sg13g2_mux2_1 _0880_ (.A0(net56),
    .A1(net288),
    .S(_0403_),
    .X(_0112_));
 sg13g2_mux2_1 _0881_ (.A0(net110),
    .A1(net285),
    .S(_0403_),
    .X(_0113_));
 sg13g2_and2_2 _0882_ (.A(net267),
    .B(net283),
    .X(_0404_));
 sg13g2_mux2_1 _0883_ (.A0(net141),
    .A1(net300),
    .S(_0404_),
    .X(_0114_));
 sg13g2_mux2_1 _0884_ (.A0(net170),
    .A1(net299),
    .S(_0404_),
    .X(_0115_));
 sg13g2_mux2_1 _0885_ (.A0(net44),
    .A1(net296),
    .S(_0404_),
    .X(_0116_));
 sg13g2_mux2_1 _0886_ (.A0(net88),
    .A1(net293),
    .S(_0404_),
    .X(_0117_));
 sg13g2_mux2_1 _0887_ (.A0(net144),
    .A1(net292),
    .S(_0404_),
    .X(_0118_));
 sg13g2_mux2_1 _0888_ (.A0(net182),
    .A1(net290),
    .S(_0404_),
    .X(_0119_));
 sg13g2_mux2_1 _0889_ (.A0(net115),
    .A1(net288),
    .S(_0404_),
    .X(_0120_));
 sg13g2_mux2_1 _0890_ (.A0(net213),
    .A1(net285),
    .S(_0404_),
    .X(_0121_));
 sg13g2_nand2_2 _0891_ (.Y(_0405_),
    .A(net265),
    .B(net283));
 sg13g2_mux2_1 _0892_ (.A0(net300),
    .A1(net244),
    .S(_0405_),
    .X(_0122_));
 sg13g2_mux2_1 _0893_ (.A0(net298),
    .A1(net247),
    .S(_0405_),
    .X(_0123_));
 sg13g2_mux2_1 _0894_ (.A0(net295),
    .A1(net246),
    .S(_0405_),
    .X(_0124_));
 sg13g2_mux2_1 _0895_ (.A0(net294),
    .A1(net209),
    .S(_0405_),
    .X(_0125_));
 sg13g2_mux2_1 _0896_ (.A0(net291),
    .A1(net227),
    .S(_0405_),
    .X(_0126_));
 sg13g2_mux2_1 _0897_ (.A0(net289),
    .A1(net241),
    .S(_0405_),
    .X(_0127_));
 sg13g2_mux2_1 _0898_ (.A0(net286),
    .A1(net233),
    .S(_0405_),
    .X(_0128_));
 sg13g2_mux2_1 _0899_ (.A0(\spi_wrapper_i.reg_data_o[7] ),
    .A1(net222),
    .S(_0405_),
    .X(_0129_));
 sg13g2_and2_2 _0900_ (.A(net273),
    .B(_0396_),
    .X(_0406_));
 sg13g2_mux2_1 _0901_ (.A0(net105),
    .A1(net301),
    .S(_0406_),
    .X(_0130_));
 sg13g2_mux2_1 _0902_ (.A0(net89),
    .A1(net298),
    .S(_0406_),
    .X(_0131_));
 sg13g2_mux2_1 _0903_ (.A0(net133),
    .A1(net295),
    .S(_0406_),
    .X(_0132_));
 sg13g2_mux2_1 _0904_ (.A0(net188),
    .A1(net294),
    .S(_0406_),
    .X(_0133_));
 sg13g2_mux2_1 _0905_ (.A0(net50),
    .A1(net291),
    .S(_0406_),
    .X(_0134_));
 sg13g2_mux2_1 _0906_ (.A0(net211),
    .A1(net289),
    .S(_0406_),
    .X(_0135_));
 sg13g2_mux2_1 _0907_ (.A0(net163),
    .A1(net286),
    .S(_0406_),
    .X(_0136_));
 sg13g2_mux2_1 _0908_ (.A0(net161),
    .A1(net284),
    .S(_0406_),
    .X(_0137_));
 sg13g2_and2_2 _0909_ (.A(net276),
    .B(net282),
    .X(_0407_));
 sg13g2_mux2_1 _0910_ (.A0(net128),
    .A1(net301),
    .S(_0407_),
    .X(_0138_));
 sg13g2_mux2_1 _0911_ (.A0(net98),
    .A1(net297),
    .S(_0407_),
    .X(_0139_));
 sg13g2_mux2_1 _0912_ (.A0(net174),
    .A1(net295),
    .S(_0407_),
    .X(_0140_));
 sg13g2_mux2_1 _0913_ (.A0(net60),
    .A1(net293),
    .S(_0407_),
    .X(_0141_));
 sg13g2_mux2_1 _0914_ (.A0(net54),
    .A1(net291),
    .S(_0407_),
    .X(_0142_));
 sg13g2_mux2_1 _0915_ (.A0(net117),
    .A1(net290),
    .S(_0407_),
    .X(_0143_));
 sg13g2_mux2_1 _0916_ (.A0(net76),
    .A1(net286),
    .S(_0407_),
    .X(_0144_));
 sg13g2_mux2_1 _0917_ (.A0(net80),
    .A1(net284),
    .S(_0407_),
    .X(_0145_));
 sg13g2_nand2_2 _0918_ (.Y(_0408_),
    .A(net280),
    .B(net282));
 sg13g2_mux2_1 _0919_ (.A0(net301),
    .A1(net217),
    .S(_0408_),
    .X(_0146_));
 sg13g2_mux2_1 _0920_ (.A0(net298),
    .A1(net219),
    .S(_0408_),
    .X(_0147_));
 sg13g2_mux2_1 _0921_ (.A0(net295),
    .A1(net196),
    .S(_0408_),
    .X(_0148_));
 sg13g2_mux2_1 _0922_ (.A0(net35),
    .A1(\config_regs[19] ),
    .S(_0408_),
    .X(_0149_));
 sg13g2_mux2_1 _0923_ (.A0(net292),
    .A1(net198),
    .S(_0408_),
    .X(_0150_));
 sg13g2_mux2_1 _0924_ (.A0(net289),
    .A1(net200),
    .S(_0408_),
    .X(_0151_));
 sg13g2_mux2_1 _0925_ (.A0(net286),
    .A1(net212),
    .S(_0408_),
    .X(_0152_));
 sg13g2_mux2_1 _0926_ (.A0(net284),
    .A1(net184),
    .S(_0408_),
    .X(_0153_));
 sg13g2_nand2_2 _0927_ (.Y(_0409_),
    .A(net271),
    .B(net283));
 sg13g2_mux2_1 _0928_ (.A0(net300),
    .A1(net234),
    .S(_0409_),
    .X(_0154_));
 sg13g2_mux2_1 _0929_ (.A0(net299),
    .A1(net340),
    .S(_0409_),
    .X(_0155_));
 sg13g2_mux2_1 _0930_ (.A0(net296),
    .A1(net226),
    .S(_0409_),
    .X(_0156_));
 sg13g2_mux2_1 _0931_ (.A0(net35),
    .A1(net162),
    .S(_0409_),
    .X(_0157_));
 sg13g2_mux2_1 _0932_ (.A0(net292),
    .A1(net204),
    .S(_0409_),
    .X(_0158_));
 sg13g2_mux2_1 _0933_ (.A0(net290),
    .A1(net236),
    .S(_0409_),
    .X(_0159_));
 sg13g2_mux2_1 _0934_ (.A0(net286),
    .A1(net243),
    .S(_0409_),
    .X(_0160_));
 sg13g2_mux2_1 _0935_ (.A0(net285),
    .A1(net205),
    .S(_0409_),
    .X(_0161_));
 sg13g2_and2_2 _0936_ (.A(net275),
    .B(net282),
    .X(_0410_));
 sg13g2_mux2_1 _0937_ (.A0(net178),
    .A1(net301),
    .S(_0410_),
    .X(_0162_));
 sg13g2_mux2_1 _0938_ (.A0(net82),
    .A1(net297),
    .S(_0410_),
    .X(_0163_));
 sg13g2_mux2_1 _0939_ (.A0(net86),
    .A1(net295),
    .S(_0410_),
    .X(_0164_));
 sg13g2_mux2_1 _0940_ (.A0(net175),
    .A1(net294),
    .S(_0410_),
    .X(_0165_));
 sg13g2_mux2_1 _0941_ (.A0(net124),
    .A1(net291),
    .S(_0410_),
    .X(_0166_));
 sg13g2_mux2_1 _0942_ (.A0(net185),
    .A1(net289),
    .S(_0410_),
    .X(_0167_));
 sg13g2_mux2_1 _0943_ (.A0(net91),
    .A1(net286),
    .S(_0410_),
    .X(_0168_));
 sg13g2_mux2_1 _0944_ (.A0(net168),
    .A1(net284),
    .S(_0410_),
    .X(_0169_));
 sg13g2_and2_2 _0945_ (.A(net262),
    .B(net283),
    .X(_0411_));
 sg13g2_mux2_1 _0946_ (.A0(net99),
    .A1(net301),
    .S(_0411_),
    .X(_0170_));
 sg13g2_mux2_1 _0947_ (.A0(net96),
    .A1(net297),
    .S(_0411_),
    .X(_0171_));
 sg13g2_mux2_1 _0948_ (.A0(net139),
    .A1(\spi_wrapper_i.reg_data_o[2] ),
    .S(_0411_),
    .X(_0172_));
 sg13g2_mux2_1 _0949_ (.A0(net132),
    .A1(net294),
    .S(_0411_),
    .X(_0173_));
 sg13g2_mux2_1 _0950_ (.A0(net63),
    .A1(net292),
    .S(_0411_),
    .X(_0174_));
 sg13g2_mux2_1 _0951_ (.A0(net61),
    .A1(net290),
    .S(_0411_),
    .X(_0175_));
 sg13g2_mux2_1 _0952_ (.A0(net119),
    .A1(net287),
    .S(_0411_),
    .X(_0176_));
 sg13g2_mux2_1 _0953_ (.A0(net65),
    .A1(net285),
    .S(_0411_),
    .X(_0177_));
 sg13g2_and2_2 _0954_ (.A(net272),
    .B(net282),
    .X(_0412_));
 sg13g2_mux2_1 _0955_ (.A0(net136),
    .A1(\spi_wrapper_i.reg_data_o[0] ),
    .S(_0412_),
    .X(_0178_));
 sg13g2_mux2_1 _0956_ (.A0(net160),
    .A1(net297),
    .S(_0412_),
    .X(_0179_));
 sg13g2_mux2_1 _0957_ (.A0(net107),
    .A1(net296),
    .S(_0412_),
    .X(_0180_));
 sg13g2_mux2_1 _0958_ (.A0(net90),
    .A1(net293),
    .S(_0412_),
    .X(_0181_));
 sg13g2_mux2_1 _0959_ (.A0(net138),
    .A1(net291),
    .S(_0412_),
    .X(_0182_));
 sg13g2_mux2_1 _0960_ (.A0(net72),
    .A1(net289),
    .S(_0412_),
    .X(_0183_));
 sg13g2_mux2_1 _0961_ (.A0(net81),
    .A1(net286),
    .S(_0412_),
    .X(_0184_));
 sg13g2_mux2_1 _0962_ (.A0(net114),
    .A1(net284),
    .S(_0412_),
    .X(_0185_));
 sg13g2_mux2_1 _0963_ (.A0(net193),
    .A1(net2),
    .S(net337),
    .X(_0186_));
 sg13g2_mux2_1 _0964_ (.A0(net208),
    .A1(net146),
    .S(net337),
    .X(_0187_));
 sg13g2_mux2_1 _0965_ (.A0(net146),
    .A1(net3),
    .S(net337),
    .X(_0188_));
 sg13g2_mux2_1 _0966_ (.A0(net215),
    .A1(net253),
    .S(net335),
    .X(_0189_));
 sg13g2_mux2_1 _0967_ (.A0(net253),
    .A1(net4),
    .S(net337),
    .X(_0190_));
 sg13g2_mux2_1 _0968_ (.A0(net187),
    .A1(net120),
    .S(net1),
    .X(_0191_));
 sg13g2_mux2_1 _0969_ (.A0(net120),
    .A1(net5),
    .S(net337),
    .X(_0192_));
 sg13g2_mux2_1 _0970_ (.A0(net202),
    .A1(net187),
    .S(net336),
    .X(_0193_));
 sg13g2_mux2_1 _0971_ (.A0(net49),
    .A1(net6),
    .S(net337),
    .X(_0194_));
 sg13g2_mux2_1 _0972_ (.A0(net194),
    .A1(net193),
    .S(net337),
    .X(_0195_));
 sg13g2_dfrbp_1 _0973_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net312),
    .D(_0020_),
    .Q_N(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .Q(_0019_));
 sg13g2_dfrbp_1 _0974_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net312),
    .D(net32),
    .Q_N(_0573_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[1] ));
 sg13g2_dfrbp_1 _0975_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net311),
    .D(net48),
    .Q_N(_0574_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_dfrbp_1 _0976_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net312),
    .D(net22),
    .Q_N(_0575_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_dfrbp_1 _0977_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net311),
    .D(_0003_),
    .Q_N(_0572_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_dfrbp_1 _0978_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net311),
    .D(_0021_),
    .Q_N(_0571_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[0] ));
 sg13g2_dfrbp_1 _0979_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net311),
    .D(net343),
    .Q_N(_0570_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ));
 sg13g2_dfrbp_1 _0980_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net311),
    .D(net250),
    .Q_N(_0569_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[2] ));
 sg13g2_dfrbp_1 _0981_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net311),
    .D(_0024_),
    .Q_N(_0568_),
    .Q(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ));
 sg13g2_dfrbp_1 _0982_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net311),
    .D(_0025_),
    .Q_N(_0567_),
    .Q(\spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_dfrbp_1 _0983_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net315),
    .D(_0026_),
    .Q_N(_0566_),
    .Q(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_dfrbp_1 _0984_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net315),
    .D(_0027_),
    .Q_N(_0565_),
    .Q(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_dfrbp_1 _0985_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net310),
    .D(_0028_),
    .Q_N(_0564_),
    .Q(\spi_wrapper_i.reg_addr[2] ));
 sg13g2_dfrbp_1 _0986_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net315),
    .D(_0029_),
    .Q_N(_0563_),
    .Q(\spi_wrapper_i.reg_addr[3] ));
 sg13g2_dfrbp_1 _0987_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net315),
    .D(_0030_),
    .Q_N(_0562_),
    .Q(\spi_wrapper_i.reg_addr[4] ));
 sg13g2_dfrbp_1 _0988_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net312),
    .D(_0031_),
    .Q_N(_0561_),
    .Q(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_dfrbp_1 _0989_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net314),
    .D(_0032_),
    .Q_N(_0560_),
    .Q(\spi_wrapper_i.reg_data_o[0] ));
 sg13g2_dfrbp_1 _0990_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net312),
    .D(net230),
    .Q_N(_0559_),
    .Q(\spi_wrapper_i.reg_data_o[1] ));
 sg13g2_dfrbp_1 _0991_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net310),
    .D(_0034_),
    .Q_N(_0558_),
    .Q(\spi_wrapper_i.reg_data_o[2] ));
 sg13g2_dfrbp_1 _0992_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net315),
    .D(_0035_),
    .Q_N(_0557_),
    .Q(\spi_wrapper_i.reg_data_o[3] ));
 sg13g2_dfrbp_1 _0993_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net310),
    .D(_0036_),
    .Q_N(_0556_),
    .Q(\spi_wrapper_i.reg_data_o[4] ));
 sg13g2_dfrbp_1 _0994_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net309),
    .D(net190),
    .Q_N(_0555_),
    .Q(\spi_wrapper_i.reg_data_o[5] ));
 sg13g2_dfrbp_1 _0995_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net309),
    .D(_0038_),
    .Q_N(_0554_),
    .Q(\spi_wrapper_i.reg_data_o[6] ));
 sg13g2_dfrbp_1 _0996_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net310),
    .D(_0039_),
    .Q_N(_0553_),
    .Q(\spi_wrapper_i.reg_data_o[7] ));
 sg13g2_dfrbp_1 _0997_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net325),
    .D(net28),
    .Q_N(_0005_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ));
 sg13g2_dfrbp_1 _0998_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net326),
    .D(net24),
    .Q_N(_0007_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ));
 sg13g2_dfrbp_1 _0999_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net326),
    .D(net34),
    .Q_N(_0009_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ));
 sg13g2_dfrbp_1 _1000_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net326),
    .D(net30),
    .Q_N(_0011_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_dfrbp_1 _1001_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net325),
    .D(net52),
    .Q_N(_0013_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_dfrbp_1 _1002_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net325),
    .D(net94),
    .Q_N(_0015_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ));
 sg13g2_dfrbp_1 _1003_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net325),
    .D(net26),
    .Q_N(_0017_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_dfrbp_1 _1004_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net314),
    .D(net159),
    .Q_N(_0552_),
    .Q(spi_miso));
 sg13g2_dfrbp_1 _1005_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net305),
    .D(_0048_),
    .Q_N(_0551_),
    .Q(\config_regs[120] ));
 sg13g2_dfrbp_1 _1006_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net317),
    .D(_0049_),
    .Q_N(_0550_),
    .Q(\config_regs[121] ));
 sg13g2_dfrbp_1 _1007_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net305),
    .D(net143),
    .Q_N(_0549_),
    .Q(\config_regs[122] ));
 sg13g2_dfrbp_1 _1008_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net321),
    .D(_0051_),
    .Q_N(_0548_),
    .Q(\config_regs[123] ));
 sg13g2_dfrbp_1 _1009_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net322),
    .D(net113),
    .Q_N(_0547_),
    .Q(\config_regs[124] ));
 sg13g2_dfrbp_1 _1010_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net322),
    .D(_0053_),
    .Q_N(_0546_),
    .Q(\config_regs[125] ));
 sg13g2_dfrbp_1 _1011_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net317),
    .D(_0054_),
    .Q_N(_0545_),
    .Q(\config_regs[126] ));
 sg13g2_dfrbp_1 _1012_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net318),
    .D(_0055_),
    .Q_N(_0544_),
    .Q(\config_regs[127] ));
 sg13g2_dfrbp_1 _1013_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net316),
    .D(_0056_),
    .Q_N(_0543_),
    .Q(spi_mosi_sync));
 sg13g2_dfrbp_1 _1014_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net314),
    .D(net39),
    .Q_N(_0542_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ));
 sg13g2_dfrbp_1 _1015_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net312),
    .D(_0058_),
    .Q_N(_0541_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ));
 sg13g2_dfrbp_1 _1016_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net310),
    .D(_0059_),
    .Q_N(_0540_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ));
 sg13g2_dfrbp_1 _1017_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net309),
    .D(net173),
    .Q_N(_0539_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ));
 sg13g2_dfrbp_1 _1018_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net309),
    .D(_0061_),
    .Q_N(_0538_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ));
 sg13g2_dfrbp_1 _1019_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net309),
    .D(_0062_),
    .Q_N(_0537_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ));
 sg13g2_dfrbp_1 _1020_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net309),
    .D(_0063_),
    .Q_N(_0536_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ));
 sg13g2_dfrbp_1 _1021_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net309),
    .D(_0064_),
    .Q_N(_0535_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ));
 sg13g2_dfrbp_1 _1022_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net311),
    .D(net181),
    .Q_N(_0534_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_dfrbp_1 _1023_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net323),
    .D(net41),
    .Q_N(_0533_),
    .Q(\config_regs[72] ));
 sg13g2_dfrbp_1 _1024_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net321),
    .D(_0067_),
    .Q_N(_0532_),
    .Q(\config_regs[73] ));
 sg13g2_dfrbp_1 _1025_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net318),
    .D(_0068_),
    .Q_N(_0531_),
    .Q(\config_regs[74] ));
 sg13g2_dfrbp_1 _1026_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net317),
    .D(_0069_),
    .Q_N(_0530_),
    .Q(\config_regs[75] ));
 sg13g2_dfrbp_1 _1027_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net322),
    .D(net102),
    .Q_N(_0529_),
    .Q(\config_regs[76] ));
 sg13g2_dfrbp_1 _1028_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net322),
    .D(net127),
    .Q_N(_0528_),
    .Q(\config_regs[77] ));
 sg13g2_dfrbp_1 _1029_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net317),
    .D(_0072_),
    .Q_N(_0527_),
    .Q(\config_regs[78] ));
 sg13g2_dfrbp_1 _1030_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net317),
    .D(_0073_),
    .Q_N(_0526_),
    .Q(\config_regs[79] ));
 sg13g2_dfrbp_1 _1031_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net306),
    .D(_0074_),
    .Q_N(_0525_),
    .Q(\config_regs[96] ));
 sg13g2_dfrbp_1 _1032_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net303),
    .D(net71),
    .Q_N(_0524_),
    .Q(\config_regs[97] ));
 sg13g2_dfrbp_1 _1033_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net304),
    .D(_0076_),
    .Q_N(_0523_),
    .Q(\config_regs[98] ));
 sg13g2_dfrbp_1 _1034_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net304),
    .D(_0077_),
    .Q_N(_0522_),
    .Q(\config_regs[99] ));
 sg13g2_dfrbp_1 _1035_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net306),
    .D(_0078_),
    .Q_N(_0521_),
    .Q(\config_regs[100] ));
 sg13g2_dfrbp_1 _1036_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net303),
    .D(net135),
    .Q_N(_0520_),
    .Q(\config_regs[101] ));
 sg13g2_dfrbp_1 _1037_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net304),
    .D(net122),
    .Q_N(_0519_),
    .Q(\config_regs[102] ));
 sg13g2_dfrbp_1 _1038_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net304),
    .D(net156),
    .Q_N(_0518_),
    .Q(\config_regs[103] ));
 sg13g2_dfrbp_1 _1039_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net319),
    .D(_0082_),
    .Q_N(_0517_),
    .Q(\config_regs[64] ));
 sg13g2_dfrbp_1 _1040_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net330),
    .D(_0083_),
    .Q_N(_0516_),
    .Q(\config_regs[65] ));
 sg13g2_dfrbp_1 _1041_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net328),
    .D(_0084_),
    .Q_N(_0515_),
    .Q(\config_regs[66] ));
 sg13g2_dfrbp_1 _1042_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net330),
    .D(_0085_),
    .Q_N(_0514_),
    .Q(\config_regs[67] ));
 sg13g2_dfrbp_1 _1043_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net319),
    .D(net240),
    .Q_N(_0513_),
    .Q(\config_regs[68] ));
 sg13g2_dfrbp_1 _1044_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net329),
    .D(net232),
    .Q_N(_0512_),
    .Q(\config_regs[69] ));
 sg13g2_dfrbp_1 _1045_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net327),
    .D(_0088_),
    .Q_N(_0511_),
    .Q(\config_regs[70] ));
 sg13g2_dfrbp_1 _1046_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net328),
    .D(net252),
    .Q_N(_0510_),
    .Q(\config_regs[71] ));
 sg13g2_dfrbp_1 _1047_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net321),
    .D(net150),
    .Q_N(_0509_),
    .Q(\config_regs[56] ));
 sg13g2_dfrbp_1 _1048_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net321),
    .D(_0091_),
    .Q_N(_0508_),
    .Q(\config_regs[57] ));
 sg13g2_dfrbp_1 _1049_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net329),
    .D(net68),
    .Q_N(_0507_),
    .Q(\config_regs[58] ));
 sg13g2_dfrbp_1 _1050_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net321),
    .D(_0093_),
    .Q_N(_0506_),
    .Q(\config_regs[59] ));
 sg13g2_dfrbp_1 _1051_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net322),
    .D(net75),
    .Q_N(_0505_),
    .Q(\config_regs[60] ));
 sg13g2_dfrbp_1 _1052_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net329),
    .D(net79),
    .Q_N(_0504_),
    .Q(\config_regs[61] ));
 sg13g2_dfrbp_1 _1053_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net328),
    .D(_0096_),
    .Q_N(_0503_),
    .Q(\config_regs[62] ));
 sg13g2_dfrbp_1 _1054_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net328),
    .D(_0097_),
    .Q_N(_0502_),
    .Q(\config_regs[63] ));
 sg13g2_dfrbp_1 _1055_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net306),
    .D(_0098_),
    .Q_N(_0501_),
    .Q(\config_regs[48] ));
 sg13g2_dfrbp_1 _1056_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net303),
    .D(net165),
    .Q_N(_0500_),
    .Q(\config_regs[49] ));
 sg13g2_dfrbp_1 _1057_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net308),
    .D(net84),
    .Q_N(_0499_),
    .Q(\config_regs[50] ));
 sg13g2_dfrbp_1 _1058_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net306),
    .D(_0101_),
    .Q_N(_0498_),
    .Q(\config_regs[51] ));
 sg13g2_dfrbp_1 _1059_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net303),
    .D(_0102_),
    .Q_N(_0497_),
    .Q(\config_regs[52] ));
 sg13g2_dfrbp_1 _1060_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net303),
    .D(net255),
    .Q_N(_0496_),
    .Q(\config_regs[53] ));
 sg13g2_dfrbp_1 _1061_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net303),
    .D(net131),
    .Q_N(_0495_),
    .Q(\config_regs[54] ));
 sg13g2_dfrbp_1 _1062_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net309),
    .D(net153),
    .Q_N(_0494_),
    .Q(\config_regs[55] ));
 sg13g2_dfrbp_1 _1063_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net322),
    .D(net43),
    .Q_N(_0493_),
    .Q(\config_regs[104] ));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net317),
    .D(_0107_),
    .Q_N(_0492_),
    .Q(\config_regs[105] ));
 sg13g2_dfrbp_1 _1065_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net324),
    .D(_0108_),
    .Q_N(_0491_),
    .Q(\config_regs[106] ));
 sg13g2_dfrbp_1 _1066_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net304),
    .D(_0109_),
    .Q_N(_0490_),
    .Q(\config_regs[107] ));
 sg13g2_dfrbp_1 _1067_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net319),
    .D(_0110_),
    .Q_N(_0489_),
    .Q(\config_regs[108] ));
 sg13g2_dfrbp_1 _1068_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net305),
    .D(net59),
    .Q_N(_0488_),
    .Q(\config_regs[109] ));
 sg13g2_dfrbp_1 _1069_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net305),
    .D(net57),
    .Q_N(_0487_),
    .Q(\config_regs[110] ));
 sg13g2_dfrbp_1 _1070_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net304),
    .D(net111),
    .Q_N(_0486_),
    .Q(\config_regs[111] ));
 sg13g2_dfrbp_1 _1071_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net304),
    .D(_0114_),
    .Q_N(_0485_),
    .Q(\config_regs[40] ));
 sg13g2_dfrbp_1 _1072_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net307),
    .D(net171),
    .Q_N(_0484_),
    .Q(\config_regs[41] ));
 sg13g2_dfrbp_1 _1073_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net303),
    .D(net45),
    .Q_N(_0483_),
    .Q(\config_regs[42] ));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net307),
    .D(_0117_),
    .Q_N(_0482_),
    .Q(\config_regs[43] ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net306),
    .D(_0118_),
    .Q_N(_0481_),
    .Q(\config_regs[44] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net303),
    .D(net183),
    .Q_N(_0480_),
    .Q(\config_regs[45] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net308),
    .D(net116),
    .Q_N(_0479_),
    .Q(\config_regs[46] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net304),
    .D(net214),
    .Q_N(_0478_),
    .Q(\config_regs[47] ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net327),
    .D(_0122_),
    .Q_N(_0477_),
    .Q(\config_regs[32] ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net327),
    .D(_0123_),
    .Q_N(_0476_),
    .Q(\config_regs[33] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net331),
    .D(_0124_),
    .Q_N(_0475_),
    .Q(\config_regs[34] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net327),
    .D(_0125_),
    .Q_N(_0474_),
    .Q(\config_regs[35] ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net324),
    .D(net228),
    .Q_N(_0473_),
    .Q(\config_regs[36] ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net324),
    .D(net242),
    .Q_N(_0472_),
    .Q(\config_regs[37] ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net320),
    .D(_0128_),
    .Q_N(_0471_),
    .Q(\config_regs[38] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net328),
    .D(net223),
    .Q_N(_0470_),
    .Q(\config_regs[39] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net323),
    .D(net106),
    .Q_N(_0469_),
    .Q(\config_regs[24] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net330),
    .D(_0131_),
    .Q_N(_0468_),
    .Q(\config_regs[25] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net331),
    .D(_0132_),
    .Q_N(_0467_),
    .Q(\config_regs[26] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net330),
    .D(_0133_),
    .Q_N(_0466_),
    .Q(\config_regs[27] ));
 sg13g2_dfrbp_1 _1091_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net323),
    .D(_0134_),
    .Q_N(_0465_),
    .Q(\config_regs[28] ));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net320),
    .D(_0135_),
    .Q_N(_0464_),
    .Q(\config_regs[29] ));
 sg13g2_dfrbp_1 _1093_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net319),
    .D(_0136_),
    .Q_N(_0463_),
    .Q(\config_regs[30] ));
 sg13g2_dfrbp_1 _1094_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net318),
    .D(_0137_),
    .Q_N(_0462_),
    .Q(\config_regs[31] ));
 sg13g2_dfrbp_1 _1095_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net321),
    .D(net129),
    .Q_N(_0461_),
    .Q(\config_regs[112] ));
 sg13g2_dfrbp_1 _1096_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net317),
    .D(_0139_),
    .Q_N(_0460_),
    .Q(\config_regs[113] ));
 sg13g2_dfrbp_1 _1097_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net324),
    .D(_0140_),
    .Q_N(_0459_),
    .Q(\config_regs[114] ));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net306),
    .D(_0141_),
    .Q_N(_0458_),
    .Q(\config_regs[115] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net324),
    .D(net55),
    .Q_N(_0457_),
    .Q(\config_regs[116] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net305),
    .D(net118),
    .Q_N(_0456_),
    .Q(\config_regs[117] ));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net319),
    .D(_0144_),
    .Q_N(_0455_),
    .Q(\config_regs[118] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net318),
    .D(_0145_),
    .Q_N(_0454_),
    .Q(\config_regs[119] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net324),
    .D(net218),
    .Q_N(_0453_),
    .Q(\config_regs[16] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net327),
    .D(net220),
    .Q_N(_0452_),
    .Q(\config_regs[17] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net328),
    .D(_0148_),
    .Q_N(_0451_),
    .Q(\config_regs[18] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net327),
    .D(net36),
    .Q_N(_0450_),
    .Q(\config_regs[19] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net319),
    .D(net199),
    .Q_N(_0449_),
    .Q(\config_regs[20] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net323),
    .D(net201),
    .Q_N(_0448_),
    .Q(\config_regs[21] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net320),
    .D(_0152_),
    .Q_N(_0447_),
    .Q(\config_regs[22] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net328),
    .D(_0153_),
    .Q_N(_0446_),
    .Q(\config_regs[23] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net307),
    .D(_0154_),
    .Q_N(_0445_),
    .Q(\config_regs[8] ));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net315),
    .D(net341),
    .Q_N(_0444_),
    .Q(\config_regs[9] ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net306),
    .D(_0156_),
    .Q_N(_0443_),
    .Q(\config_regs[10] ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net315),
    .D(_0157_),
    .Q_N(_0442_),
    .Q(\config_regs[11] ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net306),
    .D(_0158_),
    .Q_N(_0441_),
    .Q(\config_regs[12] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net307),
    .D(net237),
    .Q_N(_0440_),
    .Q(\config_regs[13] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net307),
    .D(_0160_),
    .Q_N(_0439_),
    .Q(\config_regs[14] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net315),
    .D(net206),
    .Q_N(_0438_),
    .Q(\config_regs[15] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net321),
    .D(net179),
    .Q_N(_0437_),
    .Q(\config_regs[80] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net318),
    .D(_0163_),
    .Q_N(_0436_),
    .Q(\config_regs[81] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net329),
    .D(_0164_),
    .Q_N(_0435_),
    .Q(\config_regs[82] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net318),
    .D(_0165_),
    .Q_N(_0434_),
    .Q(\config_regs[83] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net322),
    .D(net125),
    .Q_N(_0433_),
    .Q(\config_regs[84] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net323),
    .D(net186),
    .Q_N(_0432_),
    .Q(\config_regs[85] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net319),
    .D(_0168_),
    .Q_N(_0431_),
    .Q(\config_regs[86] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net328),
    .D(_0169_),
    .Q_N(_0430_),
    .Q(\config_regs[87] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net325),
    .D(net100),
    .Q_N(_0004_),
    .Q(\config_regs[0] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net325),
    .D(_0171_),
    .Q_N(_0006_),
    .Q(\config_regs[1] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net325),
    .D(net140),
    .Q_N(_0008_),
    .Q(\config_regs[2] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net325),
    .D(_0173_),
    .Q_N(_0010_),
    .Q(\config_regs[3] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net314),
    .D(_0174_),
    .Q_N(_0012_),
    .Q(\config_regs[4] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net314),
    .D(net62),
    .Q_N(_0014_),
    .Q(\config_regs[5] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net314),
    .D(_0176_),
    .Q_N(_0016_),
    .Q(\config_regs[6] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net316),
    .D(net66),
    .Q_N(_0018_),
    .Q(\config_regs[7] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net323),
    .D(net137),
    .Q_N(_0429_),
    .Q(\config_regs[88] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net321),
    .D(_0179_),
    .Q_N(_0428_),
    .Q(\config_regs[89] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net305),
    .D(net108),
    .Q_N(_0427_),
    .Q(\config_regs[90] ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net317),
    .D(_0181_),
    .Q_N(_0426_),
    .Q(\config_regs[91] ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net323),
    .D(_0182_),
    .Q_N(_0425_),
    .Q(\config_regs[92] ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net323),
    .D(net73),
    .Q_N(_0424_),
    .Q(\config_regs[93] ));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net319),
    .D(_0184_),
    .Q_N(_0423_),
    .Q(\config_regs[94] ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net305),
    .D(_0185_),
    .Q_N(_0422_),
    .Q(\config_regs[95] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net331),
    .D(_0186_),
    .Q_N(_0421_),
    .Q(\synchronizer_spi_mode_cpol.data_sync[1] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net331),
    .D(_0187_),
    .Q_N(_0420_),
    .Q(cpha_sync));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net330),
    .D(_0188_),
    .Q_N(_0419_),
    .Q(\synchronizer_spi_mode_cpha.data_sync[1] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net314),
    .D(_0189_),
    .Q_N(uio_oe[3]),
    .Q(spi_cs_n_sync));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net326),
    .D(_0190_),
    .Q_N(_0418_),
    .Q(\synchronizer_spi_cs_n_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net330),
    .D(_0191_),
    .Q_N(_0417_),
    .Q(spi_clk_sync));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net330),
    .D(_0192_),
    .Q_N(_0416_),
    .Q(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net314),
    .D(_0193_),
    .Q_N(_0415_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net326),
    .D(_0194_),
    .Q_N(_0414_),
    .Q(\synchronizer_spi_mosi_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net330),
    .D(_0195_),
    .Q_N(_0413_),
    .Q(cpol_sync));
 sg13g2_tielo tt_um_calonso88_spi_test_8 (.L_LO(net8));
 sg13g2_tielo tt_um_calonso88_spi_test_9 (.L_LO(net9));
 sg13g2_tielo tt_um_calonso88_spi_test_10 (.L_LO(net10));
 sg13g2_tielo tt_um_calonso88_spi_test_11 (.L_LO(net11));
 sg13g2_tielo tt_um_calonso88_spi_test_12 (.L_LO(net12));
 sg13g2_tielo tt_um_calonso88_spi_test_13 (.L_LO(net13));
 sg13g2_tielo tt_um_calonso88_spi_test_14 (.L_LO(net14));
 sg13g2_tielo tt_um_calonso88_spi_test_15 (.L_LO(net15));
 sg13g2_tielo tt_um_calonso88_spi_test_16 (.L_LO(net16));
 sg13g2_tielo tt_um_calonso88_spi_test_17 (.L_LO(net17));
 sg13g2_tielo tt_um_calonso88_spi_test_18 (.L_LO(net18));
 sg13g2_tielo tt_um_calonso88_spi_test_19 (.L_LO(net19));
 sg13g2_tielo tt_um_calonso88_spi_test_20 (.L_LO(net20));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1167_ (.A(spi_miso),
    .X(uio_out[3]));
 sg13g2_buf_1 _1168_ (.A(\config_regs[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1169_ (.A(\config_regs[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1170_ (.A(\config_regs[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _1171_ (.A(\config_regs[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1172_ (.A(\config_regs[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _1173_ (.A(\config_regs[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _1174_ (.A(\config_regs[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _1175_ (.A(\config_regs[7] ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(net257));
 sg13g2_buf_2 fanout257 (.A(_0228_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net259),
    .X(net258));
 sg13g2_buf_1 fanout259 (.A(_0221_),
    .X(net259));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(_0215_));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_0210_));
 sg13g2_buf_2 fanout262 (.A(_0277_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_0277_),
    .X(net263));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_0274_));
 sg13g2_buf_2 fanout265 (.A(_0274_),
    .X(net265));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_0273_));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_0270_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_0269_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_0267_));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_0266_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_0263_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_0260_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_0259_));
 sg13g2_buf_2 fanout274 (.A(_0259_),
    .X(net274));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_0257_));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_0256_));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_0254_));
 sg13g2_buf_2 fanout278 (.A(_0254_),
    .X(net278));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_0251_));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(_0248_));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(_0245_));
 sg13g2_buf_2 fanout282 (.A(net283),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_0396_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(net285));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(net338));
 sg13g2_buf_2 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net197),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(\spi_wrapper_i.reg_data_o[5] ),
    .X(net289));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(\spi_wrapper_i.reg_data_o[5] ));
 sg13g2_buf_2 fanout291 (.A(\spi_wrapper_i.reg_data_o[4] ),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(\spi_wrapper_i.reg_data_o[4] ),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(net294));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(net35));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(net296));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(net195));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(net299));
 sg13g2_buf_1 fanout298 (.A(net299),
    .X(net298));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(\spi_wrapper_i.reg_data_o[1] ));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(\spi_wrapper_i.reg_data_o[0] ));
 sg13g2_buf_2 fanout302 (.A(net345),
    .X(net302));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(net308));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(net305));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(net307));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(net307));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(net308));
 sg13g2_buf_2 fanout308 (.A(rst_n),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net313));
 sg13g2_buf_2 fanout310 (.A(net313),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(net313));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(net313));
 sg13g2_buf_2 fanout313 (.A(net316),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(net316));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(net316));
 sg13g2_buf_2 fanout316 (.A(rst_n),
    .X(net316));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(net318));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(net320));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(net320));
 sg13g2_buf_2 fanout320 (.A(net333),
    .X(net320));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(net322));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net333));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(net324));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(net333));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(net327));
 sg13g2_buf_2 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(net333));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(net332));
 sg13g2_buf_2 fanout329 (.A(net332),
    .X(net329));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(net332));
 sg13g2_buf_2 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_1 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(rst_n));
 sg13g2_buf_2 fanout334 (.A(net336),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net337),
    .X(net336));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(net1));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[6]),
    .X(net6));
 sg13g2_tielo tt_um_calonso88_spi_test_7 (.L_LO(net7));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0002_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold3 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0041_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold5 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0046_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold7 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0040_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold9 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0043_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold11 (.A(\spi_wrapper_i.spi_reg_inst.reg_rw ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0000_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold13 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0042_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold15 (.A(\spi_wrapper_i.reg_data_o[3] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0149_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold17 (.A(\spi_wrapper_i.reg_data_o_vld ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold18 (.A(spi_mosi_sync),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0057_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold20 (.A(\config_regs[72] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0066_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold22 (.A(\config_regs[104] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0106_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold24 (.A(\config_regs[42] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0116_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold26 (.A(\config_regs[120] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold27 (.A(\spi_wrapper_i.spi_reg_inst.state[2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0001_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold29 (.A(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold30 (.A(\config_regs[28] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold31 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0044_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold33 (.A(\config_regs[78] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold34 (.A(\config_regs[116] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0142_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold36 (.A(\config_regs[110] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0112_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold38 (.A(\config_regs[109] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0111_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold40 (.A(\config_regs[115] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold41 (.A(\config_regs[5] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0175_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold43 (.A(\config_regs[4] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold44 (.A(\config_regs[123] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold45 (.A(\config_regs[7] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0177_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold47 (.A(\config_regs[58] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0092_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold49 (.A(\config_regs[105] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold50 (.A(\config_regs[97] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0075_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold52 (.A(\config_regs[93] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0183_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold54 (.A(\config_regs[60] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0094_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold56 (.A(\config_regs[118] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold57 (.A(\config_regs[121] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold58 (.A(\config_regs[61] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0095_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold60 (.A(\config_regs[119] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold61 (.A(\config_regs[94] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold62 (.A(\config_regs[81] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold63 (.A(\config_regs[50] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0100_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold65 (.A(\config_regs[63] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold66 (.A(\config_regs[82] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold67 (.A(\config_regs[99] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold68 (.A(\config_regs[43] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold69 (.A(\config_regs[25] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold70 (.A(\config_regs[91] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold71 (.A(\config_regs[86] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold72 (.A(\config_regs[79] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold73 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0045_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold75 (.A(\config_regs[107] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold76 (.A(\config_regs[1] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold77 (.A(\config_regs[62] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold78 (.A(\config_regs[113] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold79 (.A(\config_regs[0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0170_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold81 (.A(\config_regs[76] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0070_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold83 (.A(\config_regs[59] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold84 (.A(\config_regs[57] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold85 (.A(\config_regs[24] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0130_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold87 (.A(\config_regs[90] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0180_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold89 (.A(\config_regs[96] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold90 (.A(\config_regs[111] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0113_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold92 (.A(\config_regs[124] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0052_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold94 (.A(\config_regs[95] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold95 (.A(\config_regs[46] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0120_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold97 (.A(\config_regs[117] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0143_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold99 (.A(\config_regs[6] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold100 (.A(\synchronizer_spi_clk_inst.data_sync[1] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold101 (.A(\config_regs[102] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0080_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold103 (.A(\config_regs[74] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold104 (.A(\config_regs[84] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0166_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold106 (.A(\config_regs[77] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0071_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold108 (.A(\config_regs[112] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0138_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold110 (.A(\config_regs[54] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0104_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold112 (.A(\config_regs[3] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold113 (.A(\config_regs[26] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold114 (.A(\config_regs[101] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0079_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold116 (.A(\config_regs[88] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0178_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold118 (.A(\config_regs[92] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold119 (.A(\config_regs[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0172_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold121 (.A(\config_regs[40] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold122 (.A(\config_regs[122] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0050_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold124 (.A(\config_regs[44] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold125 (.A(\config_regs[108] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold126 (.A(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold127 (.A(\config_regs[126] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold128 (.A(\config_regs[75] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold129 (.A(\config_regs[56] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0090_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold131 (.A(\config_regs[106] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold132 (.A(\config_regs[55] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0105_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold134 (.A(\config_regs[125] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold135 (.A(\config_regs[103] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0081_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold137 (.A(\config_regs[73] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold138 (.A(spi_miso),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0047_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold140 (.A(\config_regs[89] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold141 (.A(\config_regs[31] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold142 (.A(\config_regs[11] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold143 (.A(\config_regs[30] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold144 (.A(\config_regs[49] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0099_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold146 (.A(\config_regs[48] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold147 (.A(\config_regs[51] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold148 (.A(\config_regs[87] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold149 (.A(\config_regs[52] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold150 (.A(\config_regs[41] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0115_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold152 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0060_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold154 (.A(\config_regs[114] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold155 (.A(\config_regs[83] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold156 (.A(\config_regs[127] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold157 (.A(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold158 (.A(\config_regs[80] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0162_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold160 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0065_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold162 (.A(\config_regs[45] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0119_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold164 (.A(\config_regs[23] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold165 (.A(\config_regs[85] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0167_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold167 (.A(spi_clk_sync),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold168 (.A(\config_regs[27] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold169 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0037_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold171 (.A(\config_regs[100] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold172 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold173 (.A(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold174 (.A(cpol_sync),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold175 (.A(\spi_wrapper_i.reg_data_o[2] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold176 (.A(\config_regs[18] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold177 (.A(\spi_wrapper_i.reg_data_o[6] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold178 (.A(\config_regs[20] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0150_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold180 (.A(\config_regs[21] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0151_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold182 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold183 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold184 (.A(\config_regs[12] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold185 (.A(\config_regs[15] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0161_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold187 (.A(\spi_wrapper_i.reg_addr[2] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold188 (.A(cpha_sync),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold189 (.A(\config_regs[35] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold190 (.A(\config_regs[64] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold191 (.A(\config_regs[29] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold192 (.A(\config_regs[22] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold193 (.A(\config_regs[47] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0121_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold195 (.A(spi_cs_n_sync),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold196 (.A(\config_regs[70] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold197 (.A(\config_regs[16] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0146_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold199 (.A(\config_regs[17] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0147_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold201 (.A(\config_regs[66] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold202 (.A(\config_regs[39] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0129_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold204 (.A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold205 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold206 (.A(\config_regs[10] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold207 (.A(\config_regs[36] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0126_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold209 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0033_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold211 (.A(\config_regs[69] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0087_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold213 (.A(\config_regs[38] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold214 (.A(\config_regs[8] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold215 (.A(\config_regs[65] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold216 (.A(\config_regs[13] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0159_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold218 (.A(\config_regs[98] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold219 (.A(\config_regs[68] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0086_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold221 (.A(\config_regs[37] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0127_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold223 (.A(\config_regs[14] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold224 (.A(\config_regs[32] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold225 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold226 (.A(\config_regs[34] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold227 (.A(\config_regs[33] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold228 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[2] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0231_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0023_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold231 (.A(\config_regs[71] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0089_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold233 (.A(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold234 (.A(\config_regs[53] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0103_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold236 (.A(\spi_wrapper_i.reg_data_o[7] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold237 (.A(\spi_wrapper_i.reg_addr[1] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold238 (.A(\config_regs[9] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0155_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold240 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0022_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold242 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold243 (.A(\spi_wrapper_i.reg_addr[4] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold244 (.A(\spi_wrapper_i.reg_addr[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold245 (.A(\config_regs[67] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold246 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[3] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold247 (.A(\spi_wrapper_i.spi_reg_inst.buffer_counter[0] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold248 (.A(\spi_wrapper_i.reg_addr[0] ),
    .X(net350));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_4 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_4 FILLER_5_277 ();
 sg13g2_fill_1 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_8 FILLER_6_149 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_fill_1 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_4 FILLER_6_218 ();
 sg13g2_fill_2 FILLER_6_222 ();
 sg13g2_decap_8 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_fill_2 FILLER_7_70 ();
 sg13g2_fill_1 FILLER_7_72 ();
 sg13g2_decap_8 FILLER_7_82 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_decap_8 FILLER_7_106 ();
 sg13g2_fill_2 FILLER_7_113 ();
 sg13g2_decap_8 FILLER_7_149 ();
 sg13g2_decap_8 FILLER_7_156 ();
 sg13g2_decap_4 FILLER_7_163 ();
 sg13g2_fill_1 FILLER_7_167 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_211 ();
 sg13g2_fill_2 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_decap_4 FILLER_7_345 ();
 sg13g2_fill_1 FILLER_7_349 ();
 sg13g2_decap_8 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_4 FILLER_8_70 ();
 sg13g2_decap_4 FILLER_8_119 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_fill_2 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_194 ();
 sg13g2_decap_8 FILLER_8_204 ();
 sg13g2_decap_8 FILLER_8_211 ();
 sg13g2_decap_4 FILLER_8_228 ();
 sg13g2_fill_2 FILLER_8_267 ();
 sg13g2_fill_1 FILLER_8_269 ();
 sg13g2_fill_2 FILLER_8_280 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_309 ();
 sg13g2_fill_1 FILLER_8_311 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_fill_1 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_fill_1 FILLER_9_115 ();
 sg13g2_decap_4 FILLER_9_188 ();
 sg13g2_fill_1 FILLER_9_192 ();
 sg13g2_fill_2 FILLER_9_202 ();
 sg13g2_decap_8 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_245 ();
 sg13g2_fill_1 FILLER_9_256 ();
 sg13g2_fill_2 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_49 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_fill_2 FILLER_10_157 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_decap_4 FILLER_10_226 ();
 sg13g2_fill_1 FILLER_10_230 ();
 sg13g2_fill_2 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_4 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_46 ();
 sg13g2_decap_4 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_60 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_98 ();
 sg13g2_decap_4 FILLER_11_122 ();
 sg13g2_fill_1 FILLER_11_135 ();
 sg13g2_fill_1 FILLER_11_187 ();
 sg13g2_decap_4 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_decap_8 FILLER_11_258 ();
 sg13g2_fill_1 FILLER_11_265 ();
 sg13g2_fill_2 FILLER_11_307 ();
 sg13g2_fill_1 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_35 ();
 sg13g2_fill_2 FILLER_12_46 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_4 FILLER_12_235 ();
 sg13g2_fill_2 FILLER_12_239 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_4 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_18 ();
 sg13g2_decap_4 FILLER_13_55 ();
 sg13g2_decap_4 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_100 ();
 sg13g2_decap_4 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_189 ();
 sg13g2_decap_4 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_216 ();
 sg13g2_fill_1 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_4 FILLER_13_280 ();
 sg13g2_fill_1 FILLER_13_284 ();
 sg13g2_fill_2 FILLER_13_307 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_64 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_decap_4 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_decap_4 FILLER_14_188 ();
 sg13g2_decap_4 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_309 ();
 sg13g2_fill_1 FILLER_14_316 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_fill_1 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_114 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_decap_4 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_347 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_24 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_fill_1 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_80 ();
 sg13g2_fill_2 FILLER_16_107 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_decap_4 FILLER_16_136 ();
 sg13g2_decap_4 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_273 ();
 sg13g2_decap_4 FILLER_16_315 ();
 sg13g2_fill_1 FILLER_16_319 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_decap_4 FILLER_16_356 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_86 ();
 sg13g2_decap_4 FILLER_17_127 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_232 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_4 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_53 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_fill_1 FILLER_18_141 ();
 sg13g2_fill_1 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_decap_4 FILLER_18_235 ();
 sg13g2_decap_4 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_279 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_4 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_11 ();
 sg13g2_fill_1 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_decap_4 FILLER_19_172 ();
 sg13g2_decap_4 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_309 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_2 FILLER_19_360 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_54 ();
 sg13g2_fill_2 FILLER_20_73 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_decap_8 FILLER_20_127 ();
 sg13g2_decap_8 FILLER_20_134 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_decap_4 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_decap_8 FILLER_20_213 ();
 sg13g2_decap_4 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_decap_4 FILLER_20_247 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_decap_4 FILLER_20_349 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_80 ();
 sg13g2_fill_1 FILLER_21_87 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_fill_2 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_decap_4 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_76 ();
 sg13g2_decap_8 FILLER_22_83 ();
 sg13g2_fill_2 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_112 ();
 sg13g2_decap_4 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_decap_4 FILLER_22_241 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_decap_4 FILLER_22_261 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_2 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_4 FILLER_23_62 ();
 sg13g2_fill_2 FILLER_23_66 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_decap_8 FILLER_23_85 ();
 sg13g2_decap_4 FILLER_23_92 ();
 sg13g2_fill_1 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_127 ();
 sg13g2_decap_4 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_decap_8 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_4 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_fill_2 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_decap_4 FILLER_23_229 ();
 sg13g2_decap_4 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_259 ();
 sg13g2_decap_4 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_49 ();
 sg13g2_decap_4 FILLER_24_97 ();
 sg13g2_decap_8 FILLER_24_141 ();
 sg13g2_decap_8 FILLER_24_148 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_192 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_229 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_4 FILLER_24_302 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_104 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_decap_4 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_decap_4 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_decap_4 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_299 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_315 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_decap_4 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_107 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_214 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_decap_4 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_354 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_46 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_decap_4 FILLER_27_116 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_decap_8 FILLER_27_220 ();
 sg13g2_decap_4 FILLER_27_227 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_61 ();
 sg13g2_decap_4 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_decap_4 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_decap_4 FILLER_29_116 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_fill_1 FILLER_29_148 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_298 ();
 sg13g2_decap_4 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_322 ();
 sg13g2_decap_4 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_decap_4 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_94 ();
 sg13g2_decap_4 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_202 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_decap_4 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_298 ();
 sg13g2_decap_4 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_34 ();
 sg13g2_fill_2 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_301 ();
 sg13g2_decap_4 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_decap_4 FILLER_31_358 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_decap_4 FILLER_32_100 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_decap_4 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_190 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_decap_8 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_decap_8 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_55 ();
 sg13g2_decap_4 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_66 ();
 sg13g2_fill_2 FILLER_33_80 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_decap_4 FILLER_33_120 ();
 sg13g2_fill_2 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_fill_1 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_289 ();
 sg13g2_decap_4 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_decap_4 FILLER_33_352 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_fill_2 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_decap_4 FILLER_34_85 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_204 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_41 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_35_314 ();
 sg13g2_decap_8 FILLER_35_321 ();
 sg13g2_decap_8 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_361 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_18 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_204 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_33 ();
 sg13g2_fill_1 FILLER_37_47 ();
 sg13g2_decap_4 FILLER_37_57 ();
 sg13g2_fill_1 FILLER_37_61 ();
 sg13g2_fill_2 FILLER_37_92 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_229 ();
 sg13g2_fill_2 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_decap_4 FILLER_37_330 ();
 sg13g2_decap_4 FILLER_37_363 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_46 ();
 sg13g2_fill_2 FILLER_38_53 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_86 ();
 sg13g2_fill_1 FILLER_38_88 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_182 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_206 ();
 sg13g2_fill_2 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_fill_2 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
endmodule
