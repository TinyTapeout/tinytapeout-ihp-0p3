module tt_um_a1k0n_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire audio;
 wire hsync;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire \vgademo.a_cos[0] ;
 wire \vgademo.a_cos[10] ;
 wire \vgademo.a_cos[11] ;
 wire \vgademo.a_cos[12] ;
 wire \vgademo.a_cos[13] ;
 wire \vgademo.a_cos[14] ;
 wire \vgademo.a_cos[1] ;
 wire \vgademo.a_cos[2] ;
 wire \vgademo.a_cos[3] ;
 wire \vgademo.a_cos[4] ;
 wire \vgademo.a_cos[5] ;
 wire \vgademo.a_cos[6] ;
 wire \vgademo.a_cos[7] ;
 wire \vgademo.a_cos[8] ;
 wire \vgademo.a_cos[9] ;
 wire \vgademo.a_scrolly[10] ;
 wire \vgademo.a_scrolly[11] ;
 wire \vgademo.a_scrolly[12] ;
 wire \vgademo.a_scrolly[13] ;
 wire \vgademo.a_scrolly[3] ;
 wire \vgademo.a_scrolly[4] ;
 wire \vgademo.a_scrolly[5] ;
 wire \vgademo.a_scrolly[6] ;
 wire \vgademo.a_scrolly[7] ;
 wire \vgademo.a_scrolly[8] ;
 wire \vgademo.a_scrolly[9] ;
 wire \vgademo.a_sin[0] ;
 wire \vgademo.a_sin[10] ;
 wire \vgademo.a_sin[11] ;
 wire \vgademo.a_sin[12] ;
 wire \vgademo.a_sin[13] ;
 wire \vgademo.a_sin[14] ;
 wire \vgademo.a_sin[1] ;
 wire \vgademo.a_sin[2] ;
 wire \vgademo.a_sin[3] ;
 wire \vgademo.a_sin[4] ;
 wire \vgademo.a_sin[5] ;
 wire \vgademo.a_sin[6] ;
 wire \vgademo.a_sin[7] ;
 wire \vgademo.a_sin[8] ;
 wire \vgademo.a_sin[9] ;
 wire \vgademo.audio_beat_out[0] ;
 wire \vgademo.audio_beat_out[1] ;
 wire \vgademo.audio_beat_out[2] ;
 wire \vgademo.audio_beat_out[3] ;
 wire \vgademo.audio_beat_out[4] ;
 wire \vgademo.audio_kick_frames[0] ;
 wire \vgademo.audio_kick_frames[1] ;
 wire \vgademo.audio_kick_frames[2] ;
 wire \vgademo.audio_snare_frames[0] ;
 wire \vgademo.audio_snare_frames[1] ;
 wire \vgademo.audio_snare_frames[2] ;
 wire \vgademo.audio_snare_frames[3] ;
 wire \vgademo.audio_songpos[0] ;
 wire \vgademo.audio_songpos[1] ;
 wire \vgademo.audio_songpos[2] ;
 wire \vgademo.audio_songpos[3] ;
 wire \vgademo.audio_songpos[4] ;
 wire \vgademo.audio_songpos[5] ;
 wire \vgademo.audio_songpos[6] ;
 wire \vgademo.audio_songpos[7] ;
 wire \vgademo.b_cos[0] ;
 wire \vgademo.b_cos[10] ;
 wire \vgademo.b_cos[11] ;
 wire \vgademo.b_cos[1] ;
 wire \vgademo.b_cos[2] ;
 wire \vgademo.b_cos[3] ;
 wire \vgademo.b_cos[4] ;
 wire \vgademo.b_cos[5] ;
 wire \vgademo.b_cos[6] ;
 wire \vgademo.b_cos[7] ;
 wire \vgademo.b_cos[8] ;
 wire \vgademo.b_cos[9] ;
 wire \vgademo.b_sin[0] ;
 wire \vgademo.b_sin[10] ;
 wire \vgademo.b_sin[11] ;
 wire \vgademo.b_sin[1] ;
 wire \vgademo.b_sin[2] ;
 wire \vgademo.b_sin[3] ;
 wire \vgademo.b_sin[4] ;
 wire \vgademo.b_sin[5] ;
 wire \vgademo.b_sin[6] ;
 wire \vgademo.b_sin[7] ;
 wire \vgademo.b_sin[8] ;
 wire \vgademo.b_sin[9] ;
 wire \vgademo.bayer_j[0] ;
 wire \vgademo.bayer_j[1] ;
 wire \vgademo.h_count[0] ;
 wire \vgademo.h_count[10] ;
 wire \vgademo.h_count[1] ;
 wire \vgademo.h_count[2] ;
 wire \vgademo.h_count[3] ;
 wire \vgademo.h_count[4] ;
 wire \vgademo.h_count[5] ;
 wire \vgademo.h_count[6] ;
 wire \vgademo.h_count[7] ;
 wire \vgademo.h_count[8] ;
 wire \vgademo.h_count[9] ;
 wire \vgademo.linelfsr[0] ;
 wire \vgademo.linelfsr[10] ;
 wire \vgademo.linelfsr[11] ;
 wire \vgademo.linelfsr[12] ;
 wire \vgademo.linelfsr[1] ;
 wire \vgademo.linelfsr[2] ;
 wire \vgademo.linelfsr[3] ;
 wire \vgademo.linelfsr[4] ;
 wire \vgademo.linelfsr[5] ;
 wire \vgademo.linelfsr[6] ;
 wire \vgademo.linelfsr[7] ;
 wire \vgademo.linelfsr[8] ;
 wire \vgademo.linelfsr[9] ;
 wire \vgademo.plane_du[0] ;
 wire \vgademo.plane_du[10] ;
 wire \vgademo.plane_du[1] ;
 wire \vgademo.plane_du[2] ;
 wire \vgademo.plane_du[3] ;
 wire \vgademo.plane_du[4] ;
 wire \vgademo.plane_du[5] ;
 wire \vgademo.plane_du[6] ;
 wire \vgademo.plane_du[7] ;
 wire \vgademo.plane_du[8] ;
 wire \vgademo.plane_du[9] ;
 wire \vgademo.plane_dx[0] ;
 wire \vgademo.plane_dx[1] ;
 wire \vgademo.plane_dx[2] ;
 wire \vgademo.plane_dx[3] ;
 wire \vgademo.plane_dx_div.d[16] ;
 wire \vgademo.plane_dx_div.d[17] ;
 wire \vgademo.plane_dx_div.d[18] ;
 wire \vgademo.plane_dx_div.d[19] ;
 wire \vgademo.plane_dx_div.d[20] ;
 wire \vgademo.plane_dx_div.d[21] ;
 wire \vgademo.plane_dx_div.d[22] ;
 wire \vgademo.plane_dx_div.d[23] ;
 wire \vgademo.plane_dx_div.d[24] ;
 wire \vgademo.plane_dx_div.i[0] ;
 wire \vgademo.plane_dx_div.i[1] ;
 wire \vgademo.plane_dx_div.i[2] ;
 wire \vgademo.plane_dx_div.i[3] ;
 wire \vgademo.plane_dx_div.q[3] ;
 wire \vgademo.plane_dx_div.q[4] ;
 wire \vgademo.plane_dx_div.q[5] ;
 wire \vgademo.plane_dx_div.q[6] ;
 wire \vgademo.plane_dx_div.q[7] ;
 wire \vgademo.plane_dx_div.q[8] ;
 wire \vgademo.plane_dx_div.q[9] ;
 wire \vgademo.plane_dx_div.r[16] ;
 wire \vgademo.plane_dx_div.r[17] ;
 wire \vgademo.plane_dx_div.r[18] ;
 wire \vgademo.plane_dx_div.r[19] ;
 wire \vgademo.plane_dx_div.r[20] ;
 wire \vgademo.plane_dx_div.r[21] ;
 wire \vgademo.plane_dx_div.r[22] ;
 wire \vgademo.plane_dx_div.r[23] ;
 wire \vgademo.plane_dx_div.r[24] ;
 wire \vgademo.plane_dx_div.r[25] ;
 wire \vgademo.plane_u[0] ;
 wire \vgademo.plane_u[10] ;
 wire \vgademo.plane_u[11] ;
 wire \vgademo.plane_u[12] ;
 wire \vgademo.plane_u[13] ;
 wire \vgademo.plane_u[14] ;
 wire \vgademo.plane_u[15] ;
 wire \vgademo.plane_u[16] ;
 wire \vgademo.plane_u[17] ;
 wire \vgademo.plane_u[18] ;
 wire \vgademo.plane_u[19] ;
 wire \vgademo.plane_u[1] ;
 wire \vgademo.plane_u[20] ;
 wire \vgademo.plane_u[21] ;
 wire \vgademo.plane_u[2] ;
 wire \vgademo.plane_u[3] ;
 wire \vgademo.plane_u[4] ;
 wire \vgademo.plane_u[5] ;
 wire \vgademo.plane_u[6] ;
 wire \vgademo.plane_u[7] ;
 wire \vgademo.plane_u[8] ;
 wire \vgademo.plane_u[9] ;
 wire \vgademo.scanline_audio_sample[0] ;
 wire \vgademo.scanline_audio_sample[1] ;
 wire \vgademo.scanline_audio_sample[2] ;
 wire \vgademo.scanline_audio_sample[3] ;
 wire \vgademo.scanline_audio_sample[4] ;
 wire \vgademo.scanline_audio_sample[5] ;
 wire \vgademo.scanline_audio_sample[6] ;
 wire \vgademo.soundtrack.noise_lfsr[0] ;
 wire \vgademo.soundtrack.noise_lfsr[10] ;
 wire \vgademo.soundtrack.noise_lfsr[11] ;
 wire \vgademo.soundtrack.noise_lfsr[12] ;
 wire \vgademo.soundtrack.noise_lfsr[13] ;
 wire \vgademo.soundtrack.noise_lfsr[14] ;
 wire \vgademo.soundtrack.noise_lfsr[1] ;
 wire \vgademo.soundtrack.noise_lfsr[2] ;
 wire \vgademo.soundtrack.noise_lfsr[3] ;
 wire \vgademo.soundtrack.noise_lfsr[4] ;
 wire \vgademo.soundtrack.noise_lfsr[5] ;
 wire \vgademo.soundtrack.noise_lfsr[6] ;
 wire \vgademo.soundtrack.noise_lfsr[7] ;
 wire \vgademo.soundtrack.noise_lfsr[8] ;
 wire \vgademo.soundtrack.noise_lfsr[9] ;
 wire \vgademo.soundtrack.pulse_osc_p[0] ;
 wire \vgademo.soundtrack.pulse_osc_p[10] ;
 wire \vgademo.soundtrack.pulse_osc_p[11] ;
 wire \vgademo.soundtrack.pulse_osc_p[12] ;
 wire \vgademo.soundtrack.pulse_osc_p[13] ;
 wire \vgademo.soundtrack.pulse_osc_p[1] ;
 wire \vgademo.soundtrack.pulse_osc_p[2] ;
 wire \vgademo.soundtrack.pulse_osc_p[3] ;
 wire \vgademo.soundtrack.pulse_osc_p[4] ;
 wire \vgademo.soundtrack.pulse_osc_p[5] ;
 wire \vgademo.soundtrack.pulse_osc_p[6] ;
 wire \vgademo.soundtrack.pulse_osc_p[7] ;
 wire \vgademo.soundtrack.pulse_osc_p[8] ;
 wire \vgademo.soundtrack.pulse_osc_p[9] ;
 wire \vgademo.soundtrack.pulse_vol[0] ;
 wire \vgademo.soundtrack.pulse_vol[1] ;
 wire \vgademo.soundtrack.pulse_vol[2] ;
 wire \vgademo.soundtrack.pulse_vol[3] ;
 wire \vgademo.soundtrack.sample_div[0] ;
 wire \vgademo.soundtrack.sample_div[1] ;
 wire \vgademo.soundtrack.sample_div[2] ;
 wire \vgademo.soundtrack.sample_div[3] ;
 wire \vgademo.soundtrack.sample_div[4] ;
 wire \vgademo.soundtrack.sample_div[5] ;
 wire \vgademo.soundtrack.sample_div[6] ;
 wire \vgademo.soundtrack.sample_div[7] ;
 wire \vgademo.soundtrack.sample_div[8] ;
 wire \vgademo.soundtrack.sample_div[9] ;
 wire \vgademo.soundtrack.sample_div_[0] ;
 wire \vgademo.soundtrack.sample_div_[1] ;
 wire \vgademo.soundtrack.sample_div_[2] ;
 wire \vgademo.soundtrack.sample_div_[3] ;
 wire \vgademo.soundtrack.sample_div_[4] ;
 wire \vgademo.soundtrack.sample_div_[5] ;
 wire \vgademo.soundtrack.sample_div_[6] ;
 wire \vgademo.soundtrack.sample_div_[7] ;
 wire \vgademo.soundtrack.sample_div_[8] ;
 wire \vgademo.soundtrack.sample_div_[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[9] ;
 wire \vgademo.soundtrack.tick_div[0] ;
 wire \vgademo.soundtrack.tick_div[1] ;
 wire \vgademo.soundtrack.tick_div[2] ;
 wire \vgademo.soundtrack.tick_div[3] ;
 wire \vgademo.soundtrack.tick_div[4] ;
 wire \vgademo.soundtrack.tick_div[5] ;
 wire \vgademo.soundtrack.tick_div[6] ;
 wire \vgademo.soundtrack.tick_div[7] ;
 wire \vgademo.soundtrack.tick_div_[0] ;
 wire \vgademo.soundtrack.tri_osc_i[0] ;
 wire \vgademo.soundtrack.tri_osc_i[1] ;
 wire \vgademo.soundtrack.tri_osc_i[2] ;
 wire \vgademo.soundtrack.tri_osc_i[3] ;
 wire \vgademo.soundtrack.tri_osc_i[4] ;
 wire \vgademo.soundtrack.tri_osc_i[5] ;
 wire \vgademo.soundtrack.tri_osc_i[6] ;
 wire \vgademo.soundtrack.tri_osc_i[7] ;
 wire \vgademo.soundtrack.tri_osc_i[8] ;
 wire \vgademo.soundtrack.tri_osc_p[0] ;
 wire \vgademo.soundtrack.tri_osc_p[10] ;
 wire \vgademo.soundtrack.tri_osc_p[11] ;
 wire \vgademo.soundtrack.tri_osc_p[12] ;
 wire \vgademo.soundtrack.tri_osc_p[13] ;
 wire \vgademo.soundtrack.tri_osc_p[14] ;
 wire \vgademo.soundtrack.tri_osc_p[15] ;
 wire \vgademo.soundtrack.tri_osc_p[1] ;
 wire \vgademo.soundtrack.tri_osc_p[2] ;
 wire \vgademo.soundtrack.tri_osc_p[3] ;
 wire \vgademo.soundtrack.tri_osc_p[4] ;
 wire \vgademo.soundtrack.tri_osc_p[5] ;
 wire \vgademo.soundtrack.tri_osc_p[6] ;
 wire \vgademo.soundtrack.tri_osc_p[7] ;
 wire \vgademo.soundtrack.tri_osc_p[8] ;
 wire \vgademo.soundtrack.tri_osc_p[9] ;
 wire \vgademo.v_count[2] ;
 wire \vgademo.v_count[3] ;
 wire \vgademo.v_count[4] ;
 wire \vgademo.v_count[5] ;
 wire \vgademo.v_count[6] ;
 wire \vgademo.v_count[7] ;
 wire \vgademo.v_count[8] ;
 wire \vgademo.v_count[9] ;
 wire \vgademo.vsync ;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;

 sg13g2_inv_1 _3739_ (.Y(_3094_),
    .A(\vgademo.soundtrack.noise_lfsr[2] ));
 sg13g2_inv_1 _3740_ (.Y(_3095_),
    .A(net168));
 sg13g2_inv_1 _3741_ (.Y(_3096_),
    .A(net1011));
 sg13g2_inv_1 _3742_ (.Y(_3097_),
    .A(net591));
 sg13g2_inv_1 _3743_ (.Y(_3098_),
    .A(net544));
 sg13g2_inv_1 _3744_ (.Y(_3099_),
    .A(net557));
 sg13g2_inv_1 _3745_ (.Y(_3100_),
    .A(net209));
 sg13g2_inv_1 _3746_ (.Y(_3101_),
    .A(net331));
 sg13g2_inv_2 _3747_ (.Y(_3102_),
    .A(net948));
 sg13g2_inv_1 _3748_ (.Y(_3103_),
    .A(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_inv_1 _3749_ (.Y(_3104_),
    .A(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_inv_1 _3750_ (.Y(_3105_),
    .A(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_inv_1 _3751_ (.Y(_3106_),
    .A(net450));
 sg13g2_inv_1 _3752_ (.Y(_3107_),
    .A(\vgademo.audio_beat_out[2] ));
 sg13g2_inv_2 _3753_ (.Y(_3108_),
    .A(net1035));
 sg13g2_inv_1 _3754_ (.Y(_3109_),
    .A(net1024));
 sg13g2_inv_1 _3755_ (.Y(_3110_),
    .A(net1029));
 sg13g2_inv_1 _3756_ (.Y(_3111_),
    .A(net1021));
 sg13g2_inv_1 _3757_ (.Y(_3112_),
    .A(\vgademo.audio_songpos[6] ));
 sg13g2_inv_2 _3758_ (.Y(_3113_),
    .A(net577));
 sg13g2_inv_2 _3759_ (.Y(_3114_),
    .A(_0060_));
 sg13g2_inv_2 _3760_ (.Y(_3115_),
    .A(\vgademo.bayer_j[0] ));
 sg13g2_inv_2 _3761_ (.Y(_3116_),
    .A(\vgademo.v_count[2] ));
 sg13g2_inv_1 _3762_ (.Y(_3117_),
    .A(\vgademo.v_count[3] ));
 sg13g2_inv_1 _3763_ (.Y(_3118_),
    .A(\vgademo.v_count[5] ));
 sg13g2_inv_2 _3764_ (.Y(_3119_),
    .A(net986));
 sg13g2_inv_1 _3765_ (.Y(_3120_),
    .A(\vgademo.h_count[0] ));
 sg13g2_inv_1 _3766_ (.Y(_3121_),
    .A(net985));
 sg13g2_inv_2 _3767_ (.Y(_3122_),
    .A(\vgademo.h_count[2] ));
 sg13g2_inv_2 _3768_ (.Y(_3123_),
    .A(\vgademo.h_count[4] ));
 sg13g2_inv_1 _3769_ (.Y(_3124_),
    .A(\vgademo.h_count[5] ));
 sg13g2_inv_2 _3770_ (.Y(_3125_),
    .A(\vgademo.h_count[7] ));
 sg13g2_inv_2 _3771_ (.Y(_3126_),
    .A(net585));
 sg13g2_inv_2 _3772_ (.Y(_3127_),
    .A(net982));
 sg13g2_inv_2 _3773_ (.Y(_3128_),
    .A(_0063_));
 sg13g2_inv_4 _3774_ (.A(net980),
    .Y(_3129_));
 sg13g2_inv_2 _3775_ (.Y(_3130_),
    .A(net961));
 sg13g2_inv_2 _3776_ (.Y(_3131_),
    .A(net962));
 sg13g2_inv_1 _3777_ (.Y(_3132_),
    .A(net964));
 sg13g2_inv_4 _3778_ (.A(\vgademo.a_scrolly[8] ),
    .Y(_3133_));
 sg13g2_inv_2 _3779_ (.Y(_3134_),
    .A(net973));
 sg13g2_inv_2 _3780_ (.Y(_3135_),
    .A(net975));
 sg13g2_inv_1 _3781_ (.Y(_3136_),
    .A(net978));
 sg13g2_inv_2 _3782_ (.Y(_3137_),
    .A(_0066_));
 sg13g2_inv_1 _3783_ (.Y(_3138_),
    .A(_0064_));
 sg13g2_inv_1 _3784_ (.Y(_3139_),
    .A(_0069_));
 sg13g2_inv_1 _3785_ (.Y(_3140_),
    .A(_0078_));
 sg13g2_inv_1 _3786_ (.Y(_3141_),
    .A(\vgademo.plane_dx_div.r[20] ));
 sg13g2_inv_1 _3787_ (.Y(_3142_),
    .A(_0018_));
 sg13g2_inv_1 _3788_ (.Y(_3143_),
    .A(_0020_));
 sg13g2_inv_1 _3789_ (.Y(_3144_),
    .A(net339));
 sg13g2_inv_1 _3790_ (.Y(_3145_),
    .A(net325));
 sg13g2_inv_1 _3791_ (.Y(_3146_),
    .A(\vgademo.soundtrack.tri_osc_i[1] ));
 sg13g2_inv_1 _3792_ (.Y(_3147_),
    .A(net586));
 sg13g2_inv_1 _3793_ (.Y(_3148_),
    .A(net564));
 sg13g2_inv_1 _3794_ (.Y(_3149_),
    .A(net521));
 sg13g2_inv_1 _3795_ (.Y(_3150_),
    .A(\vgademo.soundtrack.pulse_vol[2] ));
 sg13g2_inv_1 _3796_ (.Y(_3151_),
    .A(net1001));
 sg13g2_inv_2 _3797_ (.Y(_3152_),
    .A(net994));
 sg13g2_inv_1 _3798_ (.Y(_3153_),
    .A(net996));
 sg13g2_inv_1 _3799_ (.Y(_3154_),
    .A(net528));
 sg13g2_inv_1 _3800_ (.Y(_3155_),
    .A(\vgademo.b_sin[9] ));
 sg13g2_inv_1 _3801_ (.Y(_3156_),
    .A(\vgademo.a_cos[6] ));
 sg13g2_inv_1 _3802_ (.Y(_3157_),
    .A(net443));
 sg13g2_inv_2 _3803_ (.Y(_3158_),
    .A(net946));
 sg13g2_inv_1 _3804_ (.Y(_3159_),
    .A(net515));
 sg13g2_inv_1 _3805_ (.Y(_3160_),
    .A(\vgademo.b_cos[7] ));
 sg13g2_inv_2 _3806_ (.Y(_3161_),
    .A(\vgademo.b_cos[8] ));
 sg13g2_inv_2 _3807_ (.Y(_3162_),
    .A(\vgademo.b_cos[9] ));
 sg13g2_inv_1 _3808_ (.Y(_3163_),
    .A(net951));
 sg13g2_inv_1 _3809_ (.Y(_3164_),
    .A(net385));
 sg13g2_inv_1 _3810_ (.Y(_3165_),
    .A(net365));
 sg13g2_inv_1 _3811_ (.Y(_3166_),
    .A(net448));
 sg13g2_inv_2 _3812_ (.Y(_3167_),
    .A(net529));
 sg13g2_inv_1 _3813_ (.Y(_3168_),
    .A(\vgademo.a_sin[9] ));
 sg13g2_inv_1 _3814_ (.Y(_3169_),
    .A(net523));
 sg13g2_inv_1 _3815_ (.Y(_3170_),
    .A(\vgademo.a_sin[12] ));
 sg13g2_inv_2 _3816_ (.Y(_3171_),
    .A(\vgademo.a_sin[14] ));
 sg13g2_inv_1 _3817_ (.Y(_3172_),
    .A(net383));
 sg13g2_inv_1 _3818_ (.Y(_3173_),
    .A(\vgademo.plane_du[3] ));
 sg13g2_inv_1 _3819_ (.Y(_3174_),
    .A(net318));
 sg13g2_inv_2 _3820_ (.Y(_3175_),
    .A(\vgademo.plane_du[4] ));
 sg13g2_inv_1 _3821_ (.Y(_3176_),
    .A(net337));
 sg13g2_inv_1 _3822_ (.Y(_3177_),
    .A(_0022_));
 sg13g2_inv_1 _3823_ (.Y(_3178_),
    .A(net353));
 sg13g2_inv_1 _3824_ (.Y(_3179_),
    .A(net574));
 sg13g2_inv_1 _3825_ (.Y(_3180_),
    .A(net364));
 sg13g2_inv_1 _3826_ (.Y(_3181_),
    .A(\vgademo.plane_du[7] ));
 sg13g2_inv_1 _3827_ (.Y(_3182_),
    .A(net327));
 sg13g2_inv_1 _3828_ (.Y(_3183_),
    .A(_0025_));
 sg13g2_inv_1 _3829_ (.Y(_3184_),
    .A(net435));
 sg13g2_inv_2 _3830_ (.Y(_3185_),
    .A(\vgademo.plane_du[9] ));
 sg13g2_inv_1 _3831_ (.Y(_3186_),
    .A(net373));
 sg13g2_inv_1 _3832_ (.Y(_3187_),
    .A(net296));
 sg13g2_inv_1 _3833_ (.Y(_3188_),
    .A(net360));
 sg13g2_inv_1 _3834_ (.Y(_3189_),
    .A(net381));
 sg13g2_inv_1 _3835_ (.Y(_3190_),
    .A(\vgademo.plane_u[14] ));
 sg13g2_inv_1 _3836_ (.Y(_3191_),
    .A(net580));
 sg13g2_inv_1 _3837_ (.Y(_3192_),
    .A(net465));
 sg13g2_inv_1 _3838_ (.Y(_3193_),
    .A(net445));
 sg13g2_inv_1 _3839_ (.Y(_3194_),
    .A(net328));
 sg13g2_inv_1 _3840_ (.Y(_3195_),
    .A(net399));
 sg13g2_inv_1 _3841_ (.Y(_3196_),
    .A(net234));
 sg13g2_inv_1 _3842_ (.Y(_3197_),
    .A(net1040));
 sg13g2_inv_1 _3843_ (.Y(_3198_),
    .A(net392));
 sg13g2_inv_1 _3844_ (.Y(_3199_),
    .A(net375));
 sg13g2_inv_1 _3845_ (.Y(_3200_),
    .A(net370));
 sg13g2_inv_1 _3846_ (.Y(_3201_),
    .A(\vgademo.soundtrack.pulse_osc_p[12] ));
 sg13g2_inv_1 _3847_ (.Y(_3202_),
    .A(net368));
 sg13g2_inv_1 _3848_ (.Y(_3203_),
    .A(net428));
 sg13g2_inv_1 _3849_ (.Y(_3204_),
    .A(net470));
 sg13g2_inv_1 _3850_ (.Y(_3205_),
    .A(net415));
 sg13g2_inv_1 _3851_ (.Y(_3206_),
    .A(net309));
 sg13g2_inv_1 _3852_ (.Y(_3207_),
    .A(net322));
 sg13g2_inv_1 _3853_ (.Y(_3208_),
    .A(net295));
 sg13g2_inv_1 _3854_ (.Y(_3209_),
    .A(\vgademo.scanline_audio_sample[3] ));
 sg13g2_nand2_2 _3855_ (.Y(_3210_),
    .A(\vgademo.h_count[7] ),
    .B(\vgademo.h_count[6] ));
 sg13g2_nor3_2 _3856_ (.A(_3123_),
    .B(net941),
    .C(_3210_),
    .Y(_3211_));
 sg13g2_nor4_2 _3857_ (.A(net986),
    .B(\vgademo.h_count[0] ),
    .C(net985),
    .Y(_3212_),
    .D(_3122_));
 sg13g2_inv_1 _3858_ (.Y(_3213_),
    .A(_3212_));
 sg13g2_nor2_1 _3859_ (.A(\vgademo.h_count[9] ),
    .B(net982),
    .Y(_3214_));
 sg13g2_and4_2 _3860_ (.A(\vgademo.h_count[8] ),
    .B(_3211_),
    .C(_3212_),
    .D(_3214_),
    .X(_3215_));
 sg13g2_nand4_1 _3861_ (.B(_3211_),
    .C(_3212_),
    .A(net983),
    .Y(_3216_),
    .D(_3214_));
 sg13g2_and4_1 _3862_ (.A(net983),
    .B(_3211_),
    .C(_3212_),
    .D(_3214_),
    .X(_3217_));
 sg13g2_nor2_1 _3863_ (.A(net555),
    .B(_3215_),
    .Y(_0000_));
 sg13g2_nand2_2 _3864_ (.Y(_3218_),
    .A(net986),
    .B(\vgademo.h_count[0] ));
 sg13g2_xor2_1 _3865_ (.B(net555),
    .A(net986),
    .X(_0002_));
 sg13g2_nor2_1 _3866_ (.A(net469),
    .B(_3218_),
    .Y(_3219_));
 sg13g2_and2_1 _3867_ (.A(net469),
    .B(_3218_),
    .X(_3220_));
 sg13g2_nor3_1 _3868_ (.A(_3215_),
    .B(_3219_),
    .C(_3220_),
    .Y(_0003_));
 sg13g2_xor2_1 _3869_ (.B(_3219_),
    .A(net459),
    .X(_3221_));
 sg13g2_nor2_1 _3870_ (.A(_3215_),
    .B(net460),
    .Y(_0004_));
 sg13g2_nand2_1 _3871_ (.Y(_3222_),
    .A(\vgademo.h_count[1] ),
    .B(\vgademo.h_count[2] ));
 sg13g2_nor3_2 _3872_ (.A(_3121_),
    .B(_3122_),
    .C(_3218_),
    .Y(_3223_));
 sg13g2_and2_1 _3873_ (.A(\vgademo.h_count[4] ),
    .B(_3223_),
    .X(_3224_));
 sg13g2_nor2_1 _3874_ (.A(net541),
    .B(_3223_),
    .Y(_3225_));
 sg13g2_nor3_1 _3875_ (.A(_3215_),
    .B(_3224_),
    .C(_3225_),
    .Y(_0005_));
 sg13g2_xor2_1 _3876_ (.B(_3224_),
    .A(net475),
    .X(_3226_));
 sg13g2_nor2_1 _3877_ (.A(_3217_),
    .B(_3226_),
    .Y(_0006_));
 sg13g2_nand2_2 _3878_ (.Y(_3227_),
    .A(\vgademo.h_count[5] ),
    .B(_3224_));
 sg13g2_o21ai_1 _3879_ (.B1(net931),
    .Y(_3228_),
    .A1(net552),
    .A2(_3227_));
 sg13g2_a21oi_1 _3880_ (.A1(net552),
    .A2(_3227_),
    .Y(_0007_),
    .B1(_3228_));
 sg13g2_nor3_1 _3881_ (.A(net588),
    .B(net433),
    .C(_3227_),
    .Y(_3229_));
 sg13g2_o21ai_1 _3882_ (.B1(net433),
    .Y(_3230_),
    .A1(net588),
    .A2(_3227_));
 sg13g2_nand2_1 _3883_ (.Y(_3231_),
    .A(net931),
    .B(_3230_));
 sg13g2_nor2_1 _3884_ (.A(_3229_),
    .B(_3231_),
    .Y(_0008_));
 sg13g2_o21ai_1 _3885_ (.B1(net560),
    .Y(_3232_),
    .A1(_3210_),
    .A2(_3227_));
 sg13g2_inv_1 _3886_ (.Y(_3233_),
    .A(net561));
 sg13g2_nor3_2 _3887_ (.A(net560),
    .B(_3210_),
    .C(_3227_),
    .Y(_3234_));
 sg13g2_nor3_1 _3888_ (.A(_3215_),
    .B(_3233_),
    .C(_3234_),
    .Y(_0009_));
 sg13g2_o21ai_1 _3889_ (.B1(net930),
    .Y(_3235_),
    .A1(_3196_),
    .A2(_3234_));
 sg13g2_a21oi_1 _3890_ (.A1(_3196_),
    .A2(_3234_),
    .Y(_0010_),
    .B1(_3235_));
 sg13g2_nand4_1 _3891_ (.B(\vgademo.h_count[8] ),
    .C(_3211_),
    .A(\vgademo.h_count[9] ),
    .Y(_3236_),
    .D(_3223_));
 sg13g2_o21ai_1 _3892_ (.B1(net930),
    .Y(_3237_),
    .A1(net272),
    .A2(_3236_));
 sg13g2_a21oi_1 _3893_ (.A1(net982),
    .A2(_3236_),
    .Y(_0001_),
    .B1(net273));
 sg13g2_nand2_2 _3894_ (.Y(_3238_),
    .A(\vgademo.v_count[7] ),
    .B(\vgademo.v_count[6] ));
 sg13g2_nor3_1 _3895_ (.A(net960),
    .B(_3118_),
    .C(_3238_),
    .Y(_3239_));
 sg13g2_nor2b_1 _3896_ (.A(net955),
    .B_N(\vgademo.v_count[8] ),
    .Y(_3240_));
 sg13g2_nand4_1 _3897_ (.B(\vgademo.v_count[3] ),
    .C(_3239_),
    .A(\vgademo.bayer_j[1] ),
    .Y(_3241_),
    .D(_3240_));
 sg13g2_nor2_1 _3898_ (.A(_0063_),
    .B(_3238_),
    .Y(_3242_));
 sg13g2_nand2_2 _3899_ (.Y(_3243_),
    .A(\vgademo.v_count[2] ),
    .B(\vgademo.v_count[3] ));
 sg13g2_nor2_2 _3900_ (.A(\vgademo.bayer_j[1] ),
    .B(\vgademo.bayer_j[0] ),
    .Y(_3244_));
 sg13g2_o21ai_1 _3901_ (.B1(_3242_),
    .Y(_3245_),
    .A1(_3243_),
    .A2(_3244_));
 sg13g2_or3_1 _3902_ (.A(\vgademo.bayer_j[0] ),
    .B(\vgademo.v_count[2] ),
    .C(_3242_),
    .X(_3246_));
 sg13g2_a21o_1 _3903_ (.A2(_3246_),
    .A1(_3245_),
    .B1(_3241_),
    .X(_0012_));
 sg13g2_nand2_2 _3904_ (.Y(_3247_),
    .A(_3119_),
    .B(_3122_));
 sg13g2_nand3_1 _3905_ (.B(\vgademo.h_count[4] ),
    .C(_3247_),
    .A(\vgademo.h_count[3] ),
    .Y(_3248_));
 sg13g2_nand2b_1 _3906_ (.Y(_3249_),
    .B(_3248_),
    .A_N(net984));
 sg13g2_o21ai_1 _3907_ (.B1(\vgademo.h_count[7] ),
    .Y(_3250_),
    .A1(\vgademo.h_count[5] ),
    .A2(_3249_));
 sg13g2_nand2_1 _3908_ (.Y(_3251_),
    .A(\vgademo.h_count[10] ),
    .B(_3250_));
 sg13g2_o21ai_1 _3909_ (.B1(\vgademo.h_count[10] ),
    .Y(_3252_),
    .A1(net983),
    .A2(_3211_));
 sg13g2_nor2_1 _3910_ (.A(\vgademo.h_count[3] ),
    .B(\vgademo.h_count[2] ),
    .Y(_3253_));
 sg13g2_a21oi_1 _3911_ (.A1(_3127_),
    .A2(_3253_),
    .Y(_3254_),
    .B1(\vgademo.h_count[10] ));
 sg13g2_nor3_1 _3912_ (.A(\vgademo.h_count[4] ),
    .B(_3124_),
    .C(_3210_),
    .Y(_3255_));
 sg13g2_a21oi_1 _3913_ (.A1(_3218_),
    .A2(_3253_),
    .Y(_3256_),
    .B1(_3254_));
 sg13g2_nand2_1 _3914_ (.Y(_3257_),
    .A(_3255_),
    .B(_3256_));
 sg13g2_a22oi_1 _3915_ (.Y(_3258_),
    .B1(_3252_),
    .B2(_3257_),
    .A2(_3251_),
    .A1(net983));
 sg13g2_nand2_2 _3916_ (.Y(_0011_),
    .A(_3126_),
    .B(_3258_));
 sg13g2_nor2_1 _3917_ (.A(net991),
    .B(_3150_),
    .Y(_3259_));
 sg13g2_nor2_1 _3918_ (.A(_3108_),
    .B(net1032),
    .Y(_3260_));
 sg13g2_nand2b_2 _3919_ (.Y(_3261_),
    .B(net1035),
    .A_N(net1032));
 sg13g2_nand3b_1 _3920_ (.B(net1027),
    .C(net1034),
    .Y(_3262_),
    .A_N(net1031));
 sg13g2_nor2b_1 _3921_ (.A(net1036),
    .B_N(net1034),
    .Y(_3263_));
 sg13g2_nor2b_2 _3922_ (.A(net1035),
    .B_N(net1036),
    .Y(_3264_));
 sg13g2_nor2_1 _3923_ (.A(net1036),
    .B(net1030),
    .Y(_3265_));
 sg13g2_nor2_2 _3924_ (.A(_3108_),
    .B(net1028),
    .Y(_3266_));
 sg13g2_nand2_1 _3925_ (.Y(_3267_),
    .A(net1034),
    .B(net944));
 sg13g2_nor3_1 _3926_ (.A(_3264_),
    .B(_3265_),
    .C(_3266_),
    .Y(_3268_));
 sg13g2_nor2_2 _3927_ (.A(net1027),
    .B(net1031),
    .Y(_3269_));
 sg13g2_or2_1 _3928_ (.X(_3270_),
    .B(net1030),
    .A(net1029));
 sg13g2_nor2_2 _3929_ (.A(net1023),
    .B(_3269_),
    .Y(_3271_));
 sg13g2_nor2b_1 _3930_ (.A(_3268_),
    .B_N(_3271_),
    .Y(_3272_));
 sg13g2_nand2_1 _3931_ (.Y(_3273_),
    .A(net1035),
    .B(net1032));
 sg13g2_nor2_2 _3932_ (.A(net1038),
    .B(_3273_),
    .Y(_3274_));
 sg13g2_nand3b_1 _3933_ (.B(net1034),
    .C(net1031),
    .Y(_3275_),
    .A_N(net1036));
 sg13g2_and2_1 _3934_ (.A(net1027),
    .B(_3275_),
    .X(_3276_));
 sg13g2_nand2_1 _3935_ (.Y(_3277_),
    .A(net1027),
    .B(_3275_));
 sg13g2_and2_2 _3936_ (.A(net1037),
    .B(net1034),
    .X(_3278_));
 sg13g2_nand2_2 _3937_ (.Y(_3279_),
    .A(net1036),
    .B(net1035));
 sg13g2_nor2_2 _3938_ (.A(net1036),
    .B(net1034),
    .Y(_3280_));
 sg13g2_xor2_1 _3939_ (.B(net1034),
    .A(net1036),
    .X(_3281_));
 sg13g2_and2_1 _3940_ (.A(net944),
    .B(_3281_),
    .X(_3282_));
 sg13g2_nor3_1 _3941_ (.A(_3269_),
    .B(_3276_),
    .C(_3282_),
    .Y(_3283_));
 sg13g2_nor2_1 _3942_ (.A(net1031),
    .B(_3263_),
    .Y(_3284_));
 sg13g2_nor2_1 _3943_ (.A(net1031),
    .B(_3281_),
    .Y(_3285_));
 sg13g2_mux2_1 _3944_ (.A0(_3277_),
    .A1(net1027),
    .S(_3285_),
    .X(_3286_));
 sg13g2_nor2_2 _3945_ (.A(net945),
    .B(net1020),
    .Y(_3287_));
 sg13g2_mux2_1 _3946_ (.A0(net1036),
    .A1(_3263_),
    .S(_3262_),
    .X(_3288_));
 sg13g2_nand2_1 _3947_ (.Y(_3289_),
    .A(_3287_),
    .B(_3288_));
 sg13g2_nand2_1 _3948_ (.Y(_3290_),
    .A(net1016),
    .B(_3289_));
 sg13g2_o21ai_1 _3949_ (.B1(net945),
    .Y(_3291_),
    .A1(_3283_),
    .A2(_3284_));
 sg13g2_a21oi_1 _3950_ (.A1(net1023),
    .A2(_3286_),
    .Y(_3292_),
    .B1(net942));
 sg13g2_a221oi_1 _3951_ (.B2(_3292_),
    .C1(_3290_),
    .B1(_3291_),
    .A1(net942),
    .Y(_3293_),
    .A2(_3272_));
 sg13g2_nor3_1 _3952_ (.A(net942),
    .B(_3271_),
    .C(_3280_),
    .Y(_3294_));
 sg13g2_nor2_2 _3953_ (.A(net1024),
    .B(net1021),
    .Y(_3295_));
 sg13g2_nand2_1 _3954_ (.Y(_3296_),
    .A(net945),
    .B(net942));
 sg13g2_nand2_1 _3955_ (.Y(_3297_),
    .A(net1028),
    .B(net1032));
 sg13g2_o21ai_1 _3956_ (.B1(_3297_),
    .Y(_3298_),
    .A1(_3108_),
    .A2(net944));
 sg13g2_nand2b_2 _3957_ (.Y(_3299_),
    .B(net1027),
    .A_N(net1034));
 sg13g2_inv_1 _3958_ (.Y(_3300_),
    .A(_3299_));
 sg13g2_nor2_1 _3959_ (.A(net1032),
    .B(_3299_),
    .Y(_3301_));
 sg13g2_nand2b_1 _3960_ (.Y(_3302_),
    .B(net1037),
    .A_N(net1030));
 sg13g2_nor4_1 _3961_ (.A(net945),
    .B(net1020),
    .C(_3299_),
    .D(_3302_),
    .Y(_3303_));
 sg13g2_nor2_1 _3962_ (.A(net1016),
    .B(_3303_),
    .Y(_3304_));
 sg13g2_o21ai_1 _3963_ (.B1(_3304_),
    .Y(_3305_),
    .A1(_3296_),
    .A2(_3298_));
 sg13g2_o21ai_1 _3964_ (.B1(net1019),
    .Y(_3306_),
    .A1(_3294_),
    .A2(_3305_));
 sg13g2_o21ai_1 _3965_ (.B1(\vgademo.soundtrack.pulse_osc_p[13] ),
    .Y(_3307_),
    .A1(_3293_),
    .A2(_3306_));
 sg13g2_or3_2 _3966_ (.A(_3201_),
    .B(_3293_),
    .C(_3306_),
    .X(_3308_));
 sg13g2_nand2_1 _3967_ (.Y(_3309_),
    .A(_3307_),
    .B(_3308_));
 sg13g2_nand3_1 _3968_ (.B(_3307_),
    .C(_3308_),
    .A(\vgademo.soundtrack.pulse_vol[0] ),
    .Y(_3310_));
 sg13g2_nand3_1 _3969_ (.B(_3259_),
    .C(_3310_),
    .A(net989),
    .Y(_3311_));
 sg13g2_nor2_1 _3970_ (.A(net1003),
    .B(_0040_),
    .Y(_3312_));
 sg13g2_a21oi_1 _3971_ (.A1(net1003),
    .A2(\vgademo.soundtrack.noise_lfsr[5] ),
    .Y(_3313_),
    .B1(_3312_));
 sg13g2_nor2_1 _3972_ (.A(net1000),
    .B(_3313_),
    .Y(_3314_));
 sg13g2_mux2_1 _3973_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(\vgademo.soundtrack.noise_lfsr[7] ),
    .S(net1005),
    .X(_3315_));
 sg13g2_a21oi_1 _3974_ (.A1(net1000),
    .A2(_3315_),
    .Y(_3316_),
    .B1(_3314_));
 sg13g2_nor2_1 _3975_ (.A(\vgademo.soundtrack.noise_lfsr[2] ),
    .B(net1002),
    .Y(_3317_));
 sg13g2_nor2b_1 _3976_ (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .B_N(net1002),
    .Y(_3318_));
 sg13g2_mux4_1 _3977_ (.S0(net1002),
    .A0(\vgademo.soundtrack.noise_lfsr[0] ),
    .A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(\vgademo.soundtrack.noise_lfsr[2] ),
    .A3(\vgademo.soundtrack.noise_lfsr[3] ),
    .S1(net1000),
    .X(_3319_));
 sg13g2_mux2_1 _3978_ (.A0(\vgademo.soundtrack.noise_lfsr[10] ),
    .A1(\vgademo.soundtrack.noise_lfsr[11] ),
    .S(net1003),
    .X(_3320_));
 sg13g2_nand2_1 _3979_ (.Y(_3321_),
    .A(net1000),
    .B(_3320_));
 sg13g2_nand2b_1 _3980_ (.Y(_3322_),
    .B(net1006),
    .A_N(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_o21ai_1 _3981_ (.B1(_3322_),
    .Y(_3323_),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .A2(net1005));
 sg13g2_o21ai_1 _3982_ (.B1(_3321_),
    .Y(_3324_),
    .A1(net1000),
    .A2(_3323_));
 sg13g2_nor2_1 _3983_ (.A(net998),
    .B(_3324_),
    .Y(_3325_));
 sg13g2_nand3b_1 _3984_ (.B(\vgademo.soundtrack.noise_lfsr[12] ),
    .C(net937),
    .Y(_3326_),
    .A_N(net1004));
 sg13g2_a21oi_1 _3985_ (.A1(net996),
    .A2(_3326_),
    .Y(_3327_),
    .B1(_3325_));
 sg13g2_nand2_1 _3986_ (.Y(_3328_),
    .A(net994),
    .B(_3327_));
 sg13g2_a21oi_1 _3987_ (.A1(net996),
    .A2(_3316_),
    .Y(_3329_),
    .B1(net993));
 sg13g2_o21ai_1 _3988_ (.B1(_3329_),
    .Y(_3330_),
    .A1(net996),
    .A2(_3319_));
 sg13g2_nand2_2 _3989_ (.Y(_3331_),
    .A(_3328_),
    .B(_3330_));
 sg13g2_inv_1 _3990_ (.Y(_3332_),
    .A(_3331_));
 sg13g2_nand2b_1 _3991_ (.Y(_3333_),
    .B(_3331_),
    .A_N(_3311_));
 sg13g2_and2_1 _3992_ (.A(_3311_),
    .B(_3332_),
    .X(_3334_));
 sg13g2_xnor2_1 _3993_ (.Y(_3335_),
    .A(_3311_),
    .B(_3331_));
 sg13g2_xnor2_1 _3994_ (.Y(_3336_),
    .A(net987),
    .B(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_xnor2_1 _3995_ (.Y(_3337_),
    .A(_3335_),
    .B(_3336_));
 sg13g2_nand2_1 _3996_ (.Y(_3338_),
    .A(net224),
    .B(_3337_));
 sg13g2_xor2_1 _3997_ (.B(_3337_),
    .A(net224),
    .X(\vgademo.soundtrack.sigma_delta_accum_[0] ));
 sg13g2_nand2_2 _3998_ (.Y(_3339_),
    .A(net991),
    .B(\vgademo.soundtrack.pulse_vol[2] ));
 sg13g2_inv_1 _3999_ (.Y(_3340_),
    .A(_3339_));
 sg13g2_nand2_1 _4000_ (.Y(_3341_),
    .A(net990),
    .B(_3340_));
 sg13g2_xor2_1 _4001_ (.B(_3339_),
    .A(net989),
    .X(_3342_));
 sg13g2_inv_1 _4002_ (.Y(_3343_),
    .A(_3342_));
 sg13g2_nor2_2 _4003_ (.A(net991),
    .B(\vgademo.soundtrack.pulse_vol[2] ),
    .Y(_3344_));
 sg13g2_nor2_1 _4004_ (.A(_3340_),
    .B(_3344_),
    .Y(_3345_));
 sg13g2_or2_1 _4005_ (.X(_3346_),
    .B(_3344_),
    .A(_3340_));
 sg13g2_and2_1 _4006_ (.A(net992),
    .B(\vgademo.soundtrack.pulse_vol[1] ),
    .X(_3347_));
 sg13g2_nand2_1 _4007_ (.Y(_3348_),
    .A(net992),
    .B(\vgademo.soundtrack.pulse_vol[1] ));
 sg13g2_nor2_1 _4008_ (.A(net992),
    .B(net991),
    .Y(_3349_));
 sg13g2_or2_1 _4009_ (.X(_3350_),
    .B(_3349_),
    .A(_3347_));
 sg13g2_nand3_1 _4010_ (.B(_3308_),
    .C(_3348_),
    .A(_3307_),
    .Y(_3351_));
 sg13g2_nand2_1 _4011_ (.Y(_3352_),
    .A(_3350_),
    .B(_3351_));
 sg13g2_nand4_1 _4012_ (.B(_3345_),
    .C(_3350_),
    .A(_3343_),
    .Y(_3353_),
    .D(_3351_));
 sg13g2_nor2b_1 _4013_ (.A(net1006),
    .B_N(\vgademo.soundtrack.noise_lfsr[9] ),
    .Y(_3354_));
 sg13g2_a21oi_1 _4014_ (.A1(net1003),
    .A2(\vgademo.soundtrack.noise_lfsr[10] ),
    .Y(_3355_),
    .B1(_3354_));
 sg13g2_mux2_1 _4015_ (.A0(\vgademo.soundtrack.noise_lfsr[11] ),
    .A1(\vgademo.soundtrack.noise_lfsr[12] ),
    .S(net1002),
    .X(_3356_));
 sg13g2_nor2_1 _4016_ (.A(net937),
    .B(_3356_),
    .Y(_3357_));
 sg13g2_a21oi_1 _4017_ (.A1(net937),
    .A2(_3355_),
    .Y(_3358_),
    .B1(_3357_));
 sg13g2_inv_1 _4018_ (.Y(_3359_),
    .A(_3358_));
 sg13g2_nor2_1 _4019_ (.A(net997),
    .B(_3359_),
    .Y(_3360_));
 sg13g2_nor2b_1 _4020_ (.A(net1006),
    .B_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Y(_3361_));
 sg13g2_a21oi_1 _4021_ (.A1(\vgademo.soundtrack.noise_lfsr[6] ),
    .A2(net1005),
    .Y(_3362_),
    .B1(_3361_));
 sg13g2_mux2_1 _4022_ (.A0(\vgademo.soundtrack.noise_lfsr[7] ),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .S(net1005),
    .X(_3363_));
 sg13g2_nor2_1 _4023_ (.A(net938),
    .B(_3363_),
    .Y(_3364_));
 sg13g2_a21oi_1 _4024_ (.A1(net937),
    .A2(_3362_),
    .Y(_3365_),
    .B1(_3364_));
 sg13g2_nand2b_1 _4025_ (.Y(_3366_),
    .B(net997),
    .A_N(_3365_));
 sg13g2_nor2_1 _4026_ (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .B(net1002),
    .Y(_3367_));
 sg13g2_a21oi_1 _4027_ (.A1(net1002),
    .A2(_0040_),
    .Y(_3368_),
    .B1(_3367_));
 sg13g2_a21oi_1 _4028_ (.A1(_3094_),
    .A2(net1002),
    .Y(_3369_),
    .B1(net1000));
 sg13g2_o21ai_1 _4029_ (.B1(_3369_),
    .Y(_3370_),
    .A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(net1002));
 sg13g2_a21oi_1 _4030_ (.A1(net1000),
    .A2(_3368_),
    .Y(_3371_),
    .B1(net996));
 sg13g2_a21oi_1 _4031_ (.A1(_3370_),
    .A2(_3371_),
    .Y(_3372_),
    .B1(net993));
 sg13g2_a22oi_1 _4032_ (.Y(_3373_),
    .B1(_3366_),
    .B2(_3372_),
    .A2(_3360_),
    .A1(net993));
 sg13g2_nor2_1 _4033_ (.A(_3353_),
    .B(_3373_),
    .Y(_3374_));
 sg13g2_nand2_1 _4034_ (.Y(_3375_),
    .A(_3353_),
    .B(_3373_));
 sg13g2_xnor2_1 _4035_ (.Y(_3376_),
    .A(_3353_),
    .B(_3373_));
 sg13g2_xor2_1 _4036_ (.B(\vgademo.soundtrack.tri_osc_p[2] ),
    .A(net987),
    .X(_3377_));
 sg13g2_xor2_1 _4037_ (.B(_3377_),
    .A(_3376_),
    .X(_3378_));
 sg13g2_o21ai_1 _4038_ (.B1(_3333_),
    .Y(_3379_),
    .A1(_3334_),
    .A2(_3336_));
 sg13g2_nor2b_1 _4039_ (.A(_3378_),
    .B_N(_3379_),
    .Y(_3380_));
 sg13g2_xnor2_1 _4040_ (.Y(_3381_),
    .A(_3378_),
    .B(_3379_));
 sg13g2_nand2_1 _4041_ (.Y(_3382_),
    .A(net371),
    .B(_3381_));
 sg13g2_xnor2_1 _4042_ (.Y(_3383_),
    .A(net371),
    .B(_3381_));
 sg13g2_xor2_1 _4043_ (.B(_3383_),
    .A(_3338_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[1] ));
 sg13g2_o21ai_1 _4044_ (.B1(_3382_),
    .Y(_3384_),
    .A1(_3338_),
    .A2(_3383_));
 sg13g2_a21oi_1 _4045_ (.A1(_3375_),
    .A2(_3377_),
    .Y(_3385_),
    .B1(_3374_));
 sg13g2_nand2_1 _4046_ (.Y(_3386_),
    .A(net991),
    .B(_3310_));
 sg13g2_nand4_1 _4047_ (.B(net989),
    .C(_3150_),
    .A(net991),
    .Y(_3387_),
    .D(_3310_));
 sg13g2_nand2_1 _4048_ (.Y(_3388_),
    .A(net937),
    .B(_3315_));
 sg13g2_o21ai_1 _4049_ (.B1(_3388_),
    .Y(_3389_),
    .A1(net938),
    .A2(_3323_));
 sg13g2_or2_1 _4050_ (.X(_3390_),
    .B(_3389_),
    .A(_3153_));
 sg13g2_nor3_1 _4051_ (.A(net1000),
    .B(_3317_),
    .C(_3318_),
    .Y(_3391_));
 sg13g2_o21ai_1 _4052_ (.B1(_3153_),
    .Y(_3392_),
    .A1(net937),
    .A2(_3313_));
 sg13g2_o21ai_1 _4053_ (.B1(_3390_),
    .Y(_3393_),
    .A1(_3391_),
    .A2(_3392_));
 sg13g2_nor2_1 _4054_ (.A(net993),
    .B(_3393_),
    .Y(_3394_));
 sg13g2_nor2_1 _4055_ (.A(net938),
    .B(net1004),
    .Y(_3395_));
 sg13g2_a22oi_1 _4056_ (.Y(_3396_),
    .B1(_3395_),
    .B2(\vgademo.soundtrack.noise_lfsr[12] ),
    .A2(_3320_),
    .A1(net937));
 sg13g2_nor3_1 _4057_ (.A(_3152_),
    .B(net997),
    .C(_3396_),
    .Y(_3397_));
 sg13g2_nor2_1 _4058_ (.A(_3394_),
    .B(_3397_),
    .Y(_3398_));
 sg13g2_or2_1 _4059_ (.X(_0366_),
    .B(_3398_),
    .A(_3387_));
 sg13g2_xnor2_1 _4060_ (.Y(_0367_),
    .A(_3387_),
    .B(_3398_));
 sg13g2_xnor2_1 _4061_ (.Y(_0368_),
    .A(net987),
    .B(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_xnor2_1 _4062_ (.Y(_0369_),
    .A(_0367_),
    .B(_0368_));
 sg13g2_nor2_1 _4063_ (.A(_3385_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_xor2_1 _4064_ (.B(_0369_),
    .A(_3385_),
    .X(_0371_));
 sg13g2_xor2_1 _4065_ (.B(_0371_),
    .A(_3380_),
    .X(_0372_));
 sg13g2_and2_1 _4066_ (.A(net566),
    .B(_0372_),
    .X(_0373_));
 sg13g2_or2_1 _4067_ (.X(_0374_),
    .B(_0372_),
    .A(net566));
 sg13g2_nand2b_1 _4068_ (.Y(_0375_),
    .B(_0374_),
    .A_N(_0373_));
 sg13g2_xnor2_1 _4069_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .A(_3384_),
    .B(_0375_));
 sg13g2_a21oi_1 _4070_ (.A1(_3384_),
    .A2(_0374_),
    .Y(_0376_),
    .B1(_0373_));
 sg13g2_a21oi_1 _4071_ (.A1(_3380_),
    .A2(_0371_),
    .Y(_0377_),
    .B1(_0370_));
 sg13g2_o21ai_1 _4072_ (.B1(_0366_),
    .Y(_0378_),
    .A1(_0367_),
    .A2(_0368_));
 sg13g2_nor3_1 _4073_ (.A(\vgademo.soundtrack.pulse_vol[2] ),
    .B(_3347_),
    .C(_3349_),
    .Y(_0379_));
 sg13g2_o21ai_1 _4074_ (.B1(_0379_),
    .Y(_0380_),
    .A1(net992),
    .A2(_3309_));
 sg13g2_or2_1 _4075_ (.X(_0381_),
    .B(_0380_),
    .A(_3342_));
 sg13g2_nor2_1 _4076_ (.A(net1001),
    .B(_3363_),
    .Y(_0382_));
 sg13g2_a21oi_1 _4077_ (.A1(net1001),
    .A2(_3355_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_nand2b_1 _4078_ (.Y(_0384_),
    .B(net1001),
    .A_N(_3362_));
 sg13g2_a21oi_1 _4079_ (.A1(net937),
    .A2(_3368_),
    .Y(_0385_),
    .B1(net996));
 sg13g2_a21oi_1 _4080_ (.A1(_0384_),
    .A2(_0385_),
    .Y(_0386_),
    .B1(net993));
 sg13g2_o21ai_1 _4081_ (.B1(_0386_),
    .Y(_0387_),
    .A1(_3153_),
    .A2(_0383_));
 sg13g2_nand2_1 _4082_ (.Y(_0388_),
    .A(net939),
    .B(_3356_));
 sg13g2_nand3_1 _4083_ (.B(_3153_),
    .C(_3356_),
    .A(net939),
    .Y(_0389_));
 sg13g2_o21ai_1 _4084_ (.B1(_0387_),
    .Y(_0390_),
    .A1(_3152_),
    .A2(_0389_));
 sg13g2_nand2b_1 _4085_ (.Y(_0391_),
    .B(_0390_),
    .A_N(_0381_));
 sg13g2_xor2_1 _4086_ (.B(_0390_),
    .A(_0381_),
    .X(_0392_));
 sg13g2_xor2_1 _4087_ (.B(\vgademo.soundtrack.tri_osc_p[4] ),
    .A(net987),
    .X(_0393_));
 sg13g2_inv_1 _4088_ (.Y(_0394_),
    .A(_0393_));
 sg13g2_xnor2_1 _4089_ (.Y(_0395_),
    .A(_0392_),
    .B(_0394_));
 sg13g2_nand2b_1 _4090_ (.Y(_0396_),
    .B(_0378_),
    .A_N(_0395_));
 sg13g2_xor2_1 _4091_ (.B(_0395_),
    .A(_0378_),
    .X(_0397_));
 sg13g2_xor2_1 _4092_ (.B(_0397_),
    .A(_0377_),
    .X(_0398_));
 sg13g2_nand2_1 _4093_ (.Y(_0399_),
    .A(net532),
    .B(_0398_));
 sg13g2_xnor2_1 _4094_ (.Y(_0400_),
    .A(net532),
    .B(_0398_));
 sg13g2_xor2_1 _4095_ (.B(_0400_),
    .A(_0376_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[3] ));
 sg13g2_o21ai_1 _4096_ (.B1(_0399_),
    .Y(_0401_),
    .A1(_0376_),
    .A2(_0400_));
 sg13g2_o21ai_1 _4097_ (.B1(_0396_),
    .Y(_0402_),
    .A1(_0377_),
    .A2(_0397_));
 sg13g2_o21ai_1 _4098_ (.B1(_0391_),
    .Y(_0403_),
    .A1(_0392_),
    .A2(_0394_));
 sg13g2_nand2_1 _4099_ (.Y(_0404_),
    .A(_3310_),
    .B(_3344_));
 sg13g2_nand3_1 _4100_ (.B(_3310_),
    .C(_3344_),
    .A(net989),
    .Y(_0405_));
 sg13g2_or2_1 _4101_ (.X(_0406_),
    .B(_3316_),
    .A(net996));
 sg13g2_a21oi_1 _4102_ (.A1(net996),
    .A2(_3324_),
    .Y(_0407_),
    .B1(net993));
 sg13g2_nand2b_1 _4103_ (.Y(_0408_),
    .B(_3153_),
    .A_N(_3326_));
 sg13g2_a22oi_1 _4104_ (.Y(_0409_),
    .B1(_0408_),
    .B2(net994),
    .A2(_0407_),
    .A1(_0406_));
 sg13g2_nor2b_1 _4105_ (.A(_0405_),
    .B_N(_0409_),
    .Y(_0410_));
 sg13g2_xnor2_1 _4106_ (.Y(_0411_),
    .A(_0405_),
    .B(_0409_));
 sg13g2_xor2_1 _4107_ (.B(\vgademo.soundtrack.tri_osc_p[5] ),
    .A(net988),
    .X(_0412_));
 sg13g2_xor2_1 _4108_ (.B(_0412_),
    .A(_0411_),
    .X(_0413_));
 sg13g2_xnor2_1 _4109_ (.Y(_0414_),
    .A(_0403_),
    .B(_0413_));
 sg13g2_nor2b_1 _4110_ (.A(_0414_),
    .B_N(_0402_),
    .Y(_0415_));
 sg13g2_xnor2_1 _4111_ (.Y(_0416_),
    .A(_0402_),
    .B(_0414_));
 sg13g2_and2_1 _4112_ (.A(net565),
    .B(_0416_),
    .X(_0417_));
 sg13g2_or2_1 _4113_ (.X(_0418_),
    .B(_0416_),
    .A(net565));
 sg13g2_nand2b_1 _4114_ (.Y(_0419_),
    .B(_0418_),
    .A_N(_0417_));
 sg13g2_xnor2_1 _4115_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .A(_0401_),
    .B(_0419_));
 sg13g2_a21oi_1 _4116_ (.A1(_0401_),
    .A2(_0418_),
    .Y(_0420_),
    .B1(_0417_));
 sg13g2_a21oi_1 _4117_ (.A1(_0403_),
    .A2(_0413_),
    .Y(_0421_),
    .B1(_0415_));
 sg13g2_a21o_1 _4118_ (.A2(_0412_),
    .A1(_0411_),
    .B1(_0410_),
    .X(_0422_));
 sg13g2_a21oi_1 _4119_ (.A1(net997),
    .A2(_3359_),
    .Y(_0423_),
    .B1(net993));
 sg13g2_o21ai_1 _4120_ (.B1(_0423_),
    .Y(_0424_),
    .A1(net999),
    .A2(_3365_));
 sg13g2_nand4_1 _4121_ (.B(_3346_),
    .C(_3350_),
    .A(_3343_),
    .Y(_0425_),
    .D(_3351_));
 sg13g2_nor2_1 _4122_ (.A(_0424_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_xor2_1 _4123_ (.B(_0425_),
    .A(_0424_),
    .X(_0427_));
 sg13g2_xnor2_1 _4124_ (.Y(_0428_),
    .A(\vgademo.soundtrack.tri_osc_p[15] ),
    .B(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_inv_1 _4125_ (.Y(_0429_),
    .A(_0428_));
 sg13g2_xnor2_1 _4126_ (.Y(_0430_),
    .A(_0427_),
    .B(_0428_));
 sg13g2_nand2_1 _4127_ (.Y(_0431_),
    .A(_0422_),
    .B(_0430_));
 sg13g2_xnor2_1 _4128_ (.Y(_0432_),
    .A(_0422_),
    .B(_0430_));
 sg13g2_xor2_1 _4129_ (.B(_0432_),
    .A(_0421_),
    .X(_0433_));
 sg13g2_nand2_1 _4130_ (.Y(_0434_),
    .A(net519),
    .B(_0433_));
 sg13g2_xnor2_1 _4131_ (.Y(_0435_),
    .A(net519),
    .B(_0433_));
 sg13g2_xor2_1 _4132_ (.B(_0435_),
    .A(_0420_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[5] ));
 sg13g2_o21ai_1 _4133_ (.B1(_0434_),
    .Y(_0436_),
    .A1(_0420_),
    .A2(_0435_));
 sg13g2_o21ai_1 _4134_ (.B1(_0431_),
    .Y(_0437_),
    .A1(_0421_),
    .A2(_0432_));
 sg13g2_a21oi_1 _4135_ (.A1(_0427_),
    .A2(_0429_),
    .Y(_0438_),
    .B1(_0426_));
 sg13g2_a21oi_1 _4136_ (.A1(net997),
    .A2(_3396_),
    .Y(_0439_),
    .B1(net994));
 sg13g2_o21ai_1 _4137_ (.B1(_0439_),
    .Y(_0440_),
    .A1(net997),
    .A2(_3389_));
 sg13g2_nor2_1 _4138_ (.A(net989),
    .B(_3339_),
    .Y(_0441_));
 sg13g2_nand2_1 _4139_ (.Y(_0442_),
    .A(_3310_),
    .B(_0441_));
 sg13g2_xor2_1 _4140_ (.B(_0442_),
    .A(_0440_),
    .X(_0443_));
 sg13g2_xnor2_1 _4141_ (.Y(_0444_),
    .A(net988),
    .B(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_nand2b_1 _4142_ (.Y(_0445_),
    .B(_0443_),
    .A_N(_0444_));
 sg13g2_xor2_1 _4143_ (.B(_0444_),
    .A(_0443_),
    .X(_0446_));
 sg13g2_nor2_1 _4144_ (.A(_0438_),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_xor2_1 _4145_ (.B(_0446_),
    .A(_0438_),
    .X(_0448_));
 sg13g2_xor2_1 _4146_ (.B(_0448_),
    .A(_0437_),
    .X(_0449_));
 sg13g2_and2_1 _4147_ (.A(net563),
    .B(_0449_),
    .X(_0450_));
 sg13g2_or2_1 _4148_ (.X(_0451_),
    .B(_0449_),
    .A(net563));
 sg13g2_nand2b_1 _4149_ (.Y(_0452_),
    .B(_0451_),
    .A_N(_0450_));
 sg13g2_xnor2_1 _4150_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[6] ),
    .A(_0436_),
    .B(_0452_));
 sg13g2_a21oi_1 _4151_ (.A1(_0436_),
    .A2(_0451_),
    .Y(_0453_),
    .B1(_0450_));
 sg13g2_a21oi_1 _4152_ (.A1(_0437_),
    .A2(_0448_),
    .Y(_0454_),
    .B1(_0447_));
 sg13g2_o21ai_1 _4153_ (.B1(_0445_),
    .Y(_0455_),
    .A1(_0440_),
    .A2(_0442_));
 sg13g2_o21ai_1 _4154_ (.B1(_3152_),
    .Y(_0456_),
    .A1(net997),
    .A2(_0383_));
 sg13g2_a21oi_2 _4155_ (.B1(_0456_),
    .Y(_0457_),
    .A2(_0388_),
    .A1(net997));
 sg13g2_nor3_1 _4156_ (.A(net991),
    .B(net989),
    .C(_3150_),
    .Y(_0458_));
 sg13g2_nor3_1 _4157_ (.A(net992),
    .B(net989),
    .C(_3339_),
    .Y(_0459_));
 sg13g2_a22oi_1 _4158_ (.Y(_0460_),
    .B1(_0459_),
    .B2(_3309_),
    .A2(_0458_),
    .A1(net992));
 sg13g2_nand2b_1 _4159_ (.Y(_0461_),
    .B(_0457_),
    .A_N(_0460_));
 sg13g2_xnor2_1 _4160_ (.Y(_0462_),
    .A(_0457_),
    .B(_0460_));
 sg13g2_inv_1 _4161_ (.Y(_0463_),
    .A(_0462_));
 sg13g2_xnor2_1 _4162_ (.Y(_0464_),
    .A(net988),
    .B(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_xnor2_1 _4163_ (.Y(_0465_),
    .A(_0462_),
    .B(_0464_));
 sg13g2_nand2_1 _4164_ (.Y(_0466_),
    .A(_0455_),
    .B(_0465_));
 sg13g2_xnor2_1 _4165_ (.Y(_0467_),
    .A(_0455_),
    .B(_0465_));
 sg13g2_xor2_1 _4166_ (.B(_0467_),
    .A(_0454_),
    .X(_0468_));
 sg13g2_nand2_1 _4167_ (.Y(_0469_),
    .A(\vgademo.soundtrack.sigma_delta_accum[7] ),
    .B(_0468_));
 sg13g2_xnor2_1 _4168_ (.Y(_0470_),
    .A(net516),
    .B(_0468_));
 sg13g2_xor2_1 _4169_ (.B(_0470_),
    .A(_0453_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[7] ));
 sg13g2_o21ai_1 _4170_ (.B1(_0469_),
    .Y(_0471_),
    .A1(_0453_),
    .A2(_0470_));
 sg13g2_o21ai_1 _4171_ (.B1(_0466_),
    .Y(_0472_),
    .A1(_0454_),
    .A2(_0467_));
 sg13g2_o21ai_1 _4172_ (.B1(_0461_),
    .Y(_0473_),
    .A1(_0463_),
    .A2(_0464_));
 sg13g2_inv_1 _4173_ (.Y(_0474_),
    .A(_0473_));
 sg13g2_and2_1 _4174_ (.A(_3152_),
    .B(_3327_),
    .X(_0475_));
 sg13g2_and2_1 _4175_ (.A(_3310_),
    .B(_0458_),
    .X(_0476_));
 sg13g2_nand2_1 _4176_ (.Y(_0477_),
    .A(_0475_),
    .B(_0476_));
 sg13g2_xnor2_1 _4177_ (.Y(_0478_),
    .A(_0475_),
    .B(_0476_));
 sg13g2_xnor2_1 _4178_ (.Y(_0479_),
    .A(net988),
    .B(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_xnor2_1 _4179_ (.Y(_0480_),
    .A(_0478_),
    .B(_0479_));
 sg13g2_xor2_1 _4180_ (.B(_0480_),
    .A(_0473_),
    .X(_0481_));
 sg13g2_nand2b_1 _4181_ (.Y(_0482_),
    .B(_0472_),
    .A_N(_0481_));
 sg13g2_xnor2_1 _4182_ (.Y(_0483_),
    .A(_0472_),
    .B(_0481_));
 sg13g2_xnor2_1 _4183_ (.Y(_0484_),
    .A(net511),
    .B(_0483_));
 sg13g2_nor2b_1 _4184_ (.A(_0484_),
    .B_N(_0471_),
    .Y(_0485_));
 sg13g2_xnor2_1 _4185_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[8] ),
    .A(_0471_),
    .B(_0484_));
 sg13g2_a21o_1 _4186_ (.A2(_0483_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[8] ),
    .B1(_0485_),
    .X(_0486_));
 sg13g2_o21ai_1 _4187_ (.B1(_0482_),
    .Y(_0487_),
    .A1(_0474_),
    .A2(_0480_));
 sg13g2_o21ai_1 _4188_ (.B1(_0477_),
    .Y(_0488_),
    .A1(_0478_),
    .A2(_0479_));
 sg13g2_nand2_1 _4189_ (.Y(_0489_),
    .A(_3152_),
    .B(_3360_));
 sg13g2_or3_1 _4190_ (.A(net990),
    .B(_3346_),
    .C(_3352_),
    .X(_0490_));
 sg13g2_nor2_1 _4191_ (.A(_0489_),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_xor2_1 _4192_ (.B(_0490_),
    .A(_0489_),
    .X(_0492_));
 sg13g2_xnor2_1 _4193_ (.Y(_0493_),
    .A(net988),
    .B(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_inv_1 _4194_ (.Y(_0494_),
    .A(_0493_));
 sg13g2_xnor2_1 _4195_ (.Y(_0495_),
    .A(_0492_),
    .B(_0493_));
 sg13g2_xnor2_1 _4196_ (.Y(_0496_),
    .A(_0488_),
    .B(_0495_));
 sg13g2_nor2b_1 _4197_ (.A(_0496_),
    .B_N(_0487_),
    .Y(_0497_));
 sg13g2_xnor2_1 _4198_ (.Y(_0498_),
    .A(_0487_),
    .B(_0496_));
 sg13g2_xnor2_1 _4199_ (.Y(_0499_),
    .A(net501),
    .B(_0498_));
 sg13g2_nor2b_1 _4200_ (.A(_0499_),
    .B_N(_0486_),
    .Y(_0500_));
 sg13g2_xnor2_1 _4201_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .A(_0486_),
    .B(_0499_));
 sg13g2_a21o_1 _4202_ (.A2(_0498_),
    .A1(net501),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_a21o_1 _4203_ (.A2(_0495_),
    .A1(_0488_),
    .B1(_0497_),
    .X(_0502_));
 sg13g2_a21oi_1 _4204_ (.A1(_0492_),
    .A2(_0494_),
    .Y(_0503_),
    .B1(_0491_));
 sg13g2_nor3_1 _4205_ (.A(net995),
    .B(net999),
    .C(_3396_),
    .Y(_0504_));
 sg13g2_nor3_1 _4206_ (.A(net989),
    .B(\vgademo.soundtrack.pulse_vol[2] ),
    .C(_3386_),
    .Y(_0505_));
 sg13g2_nand2_1 _4207_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_xnor2_1 _4208_ (.Y(_0507_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_xor2_1 _4209_ (.B(\vgademo.soundtrack.tri_osc_p[11] ),
    .A(net988),
    .X(_0508_));
 sg13g2_inv_1 _4210_ (.Y(_0509_),
    .A(_0508_));
 sg13g2_xnor2_1 _4211_ (.Y(_0510_),
    .A(_0507_),
    .B(_0509_));
 sg13g2_nor2_1 _4212_ (.A(_0503_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_xor2_1 _4213_ (.B(_0510_),
    .A(_0503_),
    .X(_0512_));
 sg13g2_xor2_1 _4214_ (.B(_0512_),
    .A(_0502_),
    .X(_0513_));
 sg13g2_xnor2_1 _4215_ (.Y(_0514_),
    .A(net507),
    .B(_0513_));
 sg13g2_nor2b_1 _4216_ (.A(_0514_),
    .B_N(_0501_),
    .Y(_0515_));
 sg13g2_xnor2_1 _4217_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .A(_0501_),
    .B(_0514_));
 sg13g2_a21o_1 _4218_ (.A2(_0513_),
    .A1(net507),
    .B1(_0515_),
    .X(_0516_));
 sg13g2_a21oi_1 _4219_ (.A1(_0502_),
    .A2(_0512_),
    .Y(_0517_),
    .B1(_0511_));
 sg13g2_o21ai_1 _4220_ (.B1(_0506_),
    .Y(_0518_),
    .A1(_0507_),
    .A2(_0509_));
 sg13g2_nand2b_1 _4221_ (.Y(_0519_),
    .B(_3342_),
    .A_N(_0380_));
 sg13g2_nor3_1 _4222_ (.A(net995),
    .B(_0389_),
    .C(_0519_),
    .Y(_0520_));
 sg13g2_o21ai_1 _4223_ (.B1(_0519_),
    .Y(_0521_),
    .A1(net995),
    .A2(_0389_));
 sg13g2_nor2b_1 _4224_ (.A(_0520_),
    .B_N(_0521_),
    .Y(_0522_));
 sg13g2_xor2_1 _4225_ (.B(\vgademo.soundtrack.tri_osc_p[12] ),
    .A(net988),
    .X(_0523_));
 sg13g2_xor2_1 _4226_ (.B(_0523_),
    .A(_0522_),
    .X(_0524_));
 sg13g2_nand2_1 _4227_ (.Y(_0525_),
    .A(_0518_),
    .B(_0524_));
 sg13g2_xnor2_1 _4228_ (.Y(_0526_),
    .A(_0518_),
    .B(_0524_));
 sg13g2_xor2_1 _4229_ (.B(_0526_),
    .A(_0517_),
    .X(_0527_));
 sg13g2_xnor2_1 _4230_ (.Y(_0528_),
    .A(net524),
    .B(_0527_));
 sg13g2_nor2b_1 _4231_ (.A(_0528_),
    .B_N(_0516_),
    .Y(_0529_));
 sg13g2_xnor2_1 _4232_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .A(_0516_),
    .B(_0528_));
 sg13g2_a21o_1 _4233_ (.A2(_0527_),
    .A1(net524),
    .B1(_0529_),
    .X(_0530_));
 sg13g2_o21ai_1 _4234_ (.B1(_0525_),
    .Y(_0531_),
    .A1(_0517_),
    .A2(_0526_));
 sg13g2_a21o_1 _4235_ (.A2(_0523_),
    .A1(_0522_),
    .B1(_0520_),
    .X(_0532_));
 sg13g2_nor2_2 _4236_ (.A(net993),
    .B(_0408_),
    .Y(_0533_));
 sg13g2_nor2_1 _4237_ (.A(net990),
    .B(_0404_),
    .Y(_0534_));
 sg13g2_nand2_1 _4238_ (.Y(_0535_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_xnor2_1 _4239_ (.Y(_0536_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_xnor2_1 _4240_ (.Y(_0537_),
    .A(net987),
    .B(\vgademo.soundtrack.tri_osc_p[13] ));
 sg13g2_xor2_1 _4241_ (.B(_0537_),
    .A(_0536_),
    .X(_0538_));
 sg13g2_xnor2_1 _4242_ (.Y(_0539_),
    .A(_0532_),
    .B(_0538_));
 sg13g2_nor2b_1 _4243_ (.A(_0539_),
    .B_N(_0531_),
    .Y(_0540_));
 sg13g2_xnor2_1 _4244_ (.Y(_0541_),
    .A(_0531_),
    .B(_0539_));
 sg13g2_xnor2_1 _4245_ (.Y(_0542_),
    .A(net526),
    .B(_0541_));
 sg13g2_nor2b_1 _4246_ (.A(_0542_),
    .B_N(_0530_),
    .Y(_0543_));
 sg13g2_xnor2_1 _4247_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .A(_0530_),
    .B(_0542_));
 sg13g2_a21o_1 _4248_ (.A2(_0541_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[12] ),
    .B1(_0543_),
    .X(_0544_));
 sg13g2_o21ai_1 _4249_ (.B1(_0535_),
    .Y(_0545_),
    .A1(_0536_),
    .A2(_0537_));
 sg13g2_nor4_2 _4250_ (.A(net991),
    .B(net990),
    .C(\vgademo.soundtrack.pulse_vol[2] ),
    .Y(_0546_),
    .D(_3352_));
 sg13g2_nand2b_1 _4251_ (.Y(_0547_),
    .B(net368),
    .A_N(net987));
 sg13g2_xnor2_1 _4252_ (.Y(_0548_),
    .A(\vgademo.soundtrack.tri_osc_p[14] ),
    .B(net987));
 sg13g2_nand2b_1 _4253_ (.Y(_0549_),
    .B(_0548_),
    .A_N(_0546_));
 sg13g2_xor2_1 _4254_ (.B(_0548_),
    .A(_0546_),
    .X(_0550_));
 sg13g2_and2_1 _4255_ (.A(_0545_),
    .B(_0550_),
    .X(_0551_));
 sg13g2_xor2_1 _4256_ (.B(_0550_),
    .A(_0545_),
    .X(_0552_));
 sg13g2_a21o_1 _4257_ (.A2(_0538_),
    .A1(_0532_),
    .B1(_0540_),
    .X(_0553_));
 sg13g2_xor2_1 _4258_ (.B(_0553_),
    .A(_0552_),
    .X(_0554_));
 sg13g2_xnor2_1 _4259_ (.Y(_0555_),
    .A(net513),
    .B(_0554_));
 sg13g2_nor2b_1 _4260_ (.A(_0555_),
    .B_N(_0544_),
    .Y(_0556_));
 sg13g2_xnor2_1 _4261_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .A(_0544_),
    .B(_0555_));
 sg13g2_a21o_1 _4262_ (.A2(_0554_),
    .A1(net513),
    .B1(_0556_),
    .X(_0557_));
 sg13g2_a21oi_1 _4263_ (.A1(_0552_),
    .A2(_0553_),
    .Y(_0558_),
    .B1(_0551_));
 sg13g2_nor3_2 _4264_ (.A(_0545_),
    .B(_0549_),
    .C(_0553_),
    .Y(_0559_));
 sg13g2_xor2_1 _4265_ (.B(_0558_),
    .A(_0549_),
    .X(_0560_));
 sg13g2_and2_1 _4266_ (.A(net549),
    .B(_0560_),
    .X(_0561_));
 sg13g2_xor2_1 _4267_ (.B(_0560_),
    .A(net549),
    .X(_0562_));
 sg13g2_xor2_1 _4268_ (.B(_0562_),
    .A(_0557_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[14] ));
 sg13g2_a21o_1 _4269_ (.A2(_0562_),
    .A1(_0557_),
    .B1(_0561_),
    .X(_0563_));
 sg13g2_nor2b_1 _4270_ (.A(_0559_),
    .B_N(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .Y(_0564_));
 sg13g2_xnor2_1 _4271_ (.Y(_0565_),
    .A(net554),
    .B(_0559_));
 sg13g2_xor2_1 _4272_ (.B(_0565_),
    .A(_0563_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[15] ));
 sg13g2_xor2_1 _4273_ (.B(net254),
    .A(\vgademo.soundtrack.sample_div[1] ),
    .X(\vgademo.soundtrack.sample_div_[1] ));
 sg13g2_nand3_1 _4274_ (.B(\vgademo.soundtrack.sample_div[1] ),
    .C(net254),
    .A(net453),
    .Y(_0566_));
 sg13g2_a21o_1 _4275_ (.A2(net254),
    .A1(\vgademo.soundtrack.sample_div[1] ),
    .B1(net453),
    .X(_0567_));
 sg13g2_and2_1 _4276_ (.A(_0566_),
    .B(net454),
    .X(\vgademo.soundtrack.sample_div_[2] ));
 sg13g2_nor2_1 _4277_ (.A(_3104_),
    .B(_0566_),
    .Y(_0568_));
 sg13g2_xnor2_1 _4278_ (.Y(\vgademo.soundtrack.sample_div_[3] ),
    .A(net244),
    .B(_0566_));
 sg13g2_and2_1 _4279_ (.A(net228),
    .B(_0568_),
    .X(_0569_));
 sg13g2_xor2_1 _4280_ (.B(_0568_),
    .A(net228),
    .X(\vgademo.soundtrack.sample_div_[4] ));
 sg13g2_xor2_1 _4281_ (.B(_0569_),
    .A(net270),
    .X(\vgademo.soundtrack.sample_div_[5] ));
 sg13g2_nand3_1 _4282_ (.B(net270),
    .C(_0569_),
    .A(net456),
    .Y(_0570_));
 sg13g2_a21o_1 _4283_ (.A2(_0569_),
    .A1(net270),
    .B1(net456),
    .X(_0571_));
 sg13g2_and2_1 _4284_ (.A(_0570_),
    .B(_0571_),
    .X(\vgademo.soundtrack.sample_div_[6] ));
 sg13g2_nor2_1 _4285_ (.A(_3103_),
    .B(_0570_),
    .Y(_0572_));
 sg13g2_xnor2_1 _4286_ (.Y(\vgademo.soundtrack.sample_div_[7] ),
    .A(net230),
    .B(_0570_));
 sg13g2_and2_1 _4287_ (.A(net211),
    .B(_0572_),
    .X(_0573_));
 sg13g2_xor2_1 _4288_ (.B(_0572_),
    .A(net211),
    .X(\vgademo.soundtrack.sample_div_[8] ));
 sg13g2_and2_1 _4289_ (.A(\vgademo.soundtrack.sample_div[9] ),
    .B(_0573_),
    .X(_0574_));
 sg13g2_nand2_1 _4290_ (.Y(_0575_),
    .A(\vgademo.soundtrack.sample_div[9] ),
    .B(_0573_));
 sg13g2_xor2_1 _4291_ (.B(_0573_),
    .A(net268),
    .X(\vgademo.soundtrack.sample_div_[9] ));
 sg13g2_nor4_2 _4292_ (.A(\vgademo.h_count[4] ),
    .B(\vgademo.h_count[5] ),
    .C(_3210_),
    .Y(_0576_),
    .D(_3213_));
 sg13g2_nor2_1 _4293_ (.A(\vgademo.h_count[9] ),
    .B(net983),
    .Y(_0577_));
 sg13g2_nor3_2 _4294_ (.A(\vgademo.h_count[9] ),
    .B(net983),
    .C(net982),
    .Y(_0578_));
 sg13g2_and2_1 _4295_ (.A(_0576_),
    .B(_0578_),
    .X(_0579_));
 sg13g2_nand2_2 _4296_ (.Y(_0580_),
    .A(_0576_),
    .B(_0578_));
 sg13g2_and2_1 _4297_ (.A(net1067),
    .B(_3216_),
    .X(_0581_));
 sg13g2_nand2_1 _4298_ (.Y(_0582_),
    .A(net1067),
    .B(_3216_));
 sg13g2_nor2_1 _4299_ (.A(net893),
    .B(net923),
    .Y(_0583_));
 sg13g2_nor3_1 _4300_ (.A(\vgademo.v_count[7] ),
    .B(net958),
    .C(\vgademo.v_count[8] ),
    .Y(_0584_));
 sg13g2_nand2_1 _4301_ (.Y(_0585_),
    .A(net955),
    .B(_0584_));
 sg13g2_nor3_1 _4302_ (.A(net960),
    .B(net959),
    .C(_3243_),
    .Y(_0586_));
 sg13g2_nand4_1 _4303_ (.B(_3244_),
    .C(_0584_),
    .A(net955),
    .Y(_0587_),
    .D(_0586_));
 sg13g2_nor2_1 _4304_ (.A(net930),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_or2_1 _4305_ (.X(_0589_),
    .B(_0587_),
    .A(net930));
 sg13g2_nor3_1 _4306_ (.A(net960),
    .B(_3243_),
    .C(_0585_),
    .Y(_0590_));
 sg13g2_and4_2 _4307_ (.A(_3118_),
    .B(_3217_),
    .C(_3244_),
    .D(_0590_),
    .X(_0591_));
 sg13g2_a21oi_2 _4308_ (.B1(net885),
    .Y(_0592_),
    .A2(_0591_),
    .A1(net1066));
 sg13g2_nor2_1 _4309_ (.A(_3197_),
    .B(net866),
    .Y(_0593_));
 sg13g2_nor2_1 _4310_ (.A(net1041),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_nor2_1 _4311_ (.A(net1039),
    .B(net898),
    .Y(_0595_));
 sg13g2_nor2_1 _4312_ (.A(net1041),
    .B(net898),
    .Y(_0596_));
 sg13g2_nor3_1 _4313_ (.A(net865),
    .B(_0595_),
    .C(_0596_),
    .Y(_0597_));
 sg13g2_nor2_1 _4314_ (.A(_0594_),
    .B(_0597_),
    .Y(_0112_));
 sg13g2_nor3_1 _4315_ (.A(net547),
    .B(net898),
    .C(net868),
    .Y(_0598_));
 sg13g2_a21oi_1 _4316_ (.A1(_3197_),
    .A2(net867),
    .Y(_0113_),
    .B1(_0598_));
 sg13g2_nand2_1 _4317_ (.Y(_0599_),
    .A(\vgademo.linelfsr[2] ),
    .B(net868));
 sg13g2_nand2_1 _4318_ (.Y(_0600_),
    .A(net388),
    .B(net902));
 sg13g2_o21ai_1 _4319_ (.B1(_0599_),
    .Y(_0114_),
    .A1(net868),
    .A2(_0600_));
 sg13g2_xnor2_1 _4320_ (.Y(_0601_),
    .A(net1042),
    .B(net398));
 sg13g2_a21oi_1 _4321_ (.A1(net902),
    .A2(_0601_),
    .Y(_0602_),
    .B1(net868));
 sg13g2_a21o_1 _4322_ (.A2(net867),
    .A1(net388),
    .B1(_0602_),
    .X(_0115_));
 sg13g2_xnor2_1 _4323_ (.Y(_0603_),
    .A(net1042),
    .B(net392));
 sg13g2_a21oi_1 _4324_ (.A1(net902),
    .A2(_0603_),
    .Y(_0604_),
    .B1(net867));
 sg13g2_a21o_1 _4325_ (.A2(net867),
    .A1(net398),
    .B1(_0604_),
    .X(_0116_));
 sg13g2_nor3_1 _4326_ (.A(\vgademo.linelfsr[6] ),
    .B(net898),
    .C(net867),
    .Y(_0605_));
 sg13g2_a21oi_1 _4327_ (.A1(_3198_),
    .A2(net867),
    .Y(_0117_),
    .B1(_0605_));
 sg13g2_xnor2_1 _4328_ (.Y(_0606_),
    .A(net1042),
    .B(net375));
 sg13g2_a21oi_1 _4329_ (.A1(net902),
    .A2(_0606_),
    .Y(_0607_),
    .B1(net867));
 sg13g2_a21o_1 _4330_ (.A2(net867),
    .A1(net442),
    .B1(_0607_),
    .X(_0118_));
 sg13g2_nor3_1 _4331_ (.A(\vgademo.linelfsr[8] ),
    .B(net898),
    .C(net866),
    .Y(_0608_));
 sg13g2_a21oi_1 _4332_ (.A1(_3199_),
    .A2(net866),
    .Y(_0119_),
    .B1(_0608_));
 sg13g2_xnor2_1 _4333_ (.Y(_0609_),
    .A(net1041),
    .B(net370));
 sg13g2_nor3_1 _4334_ (.A(net898),
    .B(net866),
    .C(_0609_),
    .Y(_0610_));
 sg13g2_a21o_1 _4335_ (.A2(net866),
    .A1(net384),
    .B1(_0610_),
    .X(_0120_));
 sg13g2_nor3_1 _4336_ (.A(net320),
    .B(net898),
    .C(net866),
    .Y(_0611_));
 sg13g2_a21oi_1 _4337_ (.A1(_3200_),
    .A2(net865),
    .Y(_0121_),
    .B1(_0611_));
 sg13g2_nand2_1 _4338_ (.Y(_0612_),
    .A(net320),
    .B(net865));
 sg13g2_nand2_1 _4339_ (.Y(_0613_),
    .A(\vgademo.linelfsr[11] ),
    .B(net902));
 sg13g2_o21ai_1 _4340_ (.B1(_0612_),
    .Y(_0122_),
    .A1(net865),
    .A2(_0613_));
 sg13g2_nor3_1 _4341_ (.A(\vgademo.linelfsr[12] ),
    .B(net898),
    .C(net865),
    .Y(_0614_));
 sg13g2_a21oi_1 _4342_ (.A1(_3101_),
    .A2(net865),
    .Y(_0123_),
    .B1(_0614_));
 sg13g2_nand2_1 _4343_ (.Y(_0615_),
    .A(net338),
    .B(net865));
 sg13g2_o21ai_1 _4344_ (.B1(_0615_),
    .Y(_0124_),
    .A1(net865),
    .A2(_0596_));
 sg13g2_nand3_1 _4345_ (.B(net496),
    .C(net872),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0616_));
 sg13g2_nand4_1 _4346_ (.B(net242),
    .C(\vgademo.soundtrack.tick_div[1] ),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0617_),
    .D(net872));
 sg13g2_nor2_1 _4347_ (.A(_3105_),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_and2_1 _4348_ (.A(net213),
    .B(_0618_),
    .X(_0619_));
 sg13g2_and3_2 _4349_ (.X(_0620_),
    .A(net206),
    .B(net276),
    .C(_0619_));
 sg13g2_and2_2 _4350_ (.A(net290),
    .B(_0620_),
    .X(_0621_));
 sg13g2_nand2_2 _4351_ (.Y(_0622_),
    .A(net290),
    .B(_0620_));
 sg13g2_or2_1 _4352_ (.X(_0623_),
    .B(\vgademo.audio_beat_out[0] ),
    .A(\vgademo.audio_beat_out[1] ));
 sg13g2_nor4_2 _4353_ (.A(\vgademo.audio_beat_out[3] ),
    .B(\vgademo.audio_beat_out[2] ),
    .C(net590),
    .Y(_0624_),
    .D(_0623_));
 sg13g2_or4_2 _4354_ (.A(\vgademo.audio_beat_out[3] ),
    .B(\vgademo.audio_beat_out[2] ),
    .C(\vgademo.audio_beat_out[4] ),
    .D(_0623_),
    .X(_0625_));
 sg13g2_nand2_1 _4355_ (.Y(_0626_),
    .A(_0621_),
    .B(net934));
 sg13g2_nor2_1 _4356_ (.A(net1038),
    .B(net846),
    .Y(_0627_));
 sg13g2_a21oi_1 _4357_ (.A1(_3100_),
    .A2(net846),
    .Y(_0125_),
    .B1(_0627_));
 sg13g2_nand2_1 _4358_ (.Y(_0628_),
    .A(net189),
    .B(net844));
 sg13g2_o21ai_1 _4359_ (.B1(_0628_),
    .Y(_0126_),
    .A1(_3281_),
    .A2(net844));
 sg13g2_nand2_1 _4360_ (.Y(_0629_),
    .A(net1037),
    .B(net1033));
 sg13g2_xnor2_1 _4361_ (.Y(_0630_),
    .A(net1030),
    .B(_3279_));
 sg13g2_nand2_1 _4362_ (.Y(_0631_),
    .A(net188),
    .B(net844));
 sg13g2_o21ai_1 _4363_ (.B1(_0631_),
    .Y(_0127_),
    .A1(net844),
    .A2(_0630_));
 sg13g2_nor2_1 _4364_ (.A(_3279_),
    .B(_3297_),
    .Y(_0632_));
 sg13g2_a21oi_2 _4365_ (.B1(net1028),
    .Y(_0633_),
    .A2(_3278_),
    .A1(net1032));
 sg13g2_nor2_2 _4366_ (.A(net933),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_nand2_1 _4367_ (.Y(_0635_),
    .A(net187),
    .B(net844));
 sg13g2_o21ai_1 _4368_ (.B1(_0635_),
    .Y(_0128_),
    .A1(net844),
    .A2(_0634_));
 sg13g2_nand2_2 _4369_ (.Y(_0636_),
    .A(net1024),
    .B(net1028));
 sg13g2_nor2_1 _4370_ (.A(net1023),
    .B(net933),
    .Y(_0637_));
 sg13g2_xnor2_1 _4371_ (.Y(_0638_),
    .A(net945),
    .B(net933));
 sg13g2_xnor2_1 _4372_ (.Y(_0639_),
    .A(net1025),
    .B(net933));
 sg13g2_nand2_1 _4373_ (.Y(_0640_),
    .A(net205),
    .B(net844));
 sg13g2_o21ai_1 _4374_ (.B1(_0640_),
    .Y(_0129_),
    .A1(net844),
    .A2(_0638_));
 sg13g2_nand3_1 _4375_ (.B(net1022),
    .C(_0632_),
    .A(net1025),
    .Y(_0641_));
 sg13g2_a21o_1 _4376_ (.A2(net933),
    .A1(net1025),
    .B1(net1022),
    .X(_0642_));
 sg13g2_and2_2 _4377_ (.A(_0641_),
    .B(_0642_),
    .X(_0643_));
 sg13g2_nand2_1 _4378_ (.Y(_0644_),
    .A(net200),
    .B(net845));
 sg13g2_o21ai_1 _4379_ (.B1(_0644_),
    .Y(_0130_),
    .A1(net845),
    .A2(_0643_));
 sg13g2_or2_1 _4380_ (.X(_0645_),
    .B(_0641_),
    .A(_3112_));
 sg13g2_xnor2_1 _4381_ (.Y(_0646_),
    .A(_3112_),
    .B(_0641_));
 sg13g2_mux2_1 _4382_ (.A0(_0646_),
    .A1(net279),
    .S(net845),
    .X(_0131_));
 sg13g2_xor2_1 _4383_ (.B(_0645_),
    .A(net1018),
    .X(_0647_));
 sg13g2_mux2_1 _4384_ (.A0(_0647_),
    .A1(net278),
    .S(net845),
    .X(_0132_));
 sg13g2_nor4_2 _4385_ (.A(\vgademo.plane_dx_div.i[3] ),
    .B(\vgademo.plane_dx_div.i[2] ),
    .C(\vgademo.plane_dx_div.i[1] ),
    .Y(_0648_),
    .D(\vgademo.plane_dx_div.i[0] ));
 sg13g2_nor4_2 _4386_ (.A(_3123_),
    .B(net941),
    .C(_3125_),
    .Y(_0649_),
    .D(net984));
 sg13g2_and3_1 _4387_ (.X(_0650_),
    .A(_3212_),
    .B(_0578_),
    .C(_0649_));
 sg13g2_nand3_1 _4388_ (.B(_0578_),
    .C(_0649_),
    .A(_3212_),
    .Y(_0651_));
 sg13g2_nor2_1 _4389_ (.A(_0648_),
    .B(net929),
    .Y(_0652_));
 sg13g2_and2_1 _4390_ (.A(_0648_),
    .B(net926),
    .X(_0653_));
 sg13g2_nand2_2 _4391_ (.Y(_0654_),
    .A(_0648_),
    .B(_0651_));
 sg13g2_a22oi_1 _4392_ (.Y(_0133_),
    .B1(net906),
    .B2(_3098_),
    .A2(net907),
    .A1(_3099_));
 sg13g2_a22oi_1 _4393_ (.Y(_0655_),
    .B1(net906),
    .B2(\vgademo.plane_dx[2] ),
    .A2(net907),
    .A1(net544));
 sg13g2_inv_1 _4394_ (.Y(_0134_),
    .A(net545));
 sg13g2_a22oi_1 _4395_ (.Y(_0656_),
    .B1(net906),
    .B2(net570),
    .A2(net907),
    .A1(\vgademo.plane_dx[2] ));
 sg13g2_inv_1 _4396_ (.Y(_0135_),
    .A(net571));
 sg13g2_a22oi_1 _4397_ (.Y(_0657_),
    .B1(net906),
    .B2(net203),
    .A2(net907),
    .A1(\vgademo.plane_dx[3] ));
 sg13g2_inv_1 _4398_ (.Y(_0136_),
    .A(net204));
 sg13g2_a22oi_1 _4399_ (.Y(_0658_),
    .B1(net906),
    .B2(net1013),
    .A2(net907),
    .A1(net203));
 sg13g2_inv_1 _4400_ (.Y(_0137_),
    .A(_0658_));
 sg13g2_a22oi_1 _4401_ (.Y(_0659_),
    .B1(_0653_),
    .B2(net323),
    .A2(net907),
    .A1(net1013));
 sg13g2_inv_1 _4402_ (.Y(_0138_),
    .A(net324));
 sg13g2_a22oi_1 _4403_ (.Y(_0660_),
    .B1(net906),
    .B2(net247),
    .A2(net907),
    .A1(\vgademo.plane_dx_div.q[5] ));
 sg13g2_inv_1 _4404_ (.Y(_0139_),
    .A(net248));
 sg13g2_a22oi_1 _4405_ (.Y(_0661_),
    .B1(net905),
    .B2(net201),
    .A2(net907),
    .A1(net1011));
 sg13g2_inv_1 _4406_ (.Y(_0140_),
    .A(net202));
 sg13g2_a22oi_1 _4407_ (.Y(_0662_),
    .B1(net905),
    .B2(net1009),
    .A2(_0652_),
    .A1(net201));
 sg13g2_inv_1 _4408_ (.Y(_0141_),
    .A(_0662_));
 sg13g2_a22oi_1 _4409_ (.Y(_0663_),
    .B1(net906),
    .B2(net1007),
    .A2(net908),
    .A1(net1009));
 sg13g2_inv_1 _4410_ (.Y(_0142_),
    .A(_0663_));
 sg13g2_o21ai_1 _4411_ (.B1(_0651_),
    .Y(_0143_),
    .A1(_3095_),
    .A2(_0648_));
 sg13g2_xnor2_1 _4412_ (.Y(_0664_),
    .A(\vgademo.plane_dx_div.i[1] ),
    .B(net401));
 sg13g2_nor2_1 _4413_ (.A(net929),
    .B(net402),
    .Y(_0144_));
 sg13g2_a21o_1 _4414_ (.A2(net401),
    .A1(\vgademo.plane_dx_div.i[1] ),
    .B1(net538),
    .X(_0665_));
 sg13g2_nand3_1 _4415_ (.B(\vgademo.plane_dx_div.i[1] ),
    .C(net401),
    .A(net538),
    .Y(_0666_));
 sg13g2_and3_1 _4416_ (.X(_0145_),
    .A(net926),
    .B(net539),
    .C(_0666_));
 sg13g2_xor2_1 _4417_ (.B(_0666_),
    .A(net396),
    .X(_0667_));
 sg13g2_nor2_1 _4418_ (.A(net929),
    .B(net397),
    .Y(_0146_));
 sg13g2_nor2_1 _4419_ (.A(_0622_),
    .B(net934),
    .Y(_0668_));
 sg13g2_nand2_1 _4420_ (.Y(_0669_),
    .A(_0621_),
    .B(_0625_));
 sg13g2_nor2_1 _4421_ (.A(net326),
    .B(_0668_),
    .Y(_0670_));
 sg13g2_a21oi_1 _4422_ (.A1(net326),
    .A2(_0621_),
    .Y(_0147_),
    .B1(_0670_));
 sg13g2_and3_1 _4423_ (.X(_0671_),
    .A(\vgademo.audio_beat_out[1] ),
    .B(\vgademo.audio_beat_out[0] ),
    .C(_0621_));
 sg13g2_nand3_1 _4424_ (.B(net326),
    .C(_0621_),
    .A(net575),
    .Y(_0672_));
 sg13g2_a21o_1 _4425_ (.A2(_0621_),
    .A1(net326),
    .B1(net575),
    .X(_0673_));
 sg13g2_a21o_1 _4426_ (.A2(_0673_),
    .A1(_0672_),
    .B1(_0627_),
    .X(_0148_));
 sg13g2_o21ai_1 _4427_ (.B1(net846),
    .Y(_0674_),
    .A1(net508),
    .A2(_0672_));
 sg13g2_nor2_1 _4428_ (.A(net508),
    .B(_0622_),
    .Y(_0675_));
 sg13g2_a21oi_1 _4429_ (.A1(\vgademo.audio_beat_out[2] ),
    .A2(_0622_),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_a21oi_1 _4430_ (.A1(_0672_),
    .A2(net509),
    .Y(_0149_),
    .B1(_0674_));
 sg13g2_nor2_1 _4431_ (.A(net450),
    .B(_0674_),
    .Y(_0677_));
 sg13g2_nor3_1 _4432_ (.A(_3106_),
    .B(_0062_),
    .C(_0672_),
    .Y(_0678_));
 sg13g2_nor3_1 _4433_ (.A(_0627_),
    .B(net451),
    .C(_0678_),
    .Y(_0150_));
 sg13g2_nand3_1 _4434_ (.B(\vgademo.audio_beat_out[2] ),
    .C(_0671_),
    .A(net450),
    .Y(_0679_));
 sg13g2_xor2_1 _4435_ (.B(_0679_),
    .A(net491),
    .X(_0680_));
 sg13g2_nand2b_1 _4436_ (.Y(_0151_),
    .B(net492),
    .A_N(_0627_));
 sg13g2_a221oi_1 _4437_ (.B2(net1022),
    .C1(_0639_),
    .B1(_0634_),
    .A1(net944),
    .Y(_0681_),
    .A2(_3273_));
 sg13g2_nand2_1 _4438_ (.Y(_0682_),
    .A(net1019),
    .B(_0643_));
 sg13g2_nand2b_1 _4439_ (.Y(_0683_),
    .B(_0634_),
    .A_N(_3285_));
 sg13g2_o21ai_1 _4440_ (.B1(_0682_),
    .Y(_0684_),
    .A1(_0643_),
    .A2(_0683_));
 sg13g2_a21oi_1 _4441_ (.A1(_0638_),
    .A2(_0684_),
    .Y(_0685_),
    .B1(_0622_));
 sg13g2_o21ai_1 _4442_ (.B1(_0685_),
    .Y(_0686_),
    .A1(_3278_),
    .A2(_0681_));
 sg13g2_and2_1 _4443_ (.A(_0669_),
    .B(_0686_),
    .X(_0687_));
 sg13g2_nand2b_1 _4444_ (.Y(_0688_),
    .B(_3261_),
    .A_N(_0636_));
 sg13g2_and2_1 _4445_ (.A(net1035),
    .B(_3297_),
    .X(_0689_));
 sg13g2_a21oi_1 _4446_ (.A1(_3271_),
    .A2(_0689_),
    .Y(_0690_),
    .B1(net943));
 sg13g2_nor2b_1 _4447_ (.A(net1035),
    .B_N(net1032),
    .Y(_0691_));
 sg13g2_nand2_1 _4448_ (.Y(_0692_),
    .A(_3108_),
    .B(net1032));
 sg13g2_nor2_1 _4449_ (.A(_3109_),
    .B(net1028),
    .Y(_0693_));
 sg13g2_nand2_1 _4450_ (.Y(_0694_),
    .A(net1024),
    .B(net944));
 sg13g2_nor2_1 _4451_ (.A(_0692_),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_a21oi_1 _4452_ (.A1(_3109_),
    .A2(_3261_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_a22oi_1 _4453_ (.Y(_0697_),
    .B1(_0696_),
    .B2(net943),
    .A2(_0690_),
    .A1(_0688_));
 sg13g2_inv_1 _4454_ (.Y(_0698_),
    .A(_0697_));
 sg13g2_nor2_1 _4455_ (.A(_3295_),
    .B(_0698_),
    .Y(_0699_));
 sg13g2_nor3_2 _4456_ (.A(\vgademo.audio_kick_frames[1] ),
    .B(\vgademo.audio_kick_frames[0] ),
    .C(_3114_),
    .Y(_0700_));
 sg13g2_nand3b_1 _4457_ (.B(_3113_),
    .C(_0060_),
    .Y(_0701_),
    .A_N(\vgademo.audio_kick_frames[1] ));
 sg13g2_nand2_1 _4458_ (.Y(_0702_),
    .A(net1021),
    .B(_0693_));
 sg13g2_nor2_1 _4459_ (.A(_3260_),
    .B(_0702_),
    .Y(_0703_));
 sg13g2_nor2_1 _4460_ (.A(_0697_),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_nor2b_1 _4461_ (.A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[3] ),
    .Y(_0705_));
 sg13g2_xor2_1 _4462_ (.B(\vgademo.soundtrack.tri_osc_i[3] ),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(_0706_));
 sg13g2_o21ai_1 _4463_ (.B1(_0625_),
    .Y(_0707_),
    .A1(_0700_),
    .A2(_0706_));
 sg13g2_nor2b_1 _4464_ (.A(net1027),
    .B_N(net1031),
    .Y(_0708_));
 sg13g2_nand2_1 _4465_ (.Y(_0709_),
    .A(net1030),
    .B(_3266_));
 sg13g2_nand3_1 _4466_ (.B(_3299_),
    .C(_0709_),
    .A(_3287_),
    .Y(_0710_));
 sg13g2_nor2_1 _4467_ (.A(_3260_),
    .B(_0691_),
    .Y(_0711_));
 sg13g2_nand2_2 _4468_ (.Y(_0712_),
    .A(_3261_),
    .B(_0692_));
 sg13g2_a22oi_1 _4469_ (.Y(_0713_),
    .B1(_0712_),
    .B2(net1024),
    .A2(_3299_),
    .A1(_3271_));
 sg13g2_nand2_1 _4470_ (.Y(_0714_),
    .A(net1021),
    .B(_0713_));
 sg13g2_nand2_1 _4471_ (.Y(_0715_),
    .A(_0710_),
    .B(_0714_));
 sg13g2_o21ai_1 _4472_ (.B1(_3295_),
    .Y(_0716_),
    .A1(net1028),
    .A2(_0711_));
 sg13g2_nand3_1 _4473_ (.B(_0714_),
    .C(_0716_),
    .A(_0710_),
    .Y(_0717_));
 sg13g2_or2_1 _4474_ (.X(_0718_),
    .B(_0717_),
    .A(net932));
 sg13g2_o21ai_1 _4475_ (.B1(_0717_),
    .Y(_0719_),
    .A1(_0699_),
    .A2(_0704_));
 sg13g2_a21oi_1 _4476_ (.A1(_0700_),
    .A2(_0719_),
    .Y(_0720_),
    .B1(_0707_));
 sg13g2_mux2_1 _4477_ (.A0(_0720_),
    .A1(net487),
    .S(net838),
    .X(_0152_));
 sg13g2_nand2_1 _4478_ (.Y(_0721_),
    .A(net427),
    .B(net838));
 sg13g2_xnor2_1 _4479_ (.Y(_0722_),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .B(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_nand2b_1 _4480_ (.Y(_0723_),
    .B(_0722_),
    .A_N(_0705_));
 sg13g2_xnor2_1 _4481_ (.Y(_0724_),
    .A(_0705_),
    .B(_0722_));
 sg13g2_nor2_1 _4482_ (.A(_0699_),
    .B(_0717_),
    .Y(_0725_));
 sg13g2_nand2b_1 _4483_ (.Y(_0726_),
    .B(_0725_),
    .A_N(_0704_));
 sg13g2_a21oi_1 _4484_ (.A1(_0699_),
    .A2(_0715_),
    .Y(_0727_),
    .B1(net932));
 sg13g2_a22oi_1 _4485_ (.Y(_0728_),
    .B1(_0726_),
    .B2(_0727_),
    .A2(_0724_),
    .A1(net932));
 sg13g2_o21ai_1 _4486_ (.B1(_0721_),
    .Y(_0153_),
    .A1(_0669_),
    .A2(_0728_));
 sg13g2_nor2_1 _4487_ (.A(_3269_),
    .B(_3298_),
    .Y(_0729_));
 sg13g2_inv_1 _4488_ (.Y(_0730_),
    .A(_0729_));
 sg13g2_nand2_1 _4489_ (.Y(_0731_),
    .A(net1023),
    .B(_0730_));
 sg13g2_a221oi_1 _4490_ (.B2(net1024),
    .C1(net1021),
    .B1(_0730_),
    .A1(_3261_),
    .Y(_0732_),
    .A2(_0693_));
 sg13g2_nor2_1 _4491_ (.A(_0703_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_o21ai_1 _4492_ (.B1(_0690_),
    .Y(_0734_),
    .A1(_3261_),
    .A2(_0694_));
 sg13g2_nand2_1 _4493_ (.Y(_0735_),
    .A(net943),
    .B(_0695_));
 sg13g2_nand2_1 _4494_ (.Y(_0736_),
    .A(_0734_),
    .B(_0735_));
 sg13g2_nand2_1 _4495_ (.Y(_0737_),
    .A(_0733_),
    .B(_0736_));
 sg13g2_nor2_1 _4496_ (.A(_0697_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nor2b_1 _4497_ (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[2] ),
    .Y(_0739_));
 sg13g2_xor2_1 _4498_ (.B(\vgademo.soundtrack.tri_osc_i[5] ),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .X(_0740_));
 sg13g2_o21ai_1 _4499_ (.B1(_0723_),
    .Y(_0741_),
    .A1(_3146_),
    .A2(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_nor2b_1 _4500_ (.A(_0740_),
    .B_N(_0741_),
    .Y(_0742_));
 sg13g2_xor2_1 _4501_ (.B(_0741_),
    .A(_0740_),
    .X(_0743_));
 sg13g2_o21ai_1 _4502_ (.B1(_0700_),
    .Y(_0744_),
    .A1(_0725_),
    .A2(_0738_));
 sg13g2_o21ai_1 _4503_ (.B1(_0744_),
    .Y(_0745_),
    .A1(_0700_),
    .A2(_0743_));
 sg13g2_a22oi_1 _4504_ (.Y(_0746_),
    .B1(_0745_),
    .B2(net843),
    .A2(net838),
    .A1(net434));
 sg13g2_inv_1 _4505_ (.Y(_0154_),
    .A(_0746_));
 sg13g2_nor3_1 _4506_ (.A(_0703_),
    .B(_0732_),
    .C(_0736_),
    .Y(_0747_));
 sg13g2_nand2_1 _4507_ (.Y(_0748_),
    .A(_0697_),
    .B(_0747_));
 sg13g2_or2_1 _4508_ (.X(_0749_),
    .B(_0747_),
    .A(_0697_));
 sg13g2_o21ai_1 _4509_ (.B1(_0748_),
    .Y(_0750_),
    .A1(_0693_),
    .A2(_0749_));
 sg13g2_nand2_1 _4510_ (.Y(_0751_),
    .A(_0700_),
    .B(_0717_));
 sg13g2_nor3_1 _4511_ (.A(_0697_),
    .B(_0718_),
    .C(_0737_),
    .Y(_0752_));
 sg13g2_nand2_1 _4512_ (.Y(_0753_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(_3147_));
 sg13g2_xnor2_1 _4513_ (.Y(_0754_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_o21ai_1 _4514_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0739_),
    .A2(_0742_));
 sg13g2_or3_1 _4515_ (.A(_0739_),
    .B(_0742_),
    .C(_0754_),
    .X(_0756_));
 sg13g2_nand3_1 _4516_ (.B(_0755_),
    .C(_0756_),
    .A(net932),
    .Y(_0757_));
 sg13g2_o21ai_1 _4517_ (.B1(_0757_),
    .Y(_0758_),
    .A1(_0750_),
    .A2(_0751_));
 sg13g2_or2_1 _4518_ (.X(_0759_),
    .B(_0758_),
    .A(_0752_));
 sg13g2_a22oi_1 _4519_ (.Y(_0760_),
    .B1(_0759_),
    .B2(net843),
    .A2(net838),
    .A1(net558));
 sg13g2_inv_1 _4520_ (.Y(_0155_),
    .A(_0760_));
 sg13g2_xor2_1 _4521_ (.B(\vgademo.soundtrack.tri_osc_i[7] ),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(_0761_));
 sg13g2_a21oi_1 _4522_ (.A1(_0753_),
    .A2(_0755_),
    .Y(_0762_),
    .B1(_0761_));
 sg13g2_and3_1 _4523_ (.X(_0763_),
    .A(_0753_),
    .B(_0755_),
    .C(_0761_));
 sg13g2_nor3_1 _4524_ (.A(_0700_),
    .B(_0762_),
    .C(_0763_),
    .Y(_0764_));
 sg13g2_nand2b_1 _4525_ (.Y(_0765_),
    .B(_0737_),
    .A_N(_0699_));
 sg13g2_nor2_1 _4526_ (.A(_0751_),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_nor2_1 _4527_ (.A(_0764_),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_o21ai_1 _4528_ (.B1(_0767_),
    .Y(_0768_),
    .A1(_0718_),
    .A2(_0750_));
 sg13g2_a22oi_1 _4529_ (.Y(_0769_),
    .B1(_0768_),
    .B2(net843),
    .A2(net838),
    .A1(net569));
 sg13g2_inv_1 _4530_ (.Y(_0156_),
    .A(_0769_));
 sg13g2_nand2_1 _4531_ (.Y(_0770_),
    .A(net518),
    .B(net838));
 sg13g2_a21oi_1 _4532_ (.A1(\vgademo.soundtrack.tri_osc_i[4] ),
    .A2(_3148_),
    .Y(_0771_),
    .B1(_0762_));
 sg13g2_nor2_1 _4533_ (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(_3149_),
    .Y(_0772_));
 sg13g2_nand2_1 _4534_ (.Y(_0773_),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(_3149_));
 sg13g2_nand2b_1 _4535_ (.Y(_0774_),
    .B(_0773_),
    .A_N(_0772_));
 sg13g2_a21oi_1 _4536_ (.A1(_0771_),
    .A2(_0774_),
    .Y(_0775_),
    .B1(_0700_));
 sg13g2_o21ai_1 _4537_ (.B1(_0775_),
    .Y(_0776_),
    .A1(_0771_),
    .A2(_0774_));
 sg13g2_nor2_1 _4538_ (.A(_0749_),
    .B(_0751_),
    .Y(_0777_));
 sg13g2_o21ai_1 _4539_ (.B1(_0776_),
    .Y(_0778_),
    .A1(_0718_),
    .A2(_0765_));
 sg13g2_o21ai_1 _4540_ (.B1(net843),
    .Y(_0779_),
    .A1(_0777_),
    .A2(_0778_));
 sg13g2_nand2_1 _4541_ (.Y(_0157_),
    .A(_0770_),
    .B(_0779_));
 sg13g2_o21ai_1 _4542_ (.B1(_0773_),
    .Y(_0780_),
    .A1(_0771_),
    .A2(_0772_));
 sg13g2_xnor2_1 _4543_ (.Y(_0781_),
    .A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(_0780_));
 sg13g2_nand2b_1 _4544_ (.Y(_0782_),
    .B(_0747_),
    .A_N(_0717_));
 sg13g2_nor2_1 _4545_ (.A(_0697_),
    .B(net932),
    .Y(_0783_));
 sg13g2_a22oi_1 _4546_ (.Y(_0784_),
    .B1(_0782_),
    .B2(_0783_),
    .A2(_0781_),
    .A1(_0701_));
 sg13g2_a22oi_1 _4547_ (.Y(_0158_),
    .B1(_0784_),
    .B2(net843),
    .A2(_0687_),
    .A1(_3147_));
 sg13g2_nor3_1 _4548_ (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(\vgademo.soundtrack.tri_osc_i[7] ),
    .C(_0780_),
    .Y(_0785_));
 sg13g2_o21ai_1 _4549_ (.B1(\vgademo.soundtrack.tri_osc_i[7] ),
    .Y(_0786_),
    .A1(\vgademo.soundtrack.tri_osc_i[6] ),
    .A2(_0780_));
 sg13g2_nand2b_1 _4550_ (.Y(_0787_),
    .B(_0786_),
    .A_N(_0785_));
 sg13g2_o21ai_1 _4551_ (.B1(_0700_),
    .Y(_0788_),
    .A1(_0698_),
    .A2(_0717_));
 sg13g2_a21oi_1 _4552_ (.A1(_0698_),
    .A2(_0717_),
    .Y(_0789_),
    .B1(_0788_));
 sg13g2_a21oi_1 _4553_ (.A1(net932),
    .A2(_0787_),
    .Y(_0790_),
    .B1(_0789_));
 sg13g2_a22oi_1 _4554_ (.Y(_0159_),
    .B1(_0790_),
    .B2(net843),
    .A2(_0687_),
    .A1(_3148_));
 sg13g2_o21ai_1 _4555_ (.B1(net932),
    .Y(_0791_),
    .A1(_3149_),
    .A2(_0785_));
 sg13g2_nand2_1 _4556_ (.Y(_0792_),
    .A(_0788_),
    .B(_0791_));
 sg13g2_a22oi_1 _4557_ (.Y(_0160_),
    .B1(_0792_),
    .B2(net843),
    .A2(net838),
    .A1(_3149_));
 sg13g2_nor2_1 _4558_ (.A(net1050),
    .B(net240),
    .Y(_0793_));
 sg13g2_a21oi_2 _4559_ (.B1(_0564_),
    .Y(_0794_),
    .A2(_0565_),
    .A1(_0563_));
 sg13g2_a21oi_1 _4560_ (.A1(net1049),
    .A2(_0794_),
    .Y(_0161_),
    .B1(_0793_));
 sg13g2_mux2_1 _4561_ (.A0(\vgademo.soundtrack.tick_div[0] ),
    .A1(net174),
    .S(net871),
    .X(_0162_));
 sg13g2_a21o_1 _4562_ (.A2(net871),
    .A1(\vgademo.soundtrack.tick_div[0] ),
    .B1(net496),
    .X(_0795_));
 sg13g2_and2_1 _4563_ (.A(_0616_),
    .B(net497),
    .X(_0163_));
 sg13g2_xnor2_1 _4564_ (.Y(_0164_),
    .A(net242),
    .B(_0616_));
 sg13g2_xnor2_1 _4565_ (.Y(_0165_),
    .A(net250),
    .B(_0617_));
 sg13g2_xor2_1 _4566_ (.B(_0618_),
    .A(net213),
    .X(_0166_));
 sg13g2_xor2_1 _4567_ (.B(_0619_),
    .A(net276),
    .X(_0167_));
 sg13g2_a21oi_1 _4568_ (.A1(\vgademo.soundtrack.tick_div[5] ),
    .A2(_0619_),
    .Y(_0796_),
    .B1(net206));
 sg13g2_nor2_1 _4569_ (.A(_0620_),
    .B(net207),
    .Y(_0168_));
 sg13g2_xor2_1 _4570_ (.B(_0620_),
    .A(net290),
    .X(_0169_));
 sg13g2_nand2_1 _4571_ (.Y(_0797_),
    .A(net182),
    .B(net869));
 sg13g2_o21ai_1 _4572_ (.B1(_0797_),
    .Y(_0170_),
    .A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(net869));
 sg13g2_nand2_1 _4573_ (.Y(_0798_),
    .A(net184),
    .B(net869));
 sg13g2_o21ai_1 _4574_ (.B1(_0798_),
    .Y(_0171_),
    .A1(\vgademo.soundtrack.noise_lfsr[2] ),
    .A2(net869));
 sg13g2_nand2_1 _4575_ (.Y(_0799_),
    .A(net180),
    .B(net869));
 sg13g2_o21ai_1 _4576_ (.B1(_0799_),
    .Y(_0172_),
    .A1(\vgademo.soundtrack.noise_lfsr[3] ),
    .A2(net869));
 sg13g2_mux2_1 _4577_ (.A0(net236),
    .A1(_0040_),
    .S(net871),
    .X(_0173_));
 sg13g2_mux2_1 _4578_ (.A0(net232),
    .A1(\vgademo.soundtrack.noise_lfsr[5] ),
    .S(net872),
    .X(_0174_));
 sg13g2_mux2_1 _4579_ (.A0(_0098_),
    .A1(net170),
    .S(net872),
    .X(_0175_));
 sg13g2_mux2_1 _4580_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(net291),
    .S(net871),
    .X(_0176_));
 sg13g2_mux2_1 _4581_ (.A0(_0099_),
    .A1(net176),
    .S(net871),
    .X(_0177_));
 sg13g2_mux2_1 _4582_ (.A0(net329),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net871),
    .X(_0178_));
 sg13g2_mux2_1 _4583_ (.A0(net196),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net870),
    .X(_0179_));
 sg13g2_nand2_1 _4584_ (.Y(_0800_),
    .A(_0100_),
    .B(net870));
 sg13g2_o21ai_1 _4585_ (.B1(_0800_),
    .Y(_0180_),
    .A1(net166),
    .A2(net870));
 sg13g2_nand2_1 _4586_ (.Y(_0801_),
    .A(net194),
    .B(net870));
 sg13g2_o21ai_1 _4587_ (.B1(_0801_),
    .Y(_0181_),
    .A1(\vgademo.soundtrack.noise_lfsr[12] ),
    .A2(net869));
 sg13g2_mux2_1 _4588_ (.A0(_0102_),
    .A1(net172),
    .S(net871),
    .X(_0182_));
 sg13g2_xor2_1 _4589_ (.B(\vgademo.soundtrack.noise_lfsr[14] ),
    .A(\vgademo.soundtrack.noise_lfsr[0] ),
    .X(_0802_));
 sg13g2_mux2_1 _4590_ (.A0(net225),
    .A1(_0802_),
    .S(net871),
    .X(_0183_));
 sg13g2_mux2_1 _4591_ (.A0(net307),
    .A1(\vgademo.soundtrack.noise_lfsr[14] ),
    .S(net869),
    .X(_0184_));
 sg13g2_nor4_1 _4592_ (.A(_3264_),
    .B(_3274_),
    .C(net933),
    .D(_0633_),
    .Y(_0803_));
 sg13g2_nor2_1 _4593_ (.A(_3264_),
    .B(_0691_),
    .Y(_0804_));
 sg13g2_nand2_1 _4594_ (.Y(_0805_),
    .A(net1025),
    .B(_0634_));
 sg13g2_a21oi_1 _4595_ (.A1(_0804_),
    .A2(_0805_),
    .Y(_0806_),
    .B1(_0803_));
 sg13g2_a21oi_1 _4596_ (.A1(net1029),
    .A2(net1033),
    .Y(_0807_),
    .B1(net1038));
 sg13g2_nand3_1 _4597_ (.B(net1022),
    .C(_3279_),
    .A(net1025),
    .Y(_0808_));
 sg13g2_o21ai_1 _4598_ (.B1(_0682_),
    .Y(_0809_),
    .A1(_0807_),
    .A2(_0808_));
 sg13g2_o21ai_1 _4599_ (.B1(_0809_),
    .Y(_0810_),
    .A1(_0646_),
    .A2(_0806_));
 sg13g2_o21ai_1 _4600_ (.B1(net943),
    .Y(_0811_),
    .A1(_3264_),
    .A2(_3301_));
 sg13g2_nor2_1 _4601_ (.A(_0639_),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_o21ai_1 _4602_ (.B1(_0810_),
    .Y(_0813_),
    .A1(_0638_),
    .A2(_0804_));
 sg13g2_nor2_1 _4603_ (.A(_0812_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_o21ai_1 _4604_ (.B1(_0672_),
    .Y(_0815_),
    .A1(net846),
    .A2(_0814_));
 sg13g2_nand3_1 _4605_ (.B(net1005),
    .C(net998),
    .A(net1001),
    .Y(_0816_));
 sg13g2_or2_1 _4606_ (.X(_0817_),
    .B(_0816_),
    .A(_3152_));
 sg13g2_a21oi_1 _4607_ (.A1(net1005),
    .A2(_0817_),
    .Y(_0818_),
    .B1(_0624_));
 sg13g2_nor2_1 _4608_ (.A(net261),
    .B(_0815_),
    .Y(_0819_));
 sg13g2_a21oi_1 _4609_ (.A1(_0815_),
    .A2(_0818_),
    .Y(_0185_),
    .B1(_0819_));
 sg13g2_xnor2_1 _4610_ (.Y(_0820_),
    .A(net1001),
    .B(net1005));
 sg13g2_a21oi_1 _4611_ (.A1(_0817_),
    .A2(_0820_),
    .Y(_0821_),
    .B1(net934));
 sg13g2_nor2_1 _4612_ (.A(net249),
    .B(_0815_),
    .Y(_0822_));
 sg13g2_a21oi_1 _4613_ (.A1(_0815_),
    .A2(_0821_),
    .Y(_0186_),
    .B1(_0822_));
 sg13g2_nor2_1 _4614_ (.A(net994),
    .B(_0816_),
    .Y(_0823_));
 sg13g2_a21oi_1 _4615_ (.A1(net1001),
    .A2(net1005),
    .Y(_0824_),
    .B1(net998));
 sg13g2_nor3_1 _4616_ (.A(_0624_),
    .B(_0823_),
    .C(_0824_),
    .Y(_0825_));
 sg13g2_nor2_1 _4617_ (.A(net227),
    .B(_0815_),
    .Y(_0826_));
 sg13g2_a21oi_1 _4618_ (.A1(_0815_),
    .A2(_0825_),
    .Y(_0187_),
    .B1(_0826_));
 sg13g2_nor2_1 _4619_ (.A(net216),
    .B(_0815_),
    .Y(_0827_));
 sg13g2_a21oi_1 _4620_ (.A1(_3152_),
    .A2(_0816_),
    .Y(_0828_),
    .B1(_0624_));
 sg13g2_a21oi_1 _4621_ (.A1(_0815_),
    .A2(_0828_),
    .Y(_0188_),
    .B1(_0827_));
 sg13g2_and2_1 _4622_ (.A(net1045),
    .B(net873),
    .X(_0829_));
 sg13g2_nand2_1 _4623_ (.Y(_0830_),
    .A(net1048),
    .B(net873));
 sg13g2_nor2_1 _4624_ (.A(net1020),
    .B(net1019),
    .Y(_0831_));
 sg13g2_nand3b_1 _4625_ (.B(_3299_),
    .C(net1030),
    .Y(_0832_),
    .A_N(_3282_));
 sg13g2_o21ai_1 _4626_ (.B1(_0832_),
    .Y(_0833_),
    .A1(net1030),
    .A2(_3278_));
 sg13g2_inv_1 _4627_ (.Y(_0834_),
    .A(_0833_));
 sg13g2_nor2_1 _4628_ (.A(net1023),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_o21ai_1 _4629_ (.B1(_0630_),
    .Y(_0836_),
    .A1(_3266_),
    .A2(_3300_));
 sg13g2_a21oi_1 _4630_ (.A1(net1023),
    .A2(_0836_),
    .Y(_0837_),
    .B1(_0835_));
 sg13g2_nand2_1 _4631_ (.Y(_0838_),
    .A(net1038),
    .B(net944));
 sg13g2_nand3_1 _4632_ (.B(_0691_),
    .C(_0838_),
    .A(_3295_),
    .Y(_0839_));
 sg13g2_o21ai_1 _4633_ (.B1(_0839_),
    .Y(_0840_),
    .A1(net942),
    .A2(_0837_));
 sg13g2_nor2_1 _4634_ (.A(_3280_),
    .B(_0708_),
    .Y(_0841_));
 sg13g2_nor2b_1 _4635_ (.A(_0637_),
    .B_N(_0841_),
    .Y(_0842_));
 sg13g2_a21oi_1 _4636_ (.A1(net1020),
    .A2(_0842_),
    .Y(_0843_),
    .B1(net1016));
 sg13g2_o21ai_1 _4637_ (.B1(net943),
    .Y(_0844_),
    .A1(_3109_),
    .A2(_0730_));
 sg13g2_a22oi_1 _4638_ (.Y(_0845_),
    .B1(_0843_),
    .B2(_0844_),
    .A2(_0840_),
    .A1(net1016));
 sg13g2_a21oi_1 _4639_ (.A1(net1019),
    .A2(_0845_),
    .Y(_0846_),
    .B1(_0831_));
 sg13g2_nand3b_1 _4640_ (.B(_0711_),
    .C(net1037),
    .Y(_0847_),
    .A_N(_0708_));
 sg13g2_a21oi_1 _4641_ (.A1(_3263_),
    .A2(_3269_),
    .Y(_0848_),
    .B1(net1023));
 sg13g2_a21oi_1 _4642_ (.A1(net1030),
    .A2(_3278_),
    .Y(_0849_),
    .B1(_0636_));
 sg13g2_a21oi_1 _4643_ (.A1(_0847_),
    .A2(_0848_),
    .Y(_0850_),
    .B1(_0849_));
 sg13g2_nand2b_1 _4644_ (.Y(_0851_),
    .B(net1020),
    .A_N(_0850_));
 sg13g2_nand2b_1 _4645_ (.Y(_0852_),
    .B(net944),
    .A_N(_0629_));
 sg13g2_nor3_1 _4646_ (.A(_3266_),
    .B(_3278_),
    .C(_3301_),
    .Y(_0853_));
 sg13g2_nand2_1 _4647_ (.Y(_0854_),
    .A(_0852_),
    .B(_0853_));
 sg13g2_nand2_1 _4648_ (.Y(_0855_),
    .A(_3295_),
    .B(_0854_));
 sg13g2_a21o_1 _4649_ (.A2(_3299_),
    .A1(_3267_),
    .B1(net1031),
    .X(_0856_));
 sg13g2_nand3_1 _4650_ (.B(_0852_),
    .C(_0856_),
    .A(_3287_),
    .Y(_0857_));
 sg13g2_nand3_1 _4651_ (.B(_0855_),
    .C(_0857_),
    .A(_0851_),
    .Y(_0858_));
 sg13g2_nand2_1 _4652_ (.Y(_0859_),
    .A(_3107_),
    .B(net1019));
 sg13g2_nand2_1 _4653_ (.Y(_0860_),
    .A(net1020),
    .B(_0636_));
 sg13g2_nor2_1 _4654_ (.A(_0637_),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_nor2_1 _4655_ (.A(net1017),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_nand3_1 _4656_ (.B(net1027),
    .C(_0712_),
    .A(net945),
    .Y(_0863_));
 sg13g2_nand3_1 _4657_ (.B(_0731_),
    .C(_0863_),
    .A(net942),
    .Y(_0864_));
 sg13g2_a221oi_1 _4658_ (.B2(_0864_),
    .C1(_0859_),
    .B1(_0862_),
    .A1(net1017),
    .Y(_0865_),
    .A2(_0858_));
 sg13g2_nor2_1 _4659_ (.A(\vgademo.audio_beat_out[2] ),
    .B(net1019),
    .Y(_0866_));
 sg13g2_nor2b_1 _4660_ (.A(_0702_),
    .B_N(_0866_),
    .Y(_0867_));
 sg13g2_nor2_1 _4661_ (.A(_0865_),
    .B(_0867_),
    .Y(_0868_));
 sg13g2_o21ai_1 _4662_ (.B1(_0868_),
    .Y(_0869_),
    .A1(_3107_),
    .A2(_0846_));
 sg13g2_inv_1 _4663_ (.Y(_0870_),
    .A(net857));
 sg13g2_nand3_1 _4664_ (.B(_3295_),
    .C(_0712_),
    .A(net1028),
    .Y(_0871_));
 sg13g2_o21ai_1 _4665_ (.B1(_3287_),
    .Y(_0872_),
    .A1(_3298_),
    .A2(_0633_));
 sg13g2_o21ai_1 _4666_ (.B1(net1021),
    .Y(_0873_),
    .A1(_3274_),
    .A2(_0694_));
 sg13g2_and2_1 _4667_ (.A(_0872_),
    .B(_0873_),
    .X(_0874_));
 sg13g2_o21ai_1 _4668_ (.B1(_0874_),
    .Y(_0875_),
    .A1(_3296_),
    .A2(_0854_));
 sg13g2_a22oi_1 _4669_ (.Y(_0876_),
    .B1(_0875_),
    .B2(net1017),
    .A2(_0871_),
    .A1(_0862_));
 sg13g2_nand3_1 _4670_ (.B(_3270_),
    .C(_3299_),
    .A(net1023),
    .Y(_0877_));
 sg13g2_nand3_1 _4671_ (.B(_0834_),
    .C(_0877_),
    .A(net1020),
    .Y(_0878_));
 sg13g2_nand2_1 _4672_ (.Y(_0879_),
    .A(_3261_),
    .B(_3287_));
 sg13g2_nor4_1 _4673_ (.A(_3269_),
    .B(_3282_),
    .C(net933),
    .D(_0879_),
    .Y(_0880_));
 sg13g2_a21oi_1 _4674_ (.A1(_3295_),
    .A2(net933),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_nand3_1 _4675_ (.B(_0878_),
    .C(_0881_),
    .A(net1017),
    .Y(_0882_));
 sg13g2_nand2_1 _4676_ (.Y(_0883_),
    .A(\vgademo.audio_beat_out[2] ),
    .B(net1019));
 sg13g2_o21ai_1 _4677_ (.B1(_3287_),
    .Y(_0884_),
    .A1(_3276_),
    .A2(_0708_));
 sg13g2_a21oi_1 _4678_ (.A1(_0843_),
    .A2(_0884_),
    .Y(_0885_),
    .B1(_0883_));
 sg13g2_nor2b_1 _4679_ (.A(_3295_),
    .B_N(_0866_),
    .Y(_0886_));
 sg13g2_a22oi_1 _4680_ (.Y(_0887_),
    .B1(_0886_),
    .B2(_0702_),
    .A2(_0885_),
    .A1(_0882_));
 sg13g2_o21ai_1 _4681_ (.B1(_0887_),
    .Y(_0888_),
    .A1(_0859_),
    .A2(_0876_));
 sg13g2_o21ai_1 _4682_ (.B1(net1016),
    .Y(_0889_),
    .A1(_0835_),
    .A2(_0873_));
 sg13g2_o21ai_1 _4683_ (.B1(_3112_),
    .Y(_0890_),
    .A1(net942),
    .A2(_0636_));
 sg13g2_a21o_1 _4684_ (.A2(_0860_),
    .A1(_0844_),
    .B1(net1016),
    .X(_0891_));
 sg13g2_nand3_1 _4685_ (.B(_0890_),
    .C(_0891_),
    .A(_0889_),
    .Y(_0892_));
 sg13g2_a221oi_1 _4686_ (.B2(_0848_),
    .C1(net942),
    .B1(_0847_),
    .A1(net944),
    .Y(_0893_),
    .A2(_3274_));
 sg13g2_nor2b_1 _4687_ (.A(_0893_),
    .B_N(net1016),
    .Y(_0894_));
 sg13g2_a21oi_1 _4688_ (.A1(net1020),
    .A2(_0638_),
    .Y(_0895_),
    .B1(net1016));
 sg13g2_a22oi_1 _4689_ (.Y(_0896_),
    .B1(_0895_),
    .B2(_0731_),
    .A2(_0894_),
    .A1(_0857_));
 sg13g2_a22oi_1 _4690_ (.Y(_0897_),
    .B1(_0892_),
    .B2(\vgademo.audio_beat_out[2] ),
    .A2(_0866_),
    .A1(net945));
 sg13g2_o21ai_1 _4691_ (.B1(_0897_),
    .Y(_0898_),
    .A1(_0859_),
    .A2(_0896_));
 sg13g2_nor2b_1 _4692_ (.A(_0888_),
    .B_N(_0898_),
    .Y(_0899_));
 sg13g2_or2_1 _4693_ (.X(_0900_),
    .B(_0899_),
    .A(net857));
 sg13g2_inv_1 _4694_ (.Y(_0901_),
    .A(_0900_));
 sg13g2_nor2_1 _4695_ (.A(_0888_),
    .B(_0898_),
    .Y(_0902_));
 sg13g2_inv_1 _4696_ (.Y(_0903_),
    .A(_0902_));
 sg13g2_a21oi_2 _4697_ (.B1(_0901_),
    .Y(_0904_),
    .A2(_0903_),
    .A1(net857));
 sg13g2_nor2_1 _4698_ (.A(net860),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_xnor2_1 _4699_ (.Y(_0189_),
    .A(_3205_),
    .B(_0905_));
 sg13g2_nor2_1 _4700_ (.A(_0042_),
    .B(_0901_),
    .Y(_0906_));
 sg13g2_xor2_1 _4701_ (.B(_0900_),
    .A(_0042_),
    .X(_0907_));
 sg13g2_nor3_2 _4702_ (.A(_3205_),
    .B(_0904_),
    .C(_0907_),
    .Y(_0908_));
 sg13g2_o21ai_1 _4703_ (.B1(_0907_),
    .Y(_0909_),
    .A1(_3205_),
    .A2(_0904_));
 sg13g2_nand2_1 _4704_ (.Y(_0910_),
    .A(net864),
    .B(_0909_));
 sg13g2_nand2_1 _4705_ (.Y(_0911_),
    .A(net190),
    .B(net860));
 sg13g2_o21ai_1 _4706_ (.B1(_0911_),
    .Y(_0190_),
    .A1(_0908_),
    .A2(_0910_));
 sg13g2_or2_1 _4707_ (.X(_0912_),
    .B(_0902_),
    .A(net857));
 sg13g2_nand2b_1 _4708_ (.Y(_0913_),
    .B(_0888_),
    .A_N(_0898_));
 sg13g2_nand2_2 _4709_ (.Y(_0914_),
    .A(net857),
    .B(_0913_));
 sg13g2_nand2_1 _4710_ (.Y(_0915_),
    .A(_0912_),
    .B(_0914_));
 sg13g2_nand3_1 _4711_ (.B(_0912_),
    .C(_0914_),
    .A(net309),
    .Y(_0916_));
 sg13g2_xnor2_1 _4712_ (.Y(_0917_),
    .A(\vgademo.soundtrack.pulse_osc_p[2] ),
    .B(_0915_));
 sg13g2_o21ai_1 _4713_ (.B1(_0917_),
    .Y(_0918_),
    .A1(_0906_),
    .A2(_0908_));
 sg13g2_or3_1 _4714_ (.A(_0906_),
    .B(_0908_),
    .C(_0917_),
    .X(_0919_));
 sg13g2_a21oi_1 _4715_ (.A1(_0918_),
    .A2(_0919_),
    .Y(_0920_),
    .B1(net859));
 sg13g2_a21oi_1 _4716_ (.A1(_3206_),
    .A2(net859),
    .Y(_0191_),
    .B1(_0920_));
 sg13g2_nand2_1 _4717_ (.Y(_0921_),
    .A(_0888_),
    .B(_0898_));
 sg13g2_nor2_1 _4718_ (.A(_0899_),
    .B(_0914_),
    .Y(_0922_));
 sg13g2_a21oi_1 _4719_ (.A1(_0870_),
    .A2(_0921_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_nand2b_1 _4720_ (.Y(_0924_),
    .B(\vgademo.soundtrack.pulse_osc_p[3] ),
    .A_N(_0923_));
 sg13g2_xnor2_1 _4721_ (.Y(_0925_),
    .A(_3207_),
    .B(_0923_));
 sg13g2_a21o_1 _4722_ (.A2(_0918_),
    .A1(_0916_),
    .B1(_0925_),
    .X(_0926_));
 sg13g2_nand3_1 _4723_ (.B(_0918_),
    .C(_0925_),
    .A(_0916_),
    .Y(_0927_));
 sg13g2_a21oi_1 _4724_ (.A1(_0926_),
    .A2(_0927_),
    .Y(_0928_),
    .B1(net859));
 sg13g2_a21oi_1 _4725_ (.A1(_3207_),
    .A2(net859),
    .Y(_0192_),
    .B1(_0928_));
 sg13g2_nand2b_1 _4726_ (.Y(_0929_),
    .B(_0914_),
    .A_N(_0899_));
 sg13g2_and2_1 _4727_ (.A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .B(_0929_),
    .X(_0930_));
 sg13g2_xnor2_1 _4728_ (.Y(_0931_),
    .A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .B(_0929_));
 sg13g2_a21oi_1 _4729_ (.A1(_0924_),
    .A2(_0926_),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_and3_1 _4730_ (.X(_0933_),
    .A(_0924_),
    .B(_0926_),
    .C(_0931_));
 sg13g2_nor3_1 _4731_ (.A(net859),
    .B(_0932_),
    .C(_0933_),
    .Y(_0934_));
 sg13g2_a21o_1 _4732_ (.A2(net859),
    .A1(net342),
    .B1(_0934_),
    .X(_0193_));
 sg13g2_nand2_1 _4733_ (.Y(_0935_),
    .A(_0912_),
    .B(_0921_));
 sg13g2_nand3_1 _4734_ (.B(_0912_),
    .C(_0921_),
    .A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .Y(_0936_));
 sg13g2_xnor2_1 _4735_ (.Y(_0937_),
    .A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .B(_0935_));
 sg13g2_o21ai_1 _4736_ (.B1(_0937_),
    .Y(_0938_),
    .A1(_0930_),
    .A2(_0932_));
 sg13g2_or3_1 _4737_ (.A(_0930_),
    .B(_0932_),
    .C(_0937_),
    .X(_0939_));
 sg13g2_a21oi_1 _4738_ (.A1(_0938_),
    .A2(_0939_),
    .Y(_0940_),
    .B1(net859));
 sg13g2_a21oi_1 _4739_ (.A1(_3208_),
    .A2(net859),
    .Y(_0194_),
    .B1(_0940_));
 sg13g2_nand2_1 _4740_ (.Y(_0941_),
    .A(net288),
    .B(net860));
 sg13g2_xnor2_1 _4741_ (.Y(_0942_),
    .A(net288),
    .B(net857));
 sg13g2_a21oi_1 _4742_ (.A1(_0936_),
    .A2(_0938_),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_nand3_1 _4743_ (.B(_0938_),
    .C(_0942_),
    .A(_0936_),
    .Y(_0944_));
 sg13g2_nand2_1 _4744_ (.Y(_0945_),
    .A(net864),
    .B(_0944_));
 sg13g2_o21ai_1 _4745_ (.B1(_0941_),
    .Y(_0195_),
    .A1(_0943_),
    .A2(_0945_));
 sg13g2_nor2_1 _4746_ (.A(net362),
    .B(net864),
    .Y(_0946_));
 sg13g2_nand2b_1 _4747_ (.Y(_0947_),
    .B(net857),
    .A_N(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_a21o_1 _4748_ (.A2(_0869_),
    .A1(\vgademo.soundtrack.pulse_osc_p[6] ),
    .B1(_0943_),
    .X(_0948_));
 sg13g2_a21o_1 _4749_ (.A2(_0870_),
    .A1(\vgademo.soundtrack.pulse_osc_p[7] ),
    .B1(_0948_),
    .X(_0949_));
 sg13g2_xnor2_1 _4750_ (.Y(_0950_),
    .A(net362),
    .B(net857));
 sg13g2_xnor2_1 _4751_ (.Y(_0951_),
    .A(_0948_),
    .B(_0950_));
 sg13g2_a21oi_1 _4752_ (.A1(net864),
    .A2(_0951_),
    .Y(_0196_),
    .B1(_0946_));
 sg13g2_and3_1 _4753_ (.X(_0952_),
    .A(net864),
    .B(_0947_),
    .C(_0949_));
 sg13g2_xor2_1 _4754_ (.B(_0952_),
    .A(net271),
    .X(_0197_));
 sg13g2_a21oi_1 _4755_ (.A1(\vgademo.soundtrack.pulse_osc_p[8] ),
    .A2(_0952_),
    .Y(_0953_),
    .B1(net256));
 sg13g2_and3_1 _4756_ (.X(_0954_),
    .A(\vgademo.soundtrack.pulse_osc_p[8] ),
    .B(net256),
    .C(_0952_));
 sg13g2_nor2_1 _4757_ (.A(net257),
    .B(_0954_),
    .Y(_0198_));
 sg13g2_and2_1 _4758_ (.A(net222),
    .B(_0954_),
    .X(_0955_));
 sg13g2_xor2_1 _4759_ (.B(_0954_),
    .A(net222),
    .X(_0199_));
 sg13g2_xor2_1 _4760_ (.B(_0955_),
    .A(net275),
    .X(_0200_));
 sg13g2_nand3_1 _4761_ (.B(net275),
    .C(_0955_),
    .A(net495),
    .Y(_0956_));
 sg13g2_a21o_1 _4762_ (.A2(_0955_),
    .A1(net275),
    .B1(net495),
    .X(_0957_));
 sg13g2_and2_1 _4763_ (.A(_0956_),
    .B(_0957_),
    .X(_0201_));
 sg13g2_xnor2_1 _4764_ (.Y(_0202_),
    .A(net263),
    .B(_0956_));
 sg13g2_nor2_1 _4765_ (.A(\vgademo.audio_kick_frames[0] ),
    .B(net838),
    .Y(_0958_));
 sg13g2_o21ai_1 _4766_ (.B1(_0958_),
    .Y(_0959_),
    .A1(net934),
    .A2(net932));
 sg13g2_o21ai_1 _4767_ (.B1(_0959_),
    .Y(_0203_),
    .A1(_3113_),
    .A2(net843));
 sg13g2_or2_1 _4768_ (.X(_0960_),
    .B(_0959_),
    .A(net430));
 sg13g2_nand2_1 _4769_ (.Y(_0961_),
    .A(net430),
    .B(_0959_));
 sg13g2_or2_1 _4770_ (.X(_0962_),
    .B(_0686_),
    .A(_0625_));
 sg13g2_nand3_1 _4771_ (.B(_0961_),
    .C(_0962_),
    .A(_0960_),
    .Y(_0204_));
 sg13g2_o21ai_1 _4772_ (.B1(_0962_),
    .Y(_0963_),
    .A1(net280),
    .A2(_0960_));
 sg13g2_a21o_1 _4773_ (.A2(_0960_),
    .A1(net280),
    .B1(_0963_),
    .X(_0205_));
 sg13g2_nand2_1 _4774_ (.Y(_0964_),
    .A(net1025),
    .B(_0629_));
 sg13g2_nor2_1 _4775_ (.A(_0804_),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_nand3_1 _4776_ (.B(net1033),
    .C(_3280_),
    .A(net1029),
    .Y(_0966_));
 sg13g2_a21oi_1 _4777_ (.A1(_0852_),
    .A2(_0966_),
    .Y(_0967_),
    .B1(_0638_));
 sg13g2_or3_1 _4778_ (.A(_0647_),
    .B(_0965_),
    .C(_0967_),
    .X(_0968_));
 sg13g2_nor2b_1 _4779_ (.A(_0634_),
    .B_N(_3286_),
    .Y(_0969_));
 sg13g2_o21ai_1 _4780_ (.B1(_0639_),
    .Y(_0970_),
    .A1(_0803_),
    .A2(_0969_));
 sg13g2_nand3_1 _4781_ (.B(_0638_),
    .C(_0709_),
    .A(_3281_),
    .Y(_0971_));
 sg13g2_nand3_1 _4782_ (.B(_0970_),
    .C(_0971_),
    .A(_0647_),
    .Y(_0972_));
 sg13g2_xnor2_1 _4783_ (.Y(_0973_),
    .A(net1028),
    .B(_3261_));
 sg13g2_nand2_1 _4784_ (.Y(_0974_),
    .A(net1038),
    .B(_0973_));
 sg13g2_nand2_1 _4785_ (.Y(_0975_),
    .A(_0639_),
    .B(_0974_));
 sg13g2_nand2_1 _4786_ (.Y(_0976_),
    .A(net1026),
    .B(_3279_));
 sg13g2_nand3_1 _4787_ (.B(_0975_),
    .C(_0976_),
    .A(_0643_),
    .Y(_0977_));
 sg13g2_a22oi_1 _4788_ (.Y(_0978_),
    .B1(_0977_),
    .B2(_0682_),
    .A2(_0972_),
    .A1(_0968_));
 sg13g2_nand2b_1 _4789_ (.Y(_0979_),
    .B(_0712_),
    .A_N(net1038));
 sg13g2_nand4_1 _4790_ (.B(_0973_),
    .C(_0975_),
    .A(_0647_),
    .Y(_0980_),
    .D(_0979_));
 sg13g2_nand3_1 _4791_ (.B(_3266_),
    .C(_3302_),
    .A(net945),
    .Y(_0981_));
 sg13g2_o21ai_1 _4792_ (.B1(_0981_),
    .Y(_0982_),
    .A1(_0805_),
    .A2(_0841_));
 sg13g2_o21ai_1 _4793_ (.B1(_0980_),
    .Y(_0983_),
    .A1(_0647_),
    .A2(_0982_));
 sg13g2_a21oi_1 _4794_ (.A1(_0646_),
    .A2(_0974_),
    .Y(_0984_),
    .B1(_0643_));
 sg13g2_a21o_1 _4795_ (.A2(_0984_),
    .A1(_0983_),
    .B1(_0625_),
    .X(_0985_));
 sg13g2_o21ai_1 _4796_ (.B1(_0674_),
    .Y(_0986_),
    .A1(_0978_),
    .A2(_0985_));
 sg13g2_a21oi_1 _4797_ (.A1(net992),
    .A2(_3341_),
    .Y(_0987_),
    .B1(net934));
 sg13g2_nand2_1 _4798_ (.Y(_0988_),
    .A(net178),
    .B(_0986_));
 sg13g2_o21ai_1 _4799_ (.B1(_0988_),
    .Y(_0206_),
    .A1(_0986_),
    .A2(_0987_));
 sg13g2_a21oi_1 _4800_ (.A1(_3341_),
    .A2(_3350_),
    .Y(_0989_),
    .B1(net934));
 sg13g2_nand2_1 _4801_ (.Y(_0990_),
    .A(net186),
    .B(_0986_));
 sg13g2_o21ai_1 _4802_ (.B1(_0990_),
    .Y(_0207_),
    .A1(_0986_),
    .A2(_0989_));
 sg13g2_nand2_1 _4803_ (.Y(_0991_),
    .A(net192),
    .B(_0986_));
 sg13g2_a221oi_1 _4804_ (.B2(net992),
    .C1(net934),
    .B1(_0441_),
    .A1(_3150_),
    .Y(_0992_),
    .A2(_3348_));
 sg13g2_o21ai_1 _4805_ (.B1(_0991_),
    .Y(_0208_),
    .A1(_0986_),
    .A2(_0992_));
 sg13g2_a21oi_1 _4806_ (.A1(\vgademo.soundtrack.pulse_vol[0] ),
    .A2(_3340_),
    .Y(_0993_),
    .B1(net990));
 sg13g2_nor2_1 _4807_ (.A(net934),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_nand2_1 _4808_ (.Y(_0995_),
    .A(net198),
    .B(_0986_));
 sg13g2_o21ai_1 _4809_ (.B1(_0995_),
    .Y(_0209_),
    .A1(_0986_),
    .A2(_0994_));
 sg13g2_nand2_1 _4810_ (.Y(_0996_),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B(net864));
 sg13g2_xnor2_1 _4811_ (.Y(_0210_),
    .A(net259),
    .B(_0996_));
 sg13g2_nand2_1 _4812_ (.Y(_0997_),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B(net259));
 sg13g2_xor2_1 _4813_ (.B(\vgademo.soundtrack.tri_osc_p[1] ),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(_0998_));
 sg13g2_nor2b_1 _4814_ (.A(_0997_),
    .B_N(_0998_),
    .Y(_0999_));
 sg13g2_xor2_1 _4815_ (.B(_0998_),
    .A(_0997_),
    .X(_1000_));
 sg13g2_nand2_1 _4816_ (.Y(_1001_),
    .A(net394),
    .B(net860));
 sg13g2_o21ai_1 _4817_ (.B1(_1001_),
    .Y(_0211_),
    .A1(net860),
    .A2(_1000_));
 sg13g2_nor2_1 _4818_ (.A(net416),
    .B(net862),
    .Y(_1002_));
 sg13g2_nand2_1 _4819_ (.Y(_1003_),
    .A(net592),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_xnor2_1 _4820_ (.Y(_1004_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_a21oi_1 _4821_ (.A1(\vgademo.soundtrack.tri_osc_i[1] ),
    .A2(\vgademo.soundtrack.tri_osc_p[1] ),
    .Y(_1005_),
    .B1(_0999_));
 sg13g2_or2_1 _4822_ (.X(_1006_),
    .B(_1005_),
    .A(_1004_));
 sg13g2_xnor2_1 _4823_ (.Y(_1007_),
    .A(_1004_),
    .B(_1005_));
 sg13g2_a21oi_1 _4824_ (.A1(net864),
    .A2(_1007_),
    .Y(_0212_),
    .B1(_1002_));
 sg13g2_nor2_1 _4825_ (.A(net409),
    .B(net862),
    .Y(_1008_));
 sg13g2_xnor2_1 _4826_ (.Y(_1009_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_a21oi_1 _4827_ (.A1(_1003_),
    .A2(_1006_),
    .Y(_1010_),
    .B1(_1009_));
 sg13g2_nand3_1 _4828_ (.B(_1006_),
    .C(_1009_),
    .A(net593),
    .Y(_1011_));
 sg13g2_nand2b_1 _4829_ (.Y(_1012_),
    .B(_1011_),
    .A_N(_1010_));
 sg13g2_a21oi_1 _4830_ (.A1(net862),
    .A2(_1012_),
    .Y(_0213_),
    .B1(_1008_));
 sg13g2_nor2_1 _4831_ (.A(net374),
    .B(net862),
    .Y(_1013_));
 sg13g2_nand2_1 _4832_ (.Y(_1014_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_xnor2_1 _4833_ (.Y(_1015_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_a21oi_1 _4834_ (.A1(\vgademo.soundtrack.tri_osc_i[3] ),
    .A2(\vgademo.soundtrack.tri_osc_p[3] ),
    .Y(_1016_),
    .B1(_1010_));
 sg13g2_xnor2_1 _4835_ (.Y(_1017_),
    .A(_1015_),
    .B(_1016_));
 sg13g2_a21oi_1 _4836_ (.A1(net862),
    .A2(_1017_),
    .Y(_0214_),
    .B1(_1013_));
 sg13g2_nor2_1 _4837_ (.A(net447),
    .B(net863),
    .Y(_1018_));
 sg13g2_o21ai_1 _4838_ (.B1(_1014_),
    .Y(_1019_),
    .A1(_1015_),
    .A2(_1016_));
 sg13g2_nand2_1 _4839_ (.Y(_1020_),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_xor2_1 _4840_ (.B(\vgademo.soundtrack.tri_osc_p[5] ),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(_1021_));
 sg13g2_xnor2_1 _4841_ (.Y(_1022_),
    .A(_1019_),
    .B(_1021_));
 sg13g2_a21oi_1 _4842_ (.A1(net862),
    .A2(_1022_),
    .Y(_0215_),
    .B1(_1018_));
 sg13g2_nor2_1 _4843_ (.A(_3147_),
    .B(_3204_),
    .Y(_1023_));
 sg13g2_xnor2_1 _4844_ (.Y(_1024_),
    .A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_o21ai_1 _4845_ (.B1(_1019_),
    .Y(_1025_),
    .A1(\vgademo.soundtrack.tri_osc_i[5] ),
    .A2(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_nand3_1 _4846_ (.B(_1024_),
    .C(_1025_),
    .A(_1020_),
    .Y(_1026_));
 sg13g2_a21oi_1 _4847_ (.A1(_1020_),
    .A2(_1025_),
    .Y(_1027_),
    .B1(_1024_));
 sg13g2_nand3b_1 _4848_ (.B(net863),
    .C(_1026_),
    .Y(_1028_),
    .A_N(_1027_));
 sg13g2_o21ai_1 _4849_ (.B1(_1028_),
    .Y(_0216_),
    .A1(_3204_),
    .A2(net862));
 sg13g2_nand2_1 _4850_ (.Y(_1029_),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .B(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_xor2_1 _4851_ (.B(\vgademo.soundtrack.tri_osc_p[7] ),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(_1030_));
 sg13g2_or3_1 _4852_ (.A(_1023_),
    .B(_1027_),
    .C(_1030_),
    .X(_1031_));
 sg13g2_o21ai_1 _4853_ (.B1(_1030_),
    .Y(_1032_),
    .A1(_1023_),
    .A2(_1027_));
 sg13g2_nand3_1 _4854_ (.B(_1031_),
    .C(_1032_),
    .A(net862),
    .Y(_1033_));
 sg13g2_o21ai_1 _4855_ (.B1(_1033_),
    .Y(_0217_),
    .A1(_3203_),
    .A2(net863));
 sg13g2_xnor2_1 _4856_ (.Y(_1034_),
    .A(\vgademo.soundtrack.tri_osc_i[8] ),
    .B(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_and3_1 _4857_ (.X(_1035_),
    .A(_1029_),
    .B(_1032_),
    .C(_1034_));
 sg13g2_a21oi_1 _4858_ (.A1(_1029_),
    .A2(_1032_),
    .Y(_1036_),
    .B1(_1034_));
 sg13g2_nor3_1 _4859_ (.A(net861),
    .B(_1035_),
    .C(_1036_),
    .Y(_1037_));
 sg13g2_a21o_1 _4860_ (.A2(net861),
    .A1(net420),
    .B1(_1037_),
    .X(_0218_));
 sg13g2_a21oi_1 _4861_ (.A1(\vgademo.soundtrack.tri_osc_i[8] ),
    .A2(\vgademo.soundtrack.tri_osc_p[8] ),
    .Y(_1038_),
    .B1(_1036_));
 sg13g2_nand3_1 _4862_ (.B(net863),
    .C(_1038_),
    .A(net386),
    .Y(_1039_));
 sg13g2_nor3_2 _4863_ (.A(net386),
    .B(net861),
    .C(_1038_),
    .Y(_1040_));
 sg13g2_o21ai_1 _4864_ (.B1(_1039_),
    .Y(_1041_),
    .A1(\vgademo.soundtrack.tri_osc_p[9] ),
    .A2(net863));
 sg13g2_nor2_1 _4865_ (.A(_1040_),
    .B(_1041_),
    .Y(_0219_));
 sg13g2_and2_1 _4866_ (.A(net281),
    .B(_1040_),
    .X(_1042_));
 sg13g2_xor2_1 _4867_ (.B(_1040_),
    .A(net281),
    .X(_0220_));
 sg13g2_xor2_1 _4868_ (.B(_1042_),
    .A(net440),
    .X(_0221_));
 sg13g2_nand3_1 _4869_ (.B(net440),
    .C(_1042_),
    .A(net407),
    .Y(_1043_));
 sg13g2_a21o_1 _4870_ (.A2(_1042_),
    .A1(net440),
    .B1(net407),
    .X(_1044_));
 sg13g2_and2_1 _4871_ (.A(_1043_),
    .B(_1044_),
    .X(_0222_));
 sg13g2_nand4_1 _4872_ (.B(net407),
    .C(net587),
    .A(net346),
    .Y(_1045_),
    .D(_1042_));
 sg13g2_xnor2_1 _4873_ (.Y(_0223_),
    .A(net346),
    .B(_1043_));
 sg13g2_xnor2_1 _4874_ (.Y(_0224_),
    .A(net368),
    .B(_1045_));
 sg13g2_o21ai_1 _4875_ (.B1(net987),
    .Y(_1046_),
    .A1(_3202_),
    .A2(_1045_));
 sg13g2_o21ai_1 _4876_ (.B1(_1046_),
    .Y(_0225_),
    .A1(_0547_),
    .A2(net408));
 sg13g2_nor2_1 _4877_ (.A(net971),
    .B(net975),
    .Y(_1047_));
 sg13g2_or2_1 _4878_ (.X(_1048_),
    .B(net975),
    .A(net971));
 sg13g2_or3_2 _4879_ (.A(net972),
    .B(net974),
    .C(net977),
    .X(_1049_));
 sg13g2_nand2_1 _4880_ (.Y(_1050_),
    .A(net968),
    .B(_1049_));
 sg13g2_a21oi_2 _4881_ (.B1(net967),
    .Y(_1051_),
    .A2(_1049_),
    .A1(net968));
 sg13g2_nand2_2 _4882_ (.Y(_1052_),
    .A(\vgademo.a_scrolly[10] ),
    .B(net965));
 sg13g2_nor2_1 _4883_ (.A(net940),
    .B(_1051_),
    .Y(_1053_));
 sg13g2_nor2_2 _4884_ (.A(_1051_),
    .B(_1052_),
    .Y(_1054_));
 sg13g2_nor2_2 _4885_ (.A(\vgademo.a_scrolly[12] ),
    .B(\vgademo.a_scrolly[13] ),
    .Y(_1055_));
 sg13g2_inv_1 _4886_ (.Y(_1056_),
    .A(_1055_));
 sg13g2_nor2_1 _4887_ (.A(net961),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_nand2_2 _4888_ (.Y(_1058_),
    .A(_3130_),
    .B(_1055_));
 sg13g2_nand2b_1 _4889_ (.Y(_1059_),
    .B(\vgademo.a_scrolly[3] ),
    .A_N(net977));
 sg13g2_nor3_1 _4890_ (.A(_1048_),
    .B(_1052_),
    .C(_1059_),
    .Y(_1060_));
 sg13g2_nand3b_1 _4891_ (.B(_3130_),
    .C(_0066_),
    .Y(_1061_),
    .A_N(\vgademo.a_scrolly[12] ));
 sg13g2_inv_1 _4892_ (.Y(_1062_),
    .A(_1061_));
 sg13g2_nand2b_1 _4893_ (.Y(_1063_),
    .B(net968),
    .A_N(net966));
 sg13g2_nor4_1 _4894_ (.A(_3129_),
    .B(_1049_),
    .C(_1052_),
    .D(_1063_),
    .Y(_1064_));
 sg13g2_nor2b_1 _4895_ (.A(_1061_),
    .B_N(_1064_),
    .Y(_1065_));
 sg13g2_nor2_1 _4896_ (.A(_1054_),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_nor3_2 _4897_ (.A(_1054_),
    .B(_1058_),
    .C(_1065_),
    .Y(_1067_));
 sg13g2_nor2_1 _4898_ (.A(net969),
    .B(net971),
    .Y(_1068_));
 sg13g2_nor4_2 _4899_ (.A(net969),
    .B(net972),
    .C(net974),
    .Y(_1069_),
    .D(net977));
 sg13g2_nand3_1 _4900_ (.B(_3133_),
    .C(_1069_),
    .A(net965),
    .Y(_1070_));
 sg13g2_nand2_1 _4901_ (.Y(_1071_),
    .A(net961),
    .B(net962));
 sg13g2_nor2_1 _4902_ (.A(_0065_),
    .B(_1071_),
    .Y(_1072_));
 sg13g2_nand2_1 _4903_ (.Y(_1073_),
    .A(_1070_),
    .B(_1072_));
 sg13g2_nand2b_1 _4904_ (.Y(_1074_),
    .B(net961),
    .A_N(\vgademo.a_scrolly[12] ));
 sg13g2_nor2_2 _4905_ (.A(net966),
    .B(net968),
    .Y(_1075_));
 sg13g2_nor4_1 _4906_ (.A(net967),
    .B(net968),
    .C(_3137_),
    .D(_1074_),
    .Y(_1076_));
 sg13g2_nand2_1 _4907_ (.Y(_1077_),
    .A(_1060_),
    .B(_1076_));
 sg13g2_a221oi_1 _4908_ (.B2(_1060_),
    .C1(_1056_),
    .B1(_1076_),
    .A1(_1070_),
    .Y(_1078_),
    .A2(_1072_));
 sg13g2_nand3_1 _4909_ (.B(_1073_),
    .C(_1077_),
    .A(_1055_),
    .Y(_1079_));
 sg13g2_nand2_2 _4910_ (.Y(_1080_),
    .A(net981),
    .B(net977));
 sg13g2_nand3_1 _4911_ (.B(net975),
    .C(net978),
    .A(net981),
    .Y(_1081_));
 sg13g2_nand2_1 _4912_ (.Y(_1082_),
    .A(_3134_),
    .B(_1081_));
 sg13g2_nand2b_2 _4913_ (.Y(_1083_),
    .B(net963),
    .A_N(net964));
 sg13g2_nor2_1 _4914_ (.A(_1063_),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_a21oi_1 _4915_ (.A1(_3132_),
    .A2(_3133_),
    .Y(_1085_),
    .B1(_3131_));
 sg13g2_a21oi_1 _4916_ (.A1(_1082_),
    .A2(_1084_),
    .Y(_1086_),
    .B1(_1085_));
 sg13g2_o21ai_1 _4917_ (.B1(_0067_),
    .Y(_1087_),
    .A1(_1074_),
    .A2(_1086_));
 sg13g2_and2_1 _4918_ (.A(_3137_),
    .B(_1087_),
    .X(_1088_));
 sg13g2_nand2_2 _4919_ (.Y(_1089_),
    .A(\vgademo.a_scrolly[12] ),
    .B(\vgademo.a_scrolly[13] ));
 sg13g2_nor3_1 _4920_ (.A(net966),
    .B(net968),
    .C(_1083_),
    .Y(_1090_));
 sg13g2_nand4_1 _4921_ (.B(net940),
    .C(_3134_),
    .A(net963),
    .Y(_1091_),
    .D(_1075_));
 sg13g2_nand2_1 _4922_ (.Y(_1092_),
    .A(net962),
    .B(_1091_));
 sg13g2_a221oi_1 _4923_ (.B2(net962),
    .C1(net961),
    .B1(_1091_),
    .A1(_1082_),
    .Y(_1093_),
    .A2(_1090_));
 sg13g2_or2_1 _4924_ (.X(_1094_),
    .B(_1093_),
    .A(_1089_));
 sg13g2_nand3_1 _4925_ (.B(_1087_),
    .C(_1094_),
    .A(_3137_),
    .Y(_1095_));
 sg13g2_a21oi_1 _4926_ (.A1(_1079_),
    .A2(_1095_),
    .Y(_1096_),
    .B1(_1067_));
 sg13g2_a21oi_2 _4927_ (.B1(_3115_),
    .Y(_1097_),
    .A2(_1096_),
    .A1(_0064_));
 sg13g2_and3_1 _4928_ (.X(_1098_),
    .A(_3115_),
    .B(_0064_),
    .C(_1096_));
 sg13g2_nor2_1 _4929_ (.A(_1097_),
    .B(_1098_),
    .Y(_1099_));
 sg13g2_xnor2_1 _4930_ (.Y(_1100_),
    .A(\vgademo.audio_kick_frames[0] ),
    .B(_1099_));
 sg13g2_and4_1 _4931_ (.A(_3212_),
    .B(_0578_),
    .C(_0649_),
    .D(_1100_),
    .X(_1101_));
 sg13g2_a21o_1 _4932_ (.A2(net926),
    .A1(net458),
    .B1(_1101_),
    .X(_0226_));
 sg13g2_nand2b_1 _4933_ (.Y(_1102_),
    .B(net977),
    .A_N(_1078_));
 sg13g2_nand2_1 _4934_ (.Y(_1103_),
    .A(_0069_),
    .B(_1078_));
 sg13g2_nand3b_1 _4935_ (.B(_1102_),
    .C(_1103_),
    .Y(_1104_),
    .A_N(_1067_));
 sg13g2_a21oi_2 _4936_ (.B1(_1104_),
    .Y(_1105_),
    .A2(_1095_),
    .A1(net904));
 sg13g2_xor2_1 _4937_ (.B(_1105_),
    .A(\vgademo.bayer_j[1] ),
    .X(_1106_));
 sg13g2_xnor2_1 _4938_ (.Y(_1107_),
    .A(\vgademo.bayer_j[1] ),
    .B(_1105_));
 sg13g2_xnor2_1 _4939_ (.Y(_1108_),
    .A(_0068_),
    .B(_1106_));
 sg13g2_a21o_1 _4940_ (.A2(_1099_),
    .A1(_3113_),
    .B1(_1097_),
    .X(_1109_));
 sg13g2_nand2_1 _4941_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_xor2_1 _4942_ (.B(_1109_),
    .A(_1108_),
    .X(_1111_));
 sg13g2_and2_1 _4943_ (.A(net927),
    .B(_1111_),
    .X(_1112_));
 sg13g2_a21o_1 _4944_ (.A2(net926),
    .A1(net391),
    .B1(_1112_),
    .X(_0227_));
 sg13g2_nor2_1 _4945_ (.A(_0072_),
    .B(_1105_),
    .Y(_1113_));
 sg13g2_a21oi_1 _4946_ (.A1(_0068_),
    .A2(_1107_),
    .Y(_1114_),
    .B1(_1113_));
 sg13g2_xor2_1 _4947_ (.B(net977),
    .A(net974),
    .X(_1115_));
 sg13g2_nand2_1 _4948_ (.Y(_1116_),
    .A(_1078_),
    .B(_1115_));
 sg13g2_nand2_1 _4949_ (.Y(_1117_),
    .A(_3135_),
    .B(_1079_));
 sg13g2_a221oi_1 _4950_ (.B2(_1117_),
    .C1(_1067_),
    .B1(_1116_),
    .A1(net904),
    .Y(_1118_),
    .A2(_1095_));
 sg13g2_xnor2_1 _4951_ (.Y(_1119_),
    .A(_0071_),
    .B(_1118_));
 sg13g2_nor2b_1 _4952_ (.A(_1114_),
    .B_N(_1119_),
    .Y(_1120_));
 sg13g2_xor2_1 _4953_ (.B(_1119_),
    .A(_1114_),
    .X(_1121_));
 sg13g2_inv_1 _4954_ (.Y(_1122_),
    .A(_1121_));
 sg13g2_xnor2_1 _4955_ (.Y(_1123_),
    .A(_3114_),
    .B(_1121_));
 sg13g2_nor2_1 _4956_ (.A(_1110_),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_xor2_1 _4957_ (.B(_1123_),
    .A(_1110_),
    .X(_1125_));
 sg13g2_mux2_1 _4958_ (.A0(net302),
    .A1(_1125_),
    .S(net927),
    .X(_0228_));
 sg13g2_nor2_1 _4959_ (.A(net357),
    .B(net927),
    .Y(_1126_));
 sg13g2_nand2_1 _4960_ (.Y(_1127_),
    .A(_3116_),
    .B(_1118_));
 sg13g2_o21ai_1 _4961_ (.B1(net972),
    .Y(_1128_),
    .A1(net975),
    .A2(net977));
 sg13g2_nand2_1 _4962_ (.Y(_1129_),
    .A(_1049_),
    .B(_1128_));
 sg13g2_mux2_1 _4963_ (.A0(_0075_),
    .A1(_1129_),
    .S(_1078_),
    .X(_1130_));
 sg13g2_a221oi_1 _4964_ (.B2(_1095_),
    .C1(_1130_),
    .B1(_1079_),
    .A1(_1057_),
    .Y(_1131_),
    .A2(_1066_));
 sg13g2_nand2_1 _4965_ (.Y(_1132_),
    .A(_0074_),
    .B(_1131_));
 sg13g2_xnor2_1 _4966_ (.Y(_1133_),
    .A(_0074_),
    .B(_1131_));
 sg13g2_nand2_1 _4967_ (.Y(_1134_),
    .A(_1127_),
    .B(_1133_));
 sg13g2_nor2_1 _4968_ (.A(_1127_),
    .B(_1133_),
    .Y(_1135_));
 sg13g2_xnor2_1 _4969_ (.Y(_1136_),
    .A(_1127_),
    .B(_1133_));
 sg13g2_a21oi_1 _4970_ (.A1(_0060_),
    .A2(_1122_),
    .Y(_1137_),
    .B1(_1120_));
 sg13g2_nor2_1 _4971_ (.A(_1136_),
    .B(_1137_),
    .Y(_1138_));
 sg13g2_xor2_1 _4972_ (.B(_1137_),
    .A(_1136_),
    .X(_1139_));
 sg13g2_xnor2_1 _4973_ (.Y(_1140_),
    .A(_1124_),
    .B(_1139_));
 sg13g2_a21oi_1 _4974_ (.A1(net927),
    .A2(_1140_),
    .Y(_0229_),
    .B1(_1126_));
 sg13g2_a21oi_1 _4975_ (.A1(_1124_),
    .A2(_1139_),
    .Y(_1141_),
    .B1(_1138_));
 sg13g2_and3_1 _4976_ (.X(_1142_),
    .A(_3137_),
    .B(net904),
    .C(_1087_));
 sg13g2_nand2_1 _4977_ (.Y(_1143_),
    .A(net969),
    .B(net971));
 sg13g2_nand3b_1 _4978_ (.B(_1094_),
    .C(_1143_),
    .Y(_1144_),
    .A_N(_1068_));
 sg13g2_nand2_2 _4979_ (.Y(_1145_),
    .A(_0069_),
    .B(_1047_));
 sg13g2_xnor2_1 _4980_ (.Y(_1146_),
    .A(_0078_),
    .B(_1145_));
 sg13g2_a221oi_1 _4981_ (.B2(_1078_),
    .C1(_1067_),
    .B1(_1146_),
    .A1(_1142_),
    .Y(_1147_),
    .A2(_1144_));
 sg13g2_nand2_1 _4982_ (.Y(_1148_),
    .A(_0077_),
    .B(_1147_));
 sg13g2_xnor2_1 _4983_ (.Y(_1149_),
    .A(_0077_),
    .B(_1147_));
 sg13g2_nand2_1 _4984_ (.Y(_1150_),
    .A(_1132_),
    .B(_1149_));
 sg13g2_xor2_1 _4985_ (.B(_1149_),
    .A(_1132_),
    .X(_1151_));
 sg13g2_inv_1 _4986_ (.Y(_1152_),
    .A(_1151_));
 sg13g2_xnor2_1 _4987_ (.Y(_1153_),
    .A(_1134_),
    .B(_1151_));
 sg13g2_nand2b_1 _4988_ (.Y(_1154_),
    .B(_1153_),
    .A_N(_1141_));
 sg13g2_xnor2_1 _4989_ (.Y(_1155_),
    .A(_1141_),
    .B(_1153_));
 sg13g2_mux2_1 _4990_ (.A0(net303),
    .A1(_1155_),
    .S(net927),
    .X(_0230_));
 sg13g2_nor2_1 _4991_ (.A(net355),
    .B(net928),
    .Y(_1156_));
 sg13g2_o21ai_1 _4992_ (.B1(_1154_),
    .Y(_1157_),
    .A1(_1134_),
    .A2(_1152_));
 sg13g2_xor2_1 _4993_ (.B(_1068_),
    .A(_0080_),
    .X(_1158_));
 sg13g2_o21ai_1 _4994_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_1089_),
    .A2(_1093_));
 sg13g2_nand4_1 _4995_ (.B(net904),
    .C(_1087_),
    .A(_3137_),
    .Y(_1160_),
    .D(_1159_));
 sg13g2_nand2_1 _4996_ (.Y(_1161_),
    .A(net970),
    .B(_1145_));
 sg13g2_xor2_1 _4997_ (.B(_1161_),
    .A(_0080_),
    .X(_1162_));
 sg13g2_nand2_1 _4998_ (.Y(_1163_),
    .A(_1078_),
    .B(_1162_));
 sg13g2_a21oi_2 _4999_ (.B1(_1067_),
    .Y(_1164_),
    .A2(_1163_),
    .A1(_1160_));
 sg13g2_and2_1 _5000_ (.A(net959),
    .B(_1164_),
    .X(_1165_));
 sg13g2_or2_1 _5001_ (.X(_1166_),
    .B(_1164_),
    .A(net959));
 sg13g2_nor2b_1 _5002_ (.A(_1165_),
    .B_N(_1166_),
    .Y(_1167_));
 sg13g2_nand2b_1 _5003_ (.Y(_1168_),
    .B(_1167_),
    .A_N(_1148_));
 sg13g2_xor2_1 _5004_ (.B(_1167_),
    .A(_1148_),
    .X(_1169_));
 sg13g2_inv_1 _5005_ (.Y(_1170_),
    .A(_1169_));
 sg13g2_xor2_1 _5006_ (.B(_1169_),
    .A(_1150_),
    .X(_1171_));
 sg13g2_nand2b_1 _5007_ (.Y(_1172_),
    .B(_1157_),
    .A_N(_1171_));
 sg13g2_xor2_1 _5008_ (.B(_1171_),
    .A(_1157_),
    .X(_1173_));
 sg13g2_a21oi_1 _5009_ (.A1(net927),
    .A2(_1173_),
    .Y(_0231_),
    .B1(_1156_));
 sg13g2_nor2_1 _5010_ (.A(net312),
    .B(net928),
    .Y(_1174_));
 sg13g2_o21ai_1 _5011_ (.B1(_1172_),
    .Y(_1175_),
    .A1(_1150_),
    .A2(_1170_));
 sg13g2_nor2_1 _5012_ (.A(_3128_),
    .B(_1164_),
    .Y(_1176_));
 sg13g2_a21oi_1 _5013_ (.A1(_0075_),
    .A2(_1075_),
    .Y(_1177_),
    .B1(_3132_));
 sg13g2_nand3_1 _5014_ (.B(_0075_),
    .C(_1075_),
    .A(_3132_),
    .Y(_1178_));
 sg13g2_nor2b_1 _5015_ (.A(_1177_),
    .B_N(_1178_),
    .Y(_1179_));
 sg13g2_o21ai_1 _5016_ (.B1(_1179_),
    .Y(_1180_),
    .A1(_1089_),
    .A2(_1093_));
 sg13g2_nand4_1 _5017_ (.B(net904),
    .C(_1087_),
    .A(_3137_),
    .Y(_1181_),
    .D(_1180_));
 sg13g2_nand3_1 _5018_ (.B(net969),
    .C(_1145_),
    .A(net966),
    .Y(_1182_));
 sg13g2_xnor2_1 _5019_ (.Y(_1183_),
    .A(net940),
    .B(_1182_));
 sg13g2_nand2_1 _5020_ (.Y(_1184_),
    .A(_1078_),
    .B(_1183_));
 sg13g2_a21oi_2 _5021_ (.B1(_1067_),
    .Y(_1185_),
    .A2(_1184_),
    .A1(_1181_));
 sg13g2_xnor2_1 _5022_ (.Y(_1186_),
    .A(net958),
    .B(_1185_));
 sg13g2_nand2b_1 _5023_ (.Y(_1187_),
    .B(_1186_),
    .A_N(_1176_));
 sg13g2_xnor2_1 _5024_ (.Y(_1188_),
    .A(_1176_),
    .B(_1186_));
 sg13g2_xnor2_1 _5025_ (.Y(_1189_),
    .A(_1168_),
    .B(_1188_));
 sg13g2_nor2b_1 _5026_ (.A(_1189_),
    .B_N(_1175_),
    .Y(_1190_));
 sg13g2_xor2_1 _5027_ (.B(_1189_),
    .A(_1175_),
    .X(_1191_));
 sg13g2_a21oi_1 _5028_ (.A1(net927),
    .A2(_1191_),
    .Y(_0232_),
    .B1(_1174_));
 sg13g2_a21o_1 _5029_ (.A2(_1188_),
    .A1(_1168_),
    .B1(_1190_),
    .X(_1192_));
 sg13g2_xor2_1 _5030_ (.B(_1178_),
    .A(_0015_),
    .X(_1193_));
 sg13g2_o21ai_1 _5031_ (.B1(_1193_),
    .Y(_1194_),
    .A1(_1089_),
    .A2(_1093_));
 sg13g2_nand3_1 _5032_ (.B(_1087_),
    .C(_1194_),
    .A(_3137_),
    .Y(_1195_));
 sg13g2_a21oi_1 _5033_ (.A1(_0065_),
    .A2(_1182_),
    .Y(_1196_),
    .B1(net962));
 sg13g2_nand3_1 _5034_ (.B(_0065_),
    .C(_1182_),
    .A(net962),
    .Y(_1197_));
 sg13g2_nor2_1 _5035_ (.A(net904),
    .B(_1196_),
    .Y(_1198_));
 sg13g2_a221oi_1 _5036_ (.B2(_1198_),
    .C1(_1067_),
    .B1(_1197_),
    .A1(net904),
    .Y(_1199_),
    .A2(_1195_));
 sg13g2_nand2b_1 _5037_ (.Y(_1200_),
    .B(_0014_),
    .A_N(_1199_));
 sg13g2_xnor2_1 _5038_ (.Y(_1201_),
    .A(_0014_),
    .B(_1199_));
 sg13g2_nor2b_1 _5039_ (.A(_1185_),
    .B_N(_0016_),
    .Y(_1202_));
 sg13g2_nor2_1 _5040_ (.A(_1201_),
    .B(_1202_),
    .Y(_1203_));
 sg13g2_xnor2_1 _5041_ (.Y(_1204_),
    .A(_1201_),
    .B(_1202_));
 sg13g2_nor2_1 _5042_ (.A(_1187_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_xor2_1 _5043_ (.B(_1204_),
    .A(_1187_),
    .X(_1206_));
 sg13g2_xor2_1 _5044_ (.B(_1206_),
    .A(_1192_),
    .X(_1207_));
 sg13g2_mux2_1 _5045_ (.A0(net293),
    .A1(_1207_),
    .S(net928),
    .X(_0233_));
 sg13g2_a21oi_1 _5046_ (.A1(_1192_),
    .A2(_1206_),
    .Y(_1208_),
    .B1(_1205_));
 sg13g2_xor2_1 _5047_ (.B(_1092_),
    .A(_0019_),
    .X(_1209_));
 sg13g2_a21oi_1 _5048_ (.A1(net940),
    .A2(_1182_),
    .Y(_1210_),
    .B1(_1071_));
 sg13g2_nand3_1 _5049_ (.B(_1142_),
    .C(_1209_),
    .A(_1094_),
    .Y(_1211_));
 sg13g2_o21ai_1 _5050_ (.B1(_1211_),
    .Y(_1212_),
    .A1(net904),
    .A2(_1210_));
 sg13g2_xnor2_1 _5051_ (.Y(_1213_),
    .A(_0018_),
    .B(_1212_));
 sg13g2_xnor2_1 _5052_ (.Y(_1214_),
    .A(_1200_),
    .B(_1213_));
 sg13g2_xnor2_1 _5053_ (.Y(_1215_),
    .A(_1203_),
    .B(_1214_));
 sg13g2_xnor2_1 _5054_ (.Y(_1216_),
    .A(_1208_),
    .B(_1215_));
 sg13g2_and2_1 _5055_ (.A(net928),
    .B(_1216_),
    .X(_1217_));
 sg13g2_a21o_1 _5056_ (.A2(net926),
    .A1(net314),
    .B1(_1217_),
    .X(_0234_));
 sg13g2_nor2_1 _5057_ (.A(\vgademo.a_scrolly[3] ),
    .B(net977),
    .Y(_1218_));
 sg13g2_nand2_2 _5058_ (.Y(_1219_),
    .A(_3129_),
    .B(_3136_));
 sg13g2_nor2_2 _5059_ (.A(\vgademo.a_scrolly[10] ),
    .B(net965),
    .Y(_1220_));
 sg13g2_nand2_1 _5060_ (.Y(_1221_),
    .A(_3133_),
    .B(_1220_));
 sg13g2_nand2_2 _5061_ (.Y(_1222_),
    .A(net971),
    .B(net974));
 sg13g2_a21oi_1 _5062_ (.A1(net972),
    .A2(_1219_),
    .Y(_1223_),
    .B1(_1061_));
 sg13g2_nand4_1 _5063_ (.B(_1220_),
    .C(_1222_),
    .A(_1075_),
    .Y(_1224_),
    .D(_1223_));
 sg13g2_nor3_1 _5064_ (.A(\vgademo.audio_songpos[6] ),
    .B(net1018),
    .C(_3270_),
    .Y(_1225_));
 sg13g2_nand4_1 _5065_ (.B(_3295_),
    .C(_1224_),
    .A(_3280_),
    .Y(_1226_),
    .D(_1225_));
 sg13g2_nand2_2 _5066_ (.Y(_1227_),
    .A(net920),
    .B(_1226_));
 sg13g2_a21oi_1 _5067_ (.A1(net920),
    .A2(_1226_),
    .Y(_1228_),
    .B1(net980));
 sg13g2_a21oi_1 _5068_ (.A1(net980),
    .A2(net920),
    .Y(_0235_),
    .B1(_1228_));
 sg13g2_nand2_1 _5069_ (.Y(_1229_),
    .A(net978),
    .B(net915));
 sg13g2_nand2_1 _5070_ (.Y(_1230_),
    .A(_1080_),
    .B(_1219_));
 sg13g2_o21ai_1 _5071_ (.B1(_1229_),
    .Y(_0236_),
    .A1(_1227_),
    .A2(_1230_));
 sg13g2_nand2_1 _5072_ (.Y(_1231_),
    .A(net974),
    .B(net915));
 sg13g2_xnor2_1 _5073_ (.Y(_1232_),
    .A(_3135_),
    .B(_1080_));
 sg13g2_o21ai_1 _5074_ (.B1(_1231_),
    .Y(_0237_),
    .A1(_1227_),
    .A2(_1232_));
 sg13g2_nand2_1 _5075_ (.Y(_1233_),
    .A(net971),
    .B(net909));
 sg13g2_xnor2_1 _5076_ (.Y(_1234_),
    .A(net581),
    .B(_1081_));
 sg13g2_o21ai_1 _5077_ (.B1(_1233_),
    .Y(_0238_),
    .A1(net884),
    .A2(_1234_));
 sg13g2_nand2_1 _5078_ (.Y(_1235_),
    .A(net968),
    .B(net909));
 sg13g2_xnor2_1 _5079_ (.Y(_1236_),
    .A(_3140_),
    .B(_1222_));
 sg13g2_nand2_1 _5080_ (.Y(_1237_),
    .A(net584),
    .B(_1080_));
 sg13g2_o21ai_1 _5081_ (.B1(_1237_),
    .Y(_1238_),
    .A1(_1080_),
    .A2(_1236_));
 sg13g2_o21ai_1 _5082_ (.B1(_1235_),
    .Y(_0239_),
    .A1(net884),
    .A2(_1238_));
 sg13g2_nand2_1 _5083_ (.Y(_1239_),
    .A(net967),
    .B(net909));
 sg13g2_nor3_2 _5084_ (.A(_0078_),
    .B(_1080_),
    .C(_1222_),
    .Y(_1240_));
 sg13g2_xor2_1 _5085_ (.B(_1240_),
    .A(_0080_),
    .X(_1241_));
 sg13g2_o21ai_1 _5086_ (.B1(_1239_),
    .Y(_0240_),
    .A1(net884),
    .A2(_1241_));
 sg13g2_nand2_1 _5087_ (.Y(_1242_),
    .A(net964),
    .B(net909));
 sg13g2_or3_2 _5088_ (.A(_3133_),
    .B(_1081_),
    .C(_1143_),
    .X(_1243_));
 sg13g2_nor2_1 _5089_ (.A(_0065_),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_xnor2_1 _5090_ (.Y(_1245_),
    .A(net503),
    .B(_1243_));
 sg13g2_o21ai_1 _5091_ (.B1(_1242_),
    .Y(_0241_),
    .A1(net884),
    .A2(_1245_));
 sg13g2_nand2_1 _5092_ (.Y(_1246_),
    .A(net963),
    .B(net909));
 sg13g2_xor2_1 _5093_ (.B(_1244_),
    .A(net422),
    .X(_1247_));
 sg13g2_o21ai_1 _5094_ (.B1(_1246_),
    .Y(_0242_),
    .A1(net884),
    .A2(net423));
 sg13g2_nand2_1 _5095_ (.Y(_1248_),
    .A(net238),
    .B(net909));
 sg13g2_nor2_2 _5096_ (.A(_1052_),
    .B(_1243_),
    .Y(_1249_));
 sg13g2_nand2b_1 _5097_ (.Y(_1250_),
    .B(_1249_),
    .A_N(_0019_));
 sg13g2_xor2_1 _5098_ (.B(_1249_),
    .A(_0019_),
    .X(_1251_));
 sg13g2_o21ai_1 _5099_ (.B1(_1248_),
    .Y(_0243_),
    .A1(net884),
    .A2(_1251_));
 sg13g2_nand2_1 _5100_ (.Y(_1252_),
    .A(\vgademo.a_scrolly[12] ),
    .B(net909));
 sg13g2_xnor2_1 _5101_ (.Y(_1253_),
    .A(net536),
    .B(_1250_));
 sg13g2_o21ai_1 _5102_ (.B1(_1252_),
    .Y(_0244_),
    .A1(net884),
    .A2(_1253_));
 sg13g2_nand2_1 _5103_ (.Y(_1254_),
    .A(net403),
    .B(net909));
 sg13g2_nand3_1 _5104_ (.B(net961),
    .C(_1249_),
    .A(\vgademo.a_scrolly[12] ),
    .Y(_1255_));
 sg13g2_xnor2_1 _5105_ (.Y(_1256_),
    .A(_0066_),
    .B(_1255_));
 sg13g2_o21ai_1 _5106_ (.B1(_1254_),
    .Y(_0245_),
    .A1(net884),
    .A2(_1256_));
 sg13g2_nand2_2 _5107_ (.Y(_1257_),
    .A(_3215_),
    .B(_0587_));
 sg13g2_a21oi_1 _5108_ (.A1(_3215_),
    .A2(_0587_),
    .Y(_1258_),
    .B1(net582));
 sg13g2_nand2_1 _5109_ (.Y(_1259_),
    .A(\vgademo.bayer_j[0] ),
    .B(_3215_));
 sg13g2_nor2b_1 _5110_ (.A(net583),
    .B_N(_1259_),
    .Y(_0246_));
 sg13g2_xnor2_1 _5111_ (.Y(_0247_),
    .A(\vgademo.bayer_j[1] ),
    .B(_1259_));
 sg13g2_nand2_1 _5112_ (.Y(_1260_),
    .A(net462),
    .B(net931));
 sg13g2_nand2_2 _5113_ (.Y(_1261_),
    .A(\vgademo.bayer_j[1] ),
    .B(\vgademo.bayer_j[0] ));
 sg13g2_nor2_1 _5114_ (.A(_0071_),
    .B(_1261_),
    .Y(_1262_));
 sg13g2_xnor2_1 _5115_ (.Y(_1263_),
    .A(_0071_),
    .B(_1261_));
 sg13g2_o21ai_1 _5116_ (.B1(_1260_),
    .Y(_0248_),
    .A1(_1257_),
    .A2(_1263_));
 sg13g2_nand2_1 _5117_ (.Y(_1264_),
    .A(net542),
    .B(net931));
 sg13g2_xor2_1 _5118_ (.B(_1262_),
    .A(_0074_),
    .X(_1265_));
 sg13g2_o21ai_1 _5119_ (.B1(_1264_),
    .Y(_0249_),
    .A1(_1257_),
    .A2(_1265_));
 sg13g2_nand2_1 _5120_ (.Y(_1266_),
    .A(net265),
    .B(net930));
 sg13g2_nor2_1 _5121_ (.A(_3243_),
    .B(_1261_),
    .Y(_1267_));
 sg13g2_nor3_1 _5122_ (.A(_0077_),
    .B(_3243_),
    .C(_1261_),
    .Y(_1268_));
 sg13g2_xor2_1 _5123_ (.B(_1267_),
    .A(_0077_),
    .X(_1269_));
 sg13g2_o21ai_1 _5124_ (.B1(_1266_),
    .Y(_0250_),
    .A1(_1257_),
    .A2(_1269_));
 sg13g2_nand2_1 _5125_ (.Y(_1270_),
    .A(net305),
    .B(net930));
 sg13g2_xnor2_1 _5126_ (.Y(_1271_),
    .A(_3128_),
    .B(_1268_));
 sg13g2_o21ai_1 _5127_ (.B1(_1270_),
    .Y(_0251_),
    .A1(_1257_),
    .A2(_1271_));
 sg13g2_nand2_1 _5128_ (.Y(_1272_),
    .A(net958),
    .B(net930));
 sg13g2_nand3_1 _5129_ (.B(\vgademo.v_count[5] ),
    .C(_1267_),
    .A(net265),
    .Y(_1273_));
 sg13g2_nor2_1 _5130_ (.A(_0016_),
    .B(_1273_),
    .Y(_1274_));
 sg13g2_xnor2_1 _5131_ (.Y(_1275_),
    .A(_0016_),
    .B(_1273_));
 sg13g2_o21ai_1 _5132_ (.B1(_1272_),
    .Y(_0252_),
    .A1(_1257_),
    .A2(_1275_));
 sg13g2_nand2_1 _5133_ (.Y(_1276_),
    .A(net957),
    .B(net930));
 sg13g2_xor2_1 _5134_ (.B(_1274_),
    .A(net476),
    .X(_1277_));
 sg13g2_o21ai_1 _5135_ (.B1(_1276_),
    .Y(_0253_),
    .A1(_1257_),
    .A2(net477));
 sg13g2_nand2_1 _5136_ (.Y(_1278_),
    .A(net530),
    .B(net931));
 sg13g2_o21ai_1 _5137_ (.B1(_0018_),
    .Y(_1279_),
    .A1(_3238_),
    .A2(_1273_));
 sg13g2_nor3_1 _5138_ (.A(_0018_),
    .B(_3238_),
    .C(_1273_),
    .Y(_1280_));
 sg13g2_nand2b_1 _5139_ (.Y(_1281_),
    .B(_1279_),
    .A_N(_1257_));
 sg13g2_o21ai_1 _5140_ (.B1(_1278_),
    .Y(_0254_),
    .A1(_1280_),
    .A2(_1281_));
 sg13g2_nand2_1 _5141_ (.Y(_1282_),
    .A(net955),
    .B(net931));
 sg13g2_xor2_1 _5142_ (.B(_1280_),
    .A(net412),
    .X(_1283_));
 sg13g2_o21ai_1 _5143_ (.B1(_1282_),
    .Y(_0255_),
    .A1(_1257_),
    .A2(net413));
 sg13g2_nor2_1 _5144_ (.A(\vgademo.scanline_audio_sample[3] ),
    .B(\vgademo.scanline_audio_sample[4] ),
    .Y(_1284_));
 sg13g2_nand2_1 _5145_ (.Y(_1285_),
    .A(_0043_),
    .B(_1284_));
 sg13g2_xnor2_1 _5146_ (.Y(_1286_),
    .A(\vgademo.scanline_audio_sample[6] ),
    .B(_1285_));
 sg13g2_xor2_1 _5147_ (.B(_1286_),
    .A(_0036_),
    .X(_1287_));
 sg13g2_nand2_1 _5148_ (.Y(_1288_),
    .A(_0037_),
    .B(_1287_));
 sg13g2_xnor2_1 _5149_ (.Y(_1289_),
    .A(_0043_),
    .B(_1284_));
 sg13g2_xnor2_1 _5150_ (.Y(_1290_),
    .A(_0035_),
    .B(_1289_));
 sg13g2_xnor2_1 _5151_ (.Y(_1291_),
    .A(\vgademo.scanline_audio_sample[3] ),
    .B(\vgademo.scanline_audio_sample[4] ));
 sg13g2_nand2_1 _5152_ (.Y(_1292_),
    .A(_0044_),
    .B(_1291_));
 sg13g2_xnor2_1 _5153_ (.Y(_1293_),
    .A(_0044_),
    .B(_1291_));
 sg13g2_nor3_1 _5154_ (.A(_1288_),
    .B(_1290_),
    .C(_1293_),
    .Y(_1294_));
 sg13g2_nor2b_1 _5155_ (.A(net986),
    .B_N(\vgademo.scanline_audio_sample[1] ),
    .Y(_1295_));
 sg13g2_nand2_1 _5156_ (.Y(_1296_),
    .A(_3119_),
    .B(\vgademo.scanline_audio_sample[1] ));
 sg13g2_nor2_1 _5157_ (.A(_3120_),
    .B(\vgademo.scanline_audio_sample[0] ),
    .Y(_1297_));
 sg13g2_nor2_1 _5158_ (.A(_3119_),
    .B(\vgademo.scanline_audio_sample[1] ),
    .Y(_1298_));
 sg13g2_o21ai_1 _5159_ (.B1(_1296_),
    .Y(_1299_),
    .A1(_1297_),
    .A2(_1298_));
 sg13g2_nor2_1 _5160_ (.A(_3121_),
    .B(\vgademo.scanline_audio_sample[3] ),
    .Y(_1300_));
 sg13g2_nand2_1 _5161_ (.Y(_1301_),
    .A(_3121_),
    .B(\vgademo.scanline_audio_sample[3] ));
 sg13g2_nor2b_1 _5162_ (.A(_1300_),
    .B_N(_1301_),
    .Y(_1302_));
 sg13g2_inv_1 _5163_ (.Y(_1303_),
    .A(_1302_));
 sg13g2_nand2_1 _5164_ (.Y(_1304_),
    .A(_3122_),
    .B(\vgademo.scanline_audio_sample[2] ));
 sg13g2_xor2_1 _5165_ (.B(\vgademo.scanline_audio_sample[2] ),
    .A(\vgademo.h_count[2] ),
    .X(_1305_));
 sg13g2_nor2_1 _5166_ (.A(_1302_),
    .B(_1305_),
    .Y(_1306_));
 sg13g2_a22oi_1 _5167_ (.Y(_1307_),
    .B1(_1299_),
    .B2(_1306_),
    .A2(_3209_),
    .A1(_3121_));
 sg13g2_o21ai_1 _5168_ (.B1(_1307_),
    .Y(_1308_),
    .A1(_1302_),
    .A2(_1304_));
 sg13g2_nor2_1 _5169_ (.A(_1290_),
    .B(_1292_),
    .Y(_1309_));
 sg13g2_a21oi_1 _5170_ (.A1(net941),
    .A2(_1289_),
    .Y(_1310_),
    .B1(_1309_));
 sg13g2_nor2_1 _5171_ (.A(\vgademo.h_count[7] ),
    .B(net984),
    .Y(_1311_));
 sg13g2_a22oi_1 _5172_ (.Y(_1312_),
    .B1(_1311_),
    .B2(_1286_),
    .A2(_1308_),
    .A1(_1294_));
 sg13g2_o21ai_1 _5173_ (.B1(_1312_),
    .Y(_1313_),
    .A1(_1288_),
    .A2(_1310_));
 sg13g2_nor2b_1 _5174_ (.A(net984),
    .B_N(\vgademo.scanline_audio_sample[6] ),
    .Y(_1314_));
 sg13g2_nor2b_1 _5175_ (.A(\vgademo.scanline_audio_sample[6] ),
    .B_N(net984),
    .Y(_1315_));
 sg13g2_o21ai_1 _5176_ (.B1(_0037_),
    .Y(_1316_),
    .A1(net941),
    .A2(\vgademo.scanline_audio_sample[5] ));
 sg13g2_or3_1 _5177_ (.A(_1314_),
    .B(_1315_),
    .C(_1316_),
    .X(_1317_));
 sg13g2_a22oi_1 _5178_ (.Y(_1318_),
    .B1(\vgademo.scanline_audio_sample[4] ),
    .B2(_3123_),
    .A2(\vgademo.scanline_audio_sample[5] ),
    .A1(net941));
 sg13g2_o21ai_1 _5179_ (.B1(_1318_),
    .Y(_1319_),
    .A1(_3123_),
    .A2(\vgademo.scanline_audio_sample[4] ));
 sg13g2_nor4_1 _5180_ (.A(_1303_),
    .B(_1305_),
    .C(_1317_),
    .D(_1319_),
    .Y(_1320_));
 sg13g2_and2_1 _5181_ (.A(_1301_),
    .B(_1304_),
    .X(_1321_));
 sg13g2_nor4_1 _5182_ (.A(_1300_),
    .B(_1317_),
    .C(_1319_),
    .D(_1321_),
    .Y(_1322_));
 sg13g2_a221oi_1 _5183_ (.B2(_1299_),
    .C1(_1322_),
    .B1(_1320_),
    .A1(_3125_),
    .Y(_1323_),
    .A2(_1314_));
 sg13g2_o21ai_1 _5184_ (.B1(_1323_),
    .Y(_1324_),
    .A1(_1317_),
    .A2(_1318_));
 sg13g2_nor2b_1 _5185_ (.A(\vgademo.h_count[0] ),
    .B_N(\vgademo.scanline_audio_sample[0] ),
    .Y(_1325_));
 sg13g2_nor4_2 _5186_ (.A(_1295_),
    .B(_1297_),
    .C(_1298_),
    .Y(_1326_),
    .D(_1325_));
 sg13g2_nand2_1 _5187_ (.Y(_1327_),
    .A(_1320_),
    .B(_1326_));
 sg13g2_and4_2 _5188_ (.A(net982),
    .B(_0577_),
    .C(_1324_),
    .D(_1327_),
    .X(_1328_));
 sg13g2_nand4_1 _5189_ (.B(_0577_),
    .C(_1324_),
    .A(net982),
    .Y(_1329_),
    .D(_1327_));
 sg13g2_nand3_1 _5190_ (.B(_1306_),
    .C(_1326_),
    .A(_1294_),
    .Y(_1330_));
 sg13g2_nand3_1 _5191_ (.B(_1328_),
    .C(_1330_),
    .A(_1313_),
    .Y(_1331_));
 sg13g2_inv_2 _5192_ (.Y(_1332_),
    .A(_1331_));
 sg13g2_nor2_1 _5193_ (.A(\vgademo.v_count[8] ),
    .B(net955),
    .Y(_1333_));
 sg13g2_and2_1 _5194_ (.A(_1212_),
    .B(_1333_),
    .X(_1334_));
 sg13g2_nor2b_1 _5195_ (.A(_1186_),
    .B_N(_1201_),
    .Y(_1335_));
 sg13g2_nand3b_1 _5196_ (.B(_1167_),
    .C(_1335_),
    .Y(_1336_),
    .A_N(_1149_));
 sg13g2_inv_1 _5197_ (.Y(_1337_),
    .A(_1336_));
 sg13g2_xnor2_1 _5198_ (.Y(_1338_),
    .A(_3116_),
    .B(_1118_));
 sg13g2_nor2_1 _5199_ (.A(_1133_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_nand2_1 _5200_ (.Y(_1340_),
    .A(_0072_),
    .B(_1105_));
 sg13g2_o21ai_1 _5201_ (.B1(_1340_),
    .Y(_1341_),
    .A1(_1097_),
    .A2(_1106_));
 sg13g2_a221oi_1 _5202_ (.B2(_1341_),
    .C1(_1135_),
    .B1(_1339_),
    .A1(_3117_),
    .Y(_1342_),
    .A2(_1131_));
 sg13g2_nor2_1 _5203_ (.A(net957),
    .B(_1199_),
    .Y(_1343_));
 sg13g2_nand2b_1 _5204_ (.Y(_1344_),
    .B(_1147_),
    .A_N(net960));
 sg13g2_a21oi_1 _5205_ (.A1(_1166_),
    .A2(_1344_),
    .Y(_1345_),
    .B1(_1165_));
 sg13g2_a221oi_1 _5206_ (.B2(_1345_),
    .C1(_1343_),
    .B1(_1335_),
    .A1(_1201_),
    .Y(_1346_),
    .A2(_1202_));
 sg13g2_o21ai_1 _5207_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1336_),
    .A2(_1342_));
 sg13g2_nor2_2 _5208_ (.A(net955),
    .B(_1213_),
    .Y(_1348_));
 sg13g2_a21oi_2 _5209_ (.B1(_1334_),
    .Y(_1349_),
    .A2(_1348_),
    .A1(_1347_));
 sg13g2_a21o_1 _5210_ (.A2(_1348_),
    .A1(_1347_),
    .B1(_1334_),
    .X(_1350_));
 sg13g2_nor3_1 _5211_ (.A(_1097_),
    .B(_1098_),
    .C(_1106_),
    .Y(_1351_));
 sg13g2_and4_2 _5212_ (.A(_1337_),
    .B(_1339_),
    .C(_1348_),
    .D(_1351_),
    .X(_1352_));
 sg13g2_nand4_1 _5213_ (.B(_1339_),
    .C(_1348_),
    .A(_1337_),
    .Y(_1353_),
    .D(_1351_));
 sg13g2_nor2_2 _5214_ (.A(_1349_),
    .B(_1352_),
    .Y(_1354_));
 sg13g2_nand2_1 _5215_ (.Y(_1355_),
    .A(net856),
    .B(net854));
 sg13g2_mux2_1 _5216_ (.A0(_0074_),
    .A1(_0051_),
    .S(net851),
    .X(_1356_));
 sg13g2_nor2_1 _5217_ (.A(\vgademo.b_cos[8] ),
    .B(_1356_),
    .Y(_1357_));
 sg13g2_mux2_1 _5218_ (.A0(_0071_),
    .A1(_0049_),
    .S(net851),
    .X(_1358_));
 sg13g2_xnor2_1 _5219_ (.Y(_1359_),
    .A(_3160_),
    .B(_1358_));
 sg13g2_nor2b_1 _5220_ (.A(\vgademo.bayer_j[0] ),
    .B_N(\vgademo.b_cos[5] ),
    .Y(_1360_));
 sg13g2_nor2_1 _5221_ (.A(net954),
    .B(_1360_),
    .Y(_1361_));
 sg13g2_a21oi_1 _5222_ (.A1(net954),
    .A2(_1360_),
    .Y(_1362_),
    .B1(_0072_));
 sg13g2_nor3_1 _5223_ (.A(net850),
    .B(_1361_),
    .C(_1362_),
    .Y(_1363_));
 sg13g2_nor2b_2 _5224_ (.A(\vgademo.plane_du[2] ),
    .B_N(\vgademo.b_cos[5] ),
    .Y(_1364_));
 sg13g2_nand2_1 _5225_ (.Y(_1365_),
    .A(\vgademo.b_cos[6] ),
    .B(_1364_));
 sg13g2_nor2_1 _5226_ (.A(\vgademo.b_cos[6] ),
    .B(_1364_),
    .Y(_1366_));
 sg13g2_o21ai_1 _5227_ (.B1(_0050_),
    .Y(_1367_),
    .A1(net954),
    .A2(_1364_));
 sg13g2_a21oi_1 _5228_ (.A1(_1365_),
    .A2(_1367_),
    .Y(_1368_),
    .B1(_1354_));
 sg13g2_or2_1 _5229_ (.X(_1369_),
    .B(_1368_),
    .A(_1363_));
 sg13g2_inv_1 _5230_ (.Y(_1370_),
    .A(_1369_));
 sg13g2_nand2_1 _5231_ (.Y(_1371_),
    .A(_1359_),
    .B(_1370_));
 sg13g2_o21ai_1 _5232_ (.B1(_1371_),
    .Y(_1372_),
    .A1(\vgademo.b_cos[7] ),
    .A2(_1358_));
 sg13g2_xnor2_1 _5233_ (.Y(_1373_),
    .A(_3161_),
    .B(_1356_));
 sg13g2_a21oi_1 _5234_ (.A1(_1372_),
    .A2(_1373_),
    .Y(_1374_),
    .B1(_1357_));
 sg13g2_mux2_1 _5235_ (.A0(_0077_),
    .A1(_0052_),
    .S(net851),
    .X(_1375_));
 sg13g2_xnor2_1 _5236_ (.Y(_1376_),
    .A(_3162_),
    .B(_1375_));
 sg13g2_nand2b_1 _5237_ (.Y(_1377_),
    .B(_1376_),
    .A_N(_1374_));
 sg13g2_xor2_1 _5238_ (.B(_1376_),
    .A(_1374_),
    .X(_1378_));
 sg13g2_inv_1 _5239_ (.Y(_1379_),
    .A(_1378_));
 sg13g2_xor2_1 _5240_ (.B(_1373_),
    .A(_1372_),
    .X(_1380_));
 sg13g2_nand2b_1 _5241_ (.Y(_1381_),
    .B(net966),
    .A_N(net969));
 sg13g2_nor4_1 _5242_ (.A(net963),
    .B(net940),
    .C(net972),
    .D(_1381_),
    .Y(_1382_));
 sg13g2_nand2_1 _5243_ (.Y(_1383_),
    .A(net974),
    .B(_1219_));
 sg13g2_a221oi_1 _5244_ (.B2(_1383_),
    .C1(_1220_),
    .B1(_1382_),
    .A1(_3131_),
    .Y(_1384_),
    .A2(_0080_));
 sg13g2_and4_1 _5245_ (.A(net974),
    .B(_1062_),
    .C(_1218_),
    .D(_1382_),
    .X(_1385_));
 sg13g2_nor3_2 _5246_ (.A(_1058_),
    .B(_1384_),
    .C(_1385_),
    .Y(_1386_));
 sg13g2_nor2_1 _5247_ (.A(\vgademo.a_scrolly[10] ),
    .B(_1053_),
    .Y(_1387_));
 sg13g2_nand2_1 _5248_ (.Y(_1388_),
    .A(\vgademo.a_scrolly[13] ),
    .B(net961));
 sg13g2_o21ai_1 _5249_ (.B1(_1089_),
    .Y(_1389_),
    .A1(_1387_),
    .A2(_1388_));
 sg13g2_a21oi_2 _5250_ (.B1(_1386_),
    .Y(_1390_),
    .A2(_1389_),
    .A1(_1088_));
 sg13g2_a21o_2 _5251_ (.A2(_1389_),
    .A1(_1088_),
    .B1(_1386_),
    .X(_1391_));
 sg13g2_nor2_1 _5252_ (.A(_1083_),
    .B(_1381_),
    .Y(_1392_));
 sg13g2_nor2_1 _5253_ (.A(net974),
    .B(_1059_),
    .Y(_1393_));
 sg13g2_nor3_1 _5254_ (.A(_3134_),
    .B(_1083_),
    .C(_1381_),
    .Y(_1394_));
 sg13g2_nand2_1 _5255_ (.Y(_1395_),
    .A(_1128_),
    .B(_1392_));
 sg13g2_a221oi_1 _5256_ (.B2(_1085_),
    .C1(_1058_),
    .B1(_1395_),
    .A1(_1393_),
    .Y(_1396_),
    .A2(_1394_));
 sg13g2_and3_1 _5257_ (.X(_1397_),
    .A(_0075_),
    .B(_1059_),
    .C(_1115_));
 sg13g2_a21oi_1 _5258_ (.A1(net970),
    .A2(_1049_),
    .Y(_1398_),
    .B1(_1069_));
 sg13g2_nor2b_1 _5259_ (.A(_1398_),
    .B_N(_1397_),
    .Y(_1399_));
 sg13g2_xnor2_1 _5260_ (.Y(_1400_),
    .A(_1397_),
    .B(_1398_));
 sg13g2_a221oi_1 _5261_ (.B2(_1389_),
    .C1(_1391_),
    .B1(_1400_),
    .A1(_1236_),
    .Y(_1401_),
    .A2(net903));
 sg13g2_nor2_1 _5262_ (.A(net985),
    .B(_3247_),
    .Y(_1402_));
 sg13g2_nor3_1 _5263_ (.A(net985),
    .B(\vgademo.h_count[4] ),
    .C(_3247_),
    .Y(_1403_));
 sg13g2_nor2_1 _5264_ (.A(net941),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_nand2_1 _5265_ (.Y(_1405_),
    .A(net984),
    .B(_1404_));
 sg13g2_inv_1 _5266_ (.Y(_1406_),
    .A(_1405_));
 sg13g2_nand2_1 _5267_ (.Y(_1407_),
    .A(_0037_),
    .B(_1405_));
 sg13g2_xor2_1 _5268_ (.B(_1407_),
    .A(_0038_),
    .X(_1408_));
 sg13g2_nand2_1 _5269_ (.Y(_1409_),
    .A(_0031_),
    .B(net849));
 sg13g2_o21ai_1 _5270_ (.B1(_1409_),
    .Y(_1410_),
    .A1(net850),
    .A2(_1408_));
 sg13g2_nor2b_1 _5271_ (.A(_1410_),
    .B_N(_1401_),
    .Y(_1411_));
 sg13g2_xnor2_1 _5272_ (.Y(_1412_),
    .A(_1401_),
    .B(_1410_));
 sg13g2_inv_1 _5273_ (.Y(_1413_),
    .A(_1412_));
 sg13g2_nand2_1 _5274_ (.Y(_1414_),
    .A(_1048_),
    .B(_1222_));
 sg13g2_xor2_1 _5275_ (.B(_1383_),
    .A(_0075_),
    .X(_1415_));
 sg13g2_a221oi_1 _5276_ (.B2(_1389_),
    .C1(_1391_),
    .B1(_1415_),
    .A1(net903),
    .Y(_1416_),
    .A2(_1414_));
 sg13g2_xnor2_1 _5277_ (.Y(_1417_),
    .A(_3125_),
    .B(_1405_));
 sg13g2_nor2_1 _5278_ (.A(net849),
    .B(_1417_),
    .Y(_1418_));
 sg13g2_a21oi_2 _5279_ (.B1(_1418_),
    .Y(_1419_),
    .A2(net849),
    .A1(_0046_));
 sg13g2_and2_1 _5280_ (.A(_1416_),
    .B(_1419_),
    .X(_1420_));
 sg13g2_nand2_1 _5281_ (.Y(_1421_),
    .A(_1416_),
    .B(_1419_));
 sg13g2_xnor2_1 _5282_ (.Y(_1422_),
    .A(_3135_),
    .B(_1218_));
 sg13g2_a221oi_1 _5283_ (.B2(_1389_),
    .C1(_1391_),
    .B1(_1422_),
    .A1(net975),
    .Y(_1423_),
    .A2(net903));
 sg13g2_xnor2_1 _5284_ (.Y(_1424_),
    .A(_0036_),
    .B(_1404_));
 sg13g2_nand2_1 _5285_ (.Y(_1425_),
    .A(_0030_),
    .B(net849));
 sg13g2_o21ai_1 _5286_ (.B1(_1425_),
    .Y(_1426_),
    .A1(_1355_),
    .A2(_1424_));
 sg13g2_nor2b_1 _5287_ (.A(_1426_),
    .B_N(_1423_),
    .Y(_1427_));
 sg13g2_nand2b_1 _5288_ (.Y(_1428_),
    .B(_1423_),
    .A_N(_1426_));
 sg13g2_nor2b_1 _5289_ (.A(_1088_),
    .B_N(_1389_),
    .Y(_1429_));
 sg13g2_a22oi_1 _5290_ (.Y(_1430_),
    .B1(_1429_),
    .B2(_1230_),
    .A2(_1396_),
    .A1(_3139_));
 sg13g2_or2_1 _5291_ (.X(_1431_),
    .B(_1430_),
    .A(_1386_));
 sg13g2_xnor2_1 _5292_ (.Y(_1432_),
    .A(net941),
    .B(_1403_));
 sg13g2_mux2_1 _5293_ (.A0(_0047_),
    .A1(_1432_),
    .S(_1354_),
    .X(_1433_));
 sg13g2_or2_2 _5294_ (.X(_1434_),
    .B(_1433_),
    .A(_1431_));
 sg13g2_a221oi_1 _5295_ (.B2(_0064_),
    .C1(_1391_),
    .B1(net903),
    .A1(net981),
    .Y(_1435_),
    .A2(_1389_));
 sg13g2_inv_1 _5296_ (.Y(_1436_),
    .A(_1435_));
 sg13g2_xor2_1 _5297_ (.B(_1402_),
    .A(_0044_),
    .X(_1437_));
 sg13g2_o21ai_1 _5298_ (.B1(_0029_),
    .Y(_1438_),
    .A1(_1349_),
    .A2(_1352_));
 sg13g2_nand3_1 _5299_ (.B(net854),
    .C(_1437_),
    .A(net856),
    .Y(_1439_));
 sg13g2_and3_1 _5300_ (.X(_1440_),
    .A(_1435_),
    .B(_1438_),
    .C(_1439_));
 sg13g2_nand4_1 _5301_ (.B(_3247_),
    .C(net856),
    .A(_3222_),
    .Y(_1441_),
    .D(net854));
 sg13g2_o21ai_1 _5302_ (.B1(_0028_),
    .Y(_1442_),
    .A1(_1349_),
    .A2(_1352_));
 sg13g2_nand3_1 _5303_ (.B(_1441_),
    .C(_1442_),
    .A(_1390_),
    .Y(_1443_));
 sg13g2_xnor2_1 _5304_ (.Y(_1444_),
    .A(_0034_),
    .B(_3247_));
 sg13g2_nand3_1 _5305_ (.B(net854),
    .C(_1444_),
    .A(net856),
    .Y(_1445_));
 sg13g2_o21ai_1 _5306_ (.B1(_0048_),
    .Y(_1446_),
    .A1(_1349_),
    .A2(_1352_));
 sg13g2_nand2_1 _5307_ (.Y(_1447_),
    .A(_1445_),
    .B(_1446_));
 sg13g2_nand3_1 _5308_ (.B(_1445_),
    .C(_1446_),
    .A(_1390_),
    .Y(_1448_));
 sg13g2_nand3_1 _5309_ (.B(_1438_),
    .C(_1439_),
    .A(_1436_),
    .Y(_1449_));
 sg13g2_a21o_1 _5310_ (.A2(_1439_),
    .A1(_1438_),
    .B1(_1436_),
    .X(_1450_));
 sg13g2_a22oi_1 _5311_ (.Y(_1451_),
    .B1(_1449_),
    .B2(_1450_),
    .A2(_1448_),
    .A1(_1443_));
 sg13g2_xor2_1 _5312_ (.B(_1433_),
    .A(_1431_),
    .X(_1452_));
 sg13g2_o21ai_1 _5313_ (.B1(_1452_),
    .Y(_1453_),
    .A1(_1440_),
    .A2(_1451_));
 sg13g2_xnor2_1 _5314_ (.Y(_1454_),
    .A(_1423_),
    .B(_1426_));
 sg13g2_xor2_1 _5315_ (.B(_1426_),
    .A(_1423_),
    .X(_1455_));
 sg13g2_a21oi_2 _5316_ (.B1(_1455_),
    .Y(_1456_),
    .A2(net836),
    .A1(_1434_));
 sg13g2_a21o_2 _5317_ (.A2(net836),
    .A1(_1434_),
    .B1(_1455_),
    .X(_1457_));
 sg13g2_xor2_1 _5318_ (.B(_1419_),
    .A(_1416_),
    .X(_1458_));
 sg13g2_xnor2_1 _5319_ (.Y(_1459_),
    .A(_1416_),
    .B(_1419_));
 sg13g2_a21oi_2 _5320_ (.B1(_1459_),
    .Y(_1460_),
    .A2(_1457_),
    .A1(_1428_));
 sg13g2_o21ai_1 _5321_ (.B1(_1458_),
    .Y(_1461_),
    .A1(_1427_),
    .A2(_1456_));
 sg13g2_a21oi_2 _5322_ (.B1(_1413_),
    .Y(_1462_),
    .A2(net830),
    .A1(_1421_));
 sg13g2_o21ai_1 _5323_ (.B1(_1412_),
    .Y(_1463_),
    .A1(_1420_),
    .A2(_1460_));
 sg13g2_xor2_1 _5324_ (.B(_1050_),
    .A(_0080_),
    .X(_1464_));
 sg13g2_nand2_1 _5325_ (.Y(_1465_),
    .A(_1399_),
    .B(_1464_));
 sg13g2_or2_1 _5326_ (.X(_1466_),
    .B(_1464_),
    .A(_1399_));
 sg13g2_nand3_1 _5327_ (.B(_1465_),
    .C(_1466_),
    .A(_1429_),
    .Y(_1467_));
 sg13g2_nand3_1 _5328_ (.B(_1048_),
    .C(_1222_),
    .A(_0078_),
    .Y(_1468_));
 sg13g2_or2_1 _5329_ (.X(_1469_),
    .B(_1468_),
    .A(_3133_));
 sg13g2_o21ai_1 _5330_ (.B1(net967),
    .Y(_1470_),
    .A1(net968),
    .A2(_1048_));
 sg13g2_nand2_1 _5331_ (.Y(_1471_),
    .A(_1047_),
    .B(_1075_));
 sg13g2_nand3_1 _5332_ (.B(_1470_),
    .C(_1471_),
    .A(_1468_),
    .Y(_1472_));
 sg13g2_nand3_1 _5333_ (.B(_1469_),
    .C(_1472_),
    .A(net903),
    .Y(_1473_));
 sg13g2_a21o_2 _5334_ (.A2(_1473_),
    .A1(_1467_),
    .B1(_1386_),
    .X(_1474_));
 sg13g2_nand2_1 _5335_ (.Y(_1475_),
    .A(_0045_),
    .B(net849));
 sg13g2_nor3_2 _5336_ (.A(\vgademo.h_count[7] ),
    .B(net983),
    .C(_1406_),
    .Y(_1476_));
 sg13g2_nor2_1 _5337_ (.A(_3126_),
    .B(_1476_),
    .Y(_1477_));
 sg13g2_xnor2_1 _5338_ (.Y(_1478_),
    .A(\vgademo.h_count[9] ),
    .B(_1476_));
 sg13g2_o21ai_1 _5339_ (.B1(_1475_),
    .Y(_1479_),
    .A1(net850),
    .A2(_1478_));
 sg13g2_nor2_1 _5340_ (.A(_1474_),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_xor2_1 _5341_ (.B(_1479_),
    .A(_1474_),
    .X(_1481_));
 sg13g2_o21ai_1 _5342_ (.B1(_1481_),
    .Y(_1482_),
    .A1(_1411_),
    .A2(_1462_));
 sg13g2_or3_2 _5343_ (.A(_1411_),
    .B(_1462_),
    .C(_1481_),
    .X(_1483_));
 sg13g2_and2_1 _5344_ (.A(_1482_),
    .B(_1483_),
    .X(_1484_));
 sg13g2_nand2_2 _5345_ (.Y(_1485_),
    .A(_1482_),
    .B(_1483_));
 sg13g2_nor3_2 _5346_ (.A(_1412_),
    .B(_1420_),
    .C(_1460_),
    .Y(_1486_));
 sg13g2_nand3_1 _5347_ (.B(_1421_),
    .C(net830),
    .A(_1413_),
    .Y(_1487_));
 sg13g2_nor2_1 _5348_ (.A(_1462_),
    .B(_1486_),
    .Y(_1488_));
 sg13g2_nand2_2 _5349_ (.Y(_1489_),
    .A(net825),
    .B(net824));
 sg13g2_and3_1 _5350_ (.X(_1490_),
    .A(_1434_),
    .B(net836),
    .C(_1455_));
 sg13g2_nand3_1 _5351_ (.B(net836),
    .C(_1455_),
    .A(_1434_),
    .Y(_1491_));
 sg13g2_nand3_1 _5352_ (.B(net836),
    .C(_1454_),
    .A(_1434_),
    .Y(_1492_));
 sg13g2_a21o_1 _5353_ (.A2(net836),
    .A1(_1434_),
    .B1(_1454_),
    .X(_1493_));
 sg13g2_nor2_2 _5354_ (.A(_1456_),
    .B(_1490_),
    .Y(_1494_));
 sg13g2_nand2_2 _5355_ (.Y(_1495_),
    .A(_1457_),
    .B(_1491_));
 sg13g2_or3_2 _5356_ (.A(_1440_),
    .B(_1451_),
    .C(_1452_),
    .X(_1496_));
 sg13g2_and2_2 _5357_ (.A(net837),
    .B(_1496_),
    .X(_1497_));
 sg13g2_nand2_2 _5358_ (.Y(_1498_),
    .A(net837),
    .B(_1496_));
 sg13g2_a21oi_1 _5359_ (.A1(_1441_),
    .A2(_1442_),
    .Y(_1499_),
    .B1(_1391_));
 sg13g2_xor2_1 _5360_ (.B(_1499_),
    .A(_1447_),
    .X(_1500_));
 sg13g2_and4_2 _5361_ (.A(_1443_),
    .B(_1448_),
    .C(_1449_),
    .D(_1450_),
    .X(_1501_));
 sg13g2_nor2_2 _5362_ (.A(_1451_),
    .B(_1501_),
    .Y(_1502_));
 sg13g2_nor3_2 _5363_ (.A(_1451_),
    .B(_1500_),
    .C(_1501_),
    .Y(_1503_));
 sg13g2_and2_1 _5364_ (.A(_1497_),
    .B(_1502_),
    .X(_1504_));
 sg13g2_nand3_1 _5365_ (.B(_1496_),
    .C(_1502_),
    .A(net837),
    .Y(_1505_));
 sg13g2_nor2_1 _5366_ (.A(_1500_),
    .B(_1505_),
    .Y(_1506_));
 sg13g2_nand3_1 _5367_ (.B(_1496_),
    .C(_1503_),
    .A(net836),
    .Y(_1507_));
 sg13g2_a21o_1 _5368_ (.A2(_1496_),
    .A1(net836),
    .B1(_1503_),
    .X(_1508_));
 sg13g2_and2_1 _5369_ (.A(_1507_),
    .B(_1508_),
    .X(_1509_));
 sg13g2_a22oi_1 _5370_ (.Y(_1510_),
    .B1(_1507_),
    .B2(_1508_),
    .A2(_1493_),
    .A1(_1492_));
 sg13g2_nor3_2 _5371_ (.A(_1427_),
    .B(_1456_),
    .C(_1458_),
    .Y(_1511_));
 sg13g2_nand3_1 _5372_ (.B(_1457_),
    .C(_1459_),
    .A(_1428_),
    .Y(_1512_));
 sg13g2_nor2_2 _5373_ (.A(net831),
    .B(_1511_),
    .Y(_1513_));
 sg13g2_nand2_2 _5374_ (.Y(_1514_),
    .A(net830),
    .B(_1512_));
 sg13g2_a21oi_1 _5375_ (.A1(_1457_),
    .A2(_1491_),
    .Y(_1515_),
    .B1(_1497_));
 sg13g2_or3_1 _5376_ (.A(net831),
    .B(_1511_),
    .C(_1515_),
    .X(_1516_));
 sg13g2_nor4_2 _5377_ (.A(net831),
    .B(_1510_),
    .C(_1511_),
    .Y(_1517_),
    .D(_1515_));
 sg13g2_and3_1 _5378_ (.X(_1518_),
    .A(_1457_),
    .B(_1491_),
    .C(_1508_));
 sg13g2_a21oi_2 _5379_ (.B1(_1518_),
    .Y(_1519_),
    .A2(net828),
    .A1(net829));
 sg13g2_or4_1 _5380_ (.A(_1462_),
    .B(_1486_),
    .C(_1517_),
    .D(_1519_),
    .X(_1520_));
 sg13g2_nand2_1 _5381_ (.Y(_1521_),
    .A(_1494_),
    .B(_1504_));
 sg13g2_nor3_2 _5382_ (.A(net831),
    .B(_1495_),
    .C(_1511_),
    .Y(_1522_));
 sg13g2_nand3_1 _5383_ (.B(_1494_),
    .C(_1512_),
    .A(net829),
    .Y(_1523_));
 sg13g2_nor2_1 _5384_ (.A(_1505_),
    .B(_1523_),
    .Y(_1524_));
 sg13g2_nand4_1 _5385_ (.B(_1494_),
    .C(_1504_),
    .A(net829),
    .Y(_1525_),
    .D(net828));
 sg13g2_a21oi_1 _5386_ (.A1(net825),
    .A2(_1487_),
    .Y(_1526_),
    .B1(_1525_));
 sg13g2_nor3_1 _5387_ (.A(_1456_),
    .B(_1490_),
    .C(_1507_),
    .Y(_1527_));
 sg13g2_nand3_1 _5388_ (.B(net828),
    .C(_1527_),
    .A(net830),
    .Y(_1528_));
 sg13g2_a21o_1 _5389_ (.A2(net824),
    .A1(_1463_),
    .B1(_1528_),
    .X(_1529_));
 sg13g2_and2_1 _5390_ (.A(_1520_),
    .B(_1529_),
    .X(_1530_));
 sg13g2_a221oi_1 _5391_ (.B2(_1509_),
    .C1(_1514_),
    .B1(_1494_),
    .A1(net825),
    .Y(_1531_),
    .A2(net824));
 sg13g2_xnor2_1 _5392_ (.Y(_1532_),
    .A(_1359_),
    .B(_1369_));
 sg13g2_xor2_1 _5393_ (.B(_1369_),
    .A(_1359_),
    .X(_1533_));
 sg13g2_a21oi_1 _5394_ (.A1(_1495_),
    .A2(_1505_),
    .Y(_1534_),
    .B1(net834));
 sg13g2_nand2_1 _5395_ (.Y(_1535_),
    .A(_1531_),
    .B(_1534_));
 sg13g2_o21ai_1 _5396_ (.B1(_1500_),
    .Y(_1536_),
    .A1(_1451_),
    .A2(_1501_));
 sg13g2_a21o_1 _5397_ (.A2(_1496_),
    .A1(net837),
    .B1(_1502_),
    .X(_1537_));
 sg13g2_nor2_1 _5398_ (.A(_1497_),
    .B(_1536_),
    .Y(_1538_));
 sg13g2_a221oi_1 _5399_ (.B2(net837),
    .C1(_1536_),
    .B1(_1496_),
    .A1(_1457_),
    .Y(_1539_),
    .A2(_1491_));
 sg13g2_a221oi_1 _5400_ (.B2(net829),
    .C1(_1494_),
    .B1(net828),
    .A1(net837),
    .Y(_1540_),
    .A2(_1496_));
 sg13g2_o21ai_1 _5401_ (.B1(_1539_),
    .Y(_1541_),
    .A1(net831),
    .A2(_1511_));
 sg13g2_and2_1 _5402_ (.A(_1505_),
    .B(_1537_),
    .X(_1542_));
 sg13g2_nor2_1 _5403_ (.A(_1516_),
    .B(_1542_),
    .Y(_1543_));
 sg13g2_o21ai_1 _5404_ (.B1(_1541_),
    .Y(_1544_),
    .A1(_1516_),
    .A2(_1542_));
 sg13g2_a22oi_1 _5405_ (.Y(_1545_),
    .B1(_1544_),
    .B2(net819),
    .A2(_1534_),
    .A1(_1531_));
 sg13g2_mux2_1 _5406_ (.A0(_1530_),
    .A1(_1545_),
    .S(net817),
    .X(_1546_));
 sg13g2_o21ai_1 _5407_ (.B1(_1507_),
    .Y(_1547_),
    .A1(_1456_),
    .A2(_1490_));
 sg13g2_a21o_1 _5408_ (.A2(net828),
    .A1(net829),
    .B1(_1547_),
    .X(_1548_));
 sg13g2_nor2b_1 _5409_ (.A(_1543_),
    .B_N(_1548_),
    .Y(_1549_));
 sg13g2_nor3_2 _5410_ (.A(_1485_),
    .B(_1489_),
    .C(_1549_),
    .Y(_1550_));
 sg13g2_a21o_1 _5411_ (.A2(_1513_),
    .A1(_1509_),
    .B1(net819),
    .X(_1551_));
 sg13g2_a221oi_1 _5412_ (.B2(net817),
    .C1(net834),
    .B1(_1551_),
    .A1(net819),
    .Y(_1552_),
    .A2(_1517_));
 sg13g2_nand2_1 _5413_ (.Y(_1553_),
    .A(_1497_),
    .B(_1536_));
 sg13g2_a22oi_1 _5414_ (.Y(_1554_),
    .B1(_1497_),
    .B2(_1536_),
    .A2(_1491_),
    .A1(_1457_));
 sg13g2_nand2_1 _5415_ (.Y(_1555_),
    .A(_1495_),
    .B(_1553_));
 sg13g2_or3_2 _5416_ (.A(net831),
    .B(_1511_),
    .C(_1554_),
    .X(_1556_));
 sg13g2_nand2_1 _5417_ (.Y(_1557_),
    .A(_1494_),
    .B(_1537_));
 sg13g2_nand2_1 _5418_ (.Y(_1558_),
    .A(_1514_),
    .B(_1557_));
 sg13g2_a21o_1 _5419_ (.A2(_1558_),
    .A1(_1556_),
    .B1(net819),
    .X(_1559_));
 sg13g2_nand4_1 _5420_ (.B(net824),
    .C(_1510_),
    .A(_1463_),
    .Y(_1560_),
    .D(_1513_));
 sg13g2_a21oi_1 _5421_ (.A1(_1559_),
    .A2(_1560_),
    .Y(_1561_),
    .B1(net817));
 sg13g2_a221oi_1 _5422_ (.B2(_1560_),
    .C1(net832),
    .B1(_1559_),
    .A1(_1482_),
    .Y(_1562_),
    .A2(_1483_));
 sg13g2_or3_1 _5423_ (.A(_1550_),
    .B(_1552_),
    .C(_1562_),
    .X(_1563_));
 sg13g2_nand4_1 _5424_ (.B(_1531_),
    .C(net835),
    .A(net817),
    .Y(_1564_),
    .D(_1547_));
 sg13g2_o21ai_1 _5425_ (.B1(_1564_),
    .Y(_1565_),
    .A1(net826),
    .A2(_1546_));
 sg13g2_a21o_1 _5426_ (.A2(_1563_),
    .A1(net826),
    .B1(_1565_),
    .X(_1566_));
 sg13g2_o21ai_1 _5427_ (.B1(_1377_),
    .Y(_1567_),
    .A1(\vgademo.b_cos[9] ),
    .A2(_1375_));
 sg13g2_nand2_1 _5428_ (.Y(_1568_),
    .A(_0053_),
    .B(net851));
 sg13g2_o21ai_1 _5429_ (.B1(_1568_),
    .Y(_1569_),
    .A1(_3128_),
    .A2(net851));
 sg13g2_xnor2_1 _5430_ (.Y(_1570_),
    .A(_3163_),
    .B(_1569_));
 sg13g2_nand2b_1 _5431_ (.Y(_1571_),
    .B(_1567_),
    .A_N(_1570_));
 sg13g2_xnor2_1 _5432_ (.Y(_1572_),
    .A(_1567_),
    .B(_1570_));
 sg13g2_xor2_1 _5433_ (.B(_1570_),
    .A(_1567_),
    .X(_1573_));
 sg13g2_nor3_1 _5434_ (.A(_1495_),
    .B(_1504_),
    .C(_1538_),
    .Y(_1574_));
 sg13g2_nand2_1 _5435_ (.Y(_1575_),
    .A(_1513_),
    .B(_1574_));
 sg13g2_and4_1 _5436_ (.A(_1482_),
    .B(_1483_),
    .C(net819),
    .D(_1575_),
    .X(_1576_));
 sg13g2_nand2_1 _5437_ (.Y(_1577_),
    .A(_1519_),
    .B(_1547_));
 sg13g2_a21oi_1 _5438_ (.A1(net825),
    .A2(_1487_),
    .Y(_1578_),
    .B1(_1540_));
 sg13g2_a221oi_1 _5439_ (.B2(_1522_),
    .C1(_1540_),
    .B1(_1509_),
    .A1(net825),
    .Y(_1579_),
    .A2(net824));
 sg13g2_inv_1 _5440_ (.Y(_1580_),
    .A(_1579_));
 sg13g2_a21oi_1 _5441_ (.A1(_1509_),
    .A2(_1522_),
    .Y(_1581_),
    .B1(_1540_));
 sg13g2_nand2_1 _5442_ (.Y(_1582_),
    .A(net821),
    .B(_1581_));
 sg13g2_a21o_1 _5443_ (.A2(_1582_),
    .A1(_1559_),
    .B1(net817),
    .X(_1583_));
 sg13g2_a22oi_1 _5444_ (.Y(_1584_),
    .B1(_1579_),
    .B2(net817),
    .A2(_1577_),
    .A1(_1576_));
 sg13g2_a21o_1 _5445_ (.A2(_1584_),
    .A1(_1583_),
    .B1(net835),
    .X(_1585_));
 sg13g2_and2_1 _5446_ (.A(_1494_),
    .B(_1542_),
    .X(_1586_));
 sg13g2_nand2_1 _5447_ (.Y(_1587_),
    .A(_1514_),
    .B(_1586_));
 sg13g2_nor2b_1 _5448_ (.A(_1538_),
    .B_N(_1554_),
    .Y(_1588_));
 sg13g2_a22oi_1 _5449_ (.Y(_1589_),
    .B1(_1513_),
    .B2(_1588_),
    .A2(net824),
    .A1(net825));
 sg13g2_a22oi_1 _5450_ (.Y(_1590_),
    .B1(_1587_),
    .B2(_1589_),
    .A2(_1581_),
    .A1(net819));
 sg13g2_nor2_1 _5451_ (.A(_1484_),
    .B(_1590_),
    .Y(_1591_));
 sg13g2_nand2_1 _5452_ (.Y(_1592_),
    .A(_1522_),
    .B(_1537_));
 sg13g2_o21ai_1 _5453_ (.B1(_1578_),
    .Y(_1593_),
    .A1(_1506_),
    .A2(_1592_));
 sg13g2_o21ai_1 _5454_ (.B1(_1548_),
    .Y(_1594_),
    .A1(_1556_),
    .A2(_1586_));
 sg13g2_nand2_1 _5455_ (.Y(_1595_),
    .A(net820),
    .B(_1594_));
 sg13g2_a21oi_1 _5456_ (.A1(_1593_),
    .A2(_1595_),
    .Y(_1596_),
    .B1(_1485_));
 sg13g2_o21ai_1 _5457_ (.B1(net835),
    .Y(_1597_),
    .A1(_1591_),
    .A2(_1596_));
 sg13g2_nand3_1 _5458_ (.B(_1585_),
    .C(_1597_),
    .A(net826),
    .Y(_1598_));
 sg13g2_nand2_1 _5459_ (.Y(_1599_),
    .A(_1522_),
    .B(_1553_));
 sg13g2_nand4_1 _5460_ (.B(net834),
    .C(_1577_),
    .A(net821),
    .Y(_1600_),
    .D(_1599_));
 sg13g2_o21ai_1 _5461_ (.B1(_1548_),
    .Y(_1601_),
    .A1(_1556_),
    .A2(_1574_));
 sg13g2_nand3_1 _5462_ (.B(net832),
    .C(_1601_),
    .A(net819),
    .Y(_1602_));
 sg13g2_nand3_1 _5463_ (.B(_1600_),
    .C(_1602_),
    .A(_1535_),
    .Y(_1603_));
 sg13g2_nor2_1 _5464_ (.A(net826),
    .B(_1561_),
    .Y(_1604_));
 sg13g2_and3_1 _5465_ (.X(_1605_),
    .A(_1531_),
    .B(net835),
    .C(_1555_));
 sg13g2_o21ai_1 _5466_ (.B1(net818),
    .Y(_1606_),
    .A1(_1603_),
    .A2(_1605_));
 sg13g2_a21oi_1 _5467_ (.A1(_1604_),
    .A2(_1606_),
    .Y(_1607_),
    .B1(_1378_));
 sg13g2_a221oi_1 _5468_ (.B2(_1607_),
    .C1(_1573_),
    .B1(_1598_),
    .A1(_1378_),
    .Y(_1608_),
    .A2(_1566_));
 sg13g2_o21ai_1 _5469_ (.B1(_1541_),
    .Y(_1609_),
    .A1(_1556_),
    .A2(_1586_));
 sg13g2_a22oi_1 _5470_ (.Y(_1610_),
    .B1(_1609_),
    .B2(net821),
    .A2(_1555_),
    .A1(_1531_));
 sg13g2_nand2_1 _5471_ (.Y(_1611_),
    .A(_1514_),
    .B(_1588_));
 sg13g2_and2_1 _5472_ (.A(_1576_),
    .B(_1611_),
    .X(_1612_));
 sg13g2_o21ai_1 _5473_ (.B1(_1580_),
    .Y(_1613_),
    .A1(net818),
    .A2(_1520_));
 sg13g2_nand3b_1 _5474_ (.B(net834),
    .C(net818),
    .Y(_1614_),
    .A_N(_1610_));
 sg13g2_or3_1 _5475_ (.A(net817),
    .B(_1530_),
    .C(net833),
    .X(_1615_));
 sg13g2_o21ai_1 _5476_ (.B1(net833),
    .Y(_1616_),
    .A1(_1612_),
    .A2(_1613_));
 sg13g2_nand4_1 _5477_ (.B(_1614_),
    .C(_1615_),
    .A(net827),
    .Y(_1617_),
    .D(_1616_));
 sg13g2_a21oi_1 _5478_ (.A1(net835),
    .A2(_1593_),
    .Y(_1618_),
    .B1(_1485_));
 sg13g2_and3_1 _5479_ (.X(_1619_),
    .A(net829),
    .B(net828),
    .C(_1547_));
 sg13g2_a21oi_1 _5480_ (.A1(_1514_),
    .A2(_1588_),
    .Y(_1620_),
    .B1(_1619_));
 sg13g2_o21ai_1 _5481_ (.B1(net820),
    .Y(_1621_),
    .A1(_1524_),
    .A2(_1620_));
 sg13g2_nand2b_1 _5482_ (.Y(_1622_),
    .B(_1522_),
    .A_N(_1538_));
 sg13g2_o21ai_1 _5483_ (.B1(_1578_),
    .Y(_1623_),
    .A1(_1506_),
    .A2(_1622_));
 sg13g2_nand3_1 _5484_ (.B(_1621_),
    .C(_1623_),
    .A(net832),
    .Y(_1624_));
 sg13g2_o21ai_1 _5485_ (.B1(_1624_),
    .Y(_1625_),
    .A1(_1612_),
    .A2(_1618_));
 sg13g2_nor2_1 _5486_ (.A(_1498_),
    .B(_1503_),
    .Y(_1626_));
 sg13g2_a221oi_1 _5487_ (.B2(_1495_),
    .C1(_1518_),
    .B1(_1626_),
    .A1(net829),
    .Y(_1627_),
    .A2(net828));
 sg13g2_nor4_2 _5488_ (.A(_1462_),
    .B(_1486_),
    .C(_1517_),
    .Y(_1628_),
    .D(_1627_));
 sg13g2_nor2_1 _5489_ (.A(_1579_),
    .B(_1628_),
    .Y(_1629_));
 sg13g2_nor2_1 _5490_ (.A(net818),
    .B(_1629_),
    .Y(_1630_));
 sg13g2_nor2_1 _5491_ (.A(net826),
    .B(_1630_),
    .Y(_1631_));
 sg13g2_a21oi_1 _5492_ (.A1(_1625_),
    .A2(_1631_),
    .Y(_1632_),
    .B1(_1378_));
 sg13g2_nand3b_1 _5493_ (.B(net819),
    .C(_1516_),
    .Y(_1633_),
    .A_N(_1519_));
 sg13g2_a21oi_1 _5494_ (.A1(_1528_),
    .A2(_1633_),
    .Y(_1634_),
    .B1(net817));
 sg13g2_inv_1 _5495_ (.Y(_1635_),
    .A(_1634_));
 sg13g2_nand3_1 _5496_ (.B(net828),
    .C(_1518_),
    .A(net829),
    .Y(_1636_));
 sg13g2_a21oi_1 _5497_ (.A1(net825),
    .A2(net824),
    .Y(_1637_),
    .B1(_1636_));
 sg13g2_o21ai_1 _5498_ (.B1(_1541_),
    .Y(_1638_),
    .A1(_1514_),
    .A2(_1557_));
 sg13g2_a21oi_1 _5499_ (.A1(net820),
    .A2(_1638_),
    .Y(_1639_),
    .B1(_1637_));
 sg13g2_nor2_1 _5500_ (.A(net834),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_or4_2 _5501_ (.A(net831),
    .B(_1495_),
    .C(_1511_),
    .D(_1553_),
    .X(_1641_));
 sg13g2_or2_1 _5502_ (.X(_1642_),
    .B(_1641_),
    .A(net832));
 sg13g2_o21ai_1 _5503_ (.B1(_1541_),
    .Y(_1643_),
    .A1(_1498_),
    .A2(_1523_));
 sg13g2_nand3_1 _5504_ (.B(net834),
    .C(_1643_),
    .A(net820),
    .Y(_1644_));
 sg13g2_o21ai_1 _5505_ (.B1(_1644_),
    .Y(_1645_),
    .A1(net820),
    .A2(_1642_));
 sg13g2_nor3_1 _5506_ (.A(net826),
    .B(_1640_),
    .C(_1645_),
    .Y(_1646_));
 sg13g2_a21oi_1 _5507_ (.A1(_1541_),
    .A2(_1641_),
    .Y(_1647_),
    .B1(_1489_));
 sg13g2_nand2b_1 _5508_ (.Y(_1648_),
    .B(net826),
    .A_N(_1526_));
 sg13g2_o21ai_1 _5509_ (.B1(net818),
    .Y(_1649_),
    .A1(_1647_),
    .A2(_1648_));
 sg13g2_o21ai_1 _5510_ (.B1(_1635_),
    .Y(_1650_),
    .A1(_1646_),
    .A2(_1649_));
 sg13g2_a221oi_1 _5511_ (.B2(_1378_),
    .C1(_1572_),
    .B1(_1650_),
    .A1(_1617_),
    .Y(_1651_),
    .A2(_1632_));
 sg13g2_o21ai_1 _5512_ (.B1(_1571_),
    .Y(_1652_),
    .A1(_3163_),
    .A2(_1569_));
 sg13g2_nand2b_2 _5513_ (.Y(_1653_),
    .B(net952),
    .A_N(\vgademo.b_cos[11] ));
 sg13g2_xnor2_1 _5514_ (.Y(_1654_),
    .A(net951),
    .B(\vgademo.b_cos[11] ));
 sg13g2_xor2_1 _5515_ (.B(\vgademo.b_cos[11] ),
    .A(net951),
    .X(_1655_));
 sg13g2_mux2_1 _5516_ (.A0(net958),
    .A1(\vgademo.plane_du[8] ),
    .S(net851),
    .X(_1656_));
 sg13g2_xnor2_1 _5517_ (.Y(_1657_),
    .A(_1654_),
    .B(_1656_));
 sg13g2_xnor2_1 _5518_ (.Y(_1658_),
    .A(_1652_),
    .B(_1657_));
 sg13g2_inv_1 _5519_ (.Y(_1659_),
    .A(_1658_));
 sg13g2_nor3_1 _5520_ (.A(_1608_),
    .B(_1651_),
    .C(_1659_),
    .Y(_1660_));
 sg13g2_a21oi_1 _5521_ (.A1(_1463_),
    .A2(net824),
    .Y(_1661_),
    .B1(_1627_));
 sg13g2_nand3_1 _5522_ (.B(_1483_),
    .C(_1661_),
    .A(_1482_),
    .Y(_1662_));
 sg13g2_o21ai_1 _5523_ (.B1(_1662_),
    .Y(_1663_),
    .A1(net818),
    .A2(_1629_));
 sg13g2_o21ai_1 _5524_ (.B1(net834),
    .Y(_1664_),
    .A1(_1612_),
    .A2(_1663_));
 sg13g2_nand3_1 _5525_ (.B(_1514_),
    .C(_1626_),
    .A(_1495_),
    .Y(_1665_));
 sg13g2_nand2b_1 _5526_ (.Y(_1666_),
    .B(_1489_),
    .A_N(_1665_));
 sg13g2_a21oi_1 _5527_ (.A1(net821),
    .A2(_1609_),
    .Y(_1667_),
    .B1(_1637_));
 sg13g2_nand3_1 _5528_ (.B(_1666_),
    .C(_1667_),
    .A(net818),
    .Y(_1668_));
 sg13g2_nor4_1 _5529_ (.A(net831),
    .B(_1511_),
    .C(_1527_),
    .D(_1539_),
    .Y(_1669_));
 sg13g2_a221oi_1 _5530_ (.B2(_1521_),
    .C1(_1669_),
    .B1(_1514_),
    .A1(net825),
    .Y(_1670_),
    .A2(_1487_));
 sg13g2_nor2_1 _5531_ (.A(_1628_),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_a21oi_1 _5532_ (.A1(_1485_),
    .A2(_1671_),
    .Y(_1672_),
    .B1(net835));
 sg13g2_a21oi_1 _5533_ (.A1(_1668_),
    .A2(_1672_),
    .Y(_1673_),
    .B1(net827));
 sg13g2_nand2_1 _5534_ (.Y(_1674_),
    .A(net833),
    .B(_1612_));
 sg13g2_nor2b_1 _5535_ (.A(_1620_),
    .B_N(_1641_),
    .Y(_1675_));
 sg13g2_nor4_1 _5536_ (.A(_1485_),
    .B(_1489_),
    .C(net833),
    .D(_1675_),
    .Y(_1676_));
 sg13g2_nand2_1 _5537_ (.Y(_1677_),
    .A(net826),
    .B(_1662_));
 sg13g2_nor3_1 _5538_ (.A(_1630_),
    .B(_1676_),
    .C(_1677_),
    .Y(_1678_));
 sg13g2_a221oi_1 _5539_ (.B2(_1678_),
    .C1(_1378_),
    .B1(_1674_),
    .A1(_1664_),
    .Y(_1679_),
    .A2(_1673_));
 sg13g2_o21ai_1 _5540_ (.B1(_1560_),
    .Y(_1680_),
    .A1(_1489_),
    .A2(_1665_));
 sg13g2_o21ai_1 _5541_ (.B1(_1485_),
    .Y(_1681_),
    .A1(_1670_),
    .A2(_1680_));
 sg13g2_a21o_1 _5542_ (.A2(_1665_),
    .A1(_1525_),
    .B1(net820),
    .X(_1682_));
 sg13g2_nor3_1 _5543_ (.A(_1485_),
    .B(net832),
    .C(_1682_),
    .Y(_1683_));
 sg13g2_nor3_1 _5544_ (.A(net827),
    .B(_1550_),
    .C(_1683_),
    .Y(_1684_));
 sg13g2_mux2_1 _5545_ (.A0(_1590_),
    .A1(_1623_),
    .S(_1484_),
    .X(_1685_));
 sg13g2_mux2_1 _5546_ (.A0(_1681_),
    .A1(_1685_),
    .S(net832),
    .X(_1686_));
 sg13g2_a21o_1 _5547_ (.A2(_1665_),
    .A1(_1642_),
    .B1(net821),
    .X(_1687_));
 sg13g2_a22oi_1 _5548_ (.Y(_1688_),
    .B1(_1544_),
    .B2(net821),
    .A2(net832),
    .A1(_1526_));
 sg13g2_a21oi_1 _5549_ (.A1(_1687_),
    .A2(_1688_),
    .Y(_1689_),
    .B1(_1485_));
 sg13g2_nor2b_1 _5550_ (.A(_1689_),
    .B_N(net827),
    .Y(_1690_));
 sg13g2_a221oi_1 _5551_ (.B2(_1681_),
    .C1(_1379_),
    .B1(_1690_),
    .A1(_1684_),
    .Y(_1691_),
    .A2(_1686_));
 sg13g2_nor3_1 _5552_ (.A(_1572_),
    .B(_1679_),
    .C(_1691_),
    .Y(_1692_));
 sg13g2_nand2_1 _5553_ (.Y(_1693_),
    .A(net833),
    .B(_1647_));
 sg13g2_a21oi_1 _5554_ (.A1(_1644_),
    .A2(_1693_),
    .Y(_1694_),
    .B1(net827));
 sg13g2_nor2_1 _5555_ (.A(net832),
    .B(_1622_),
    .Y(_1695_));
 sg13g2_o21ai_1 _5556_ (.B1(_1541_),
    .Y(_1696_),
    .A1(net834),
    .A2(_1636_));
 sg13g2_and2_1 _5557_ (.A(net820),
    .B(_1696_),
    .X(_1697_));
 sg13g2_o21ai_1 _5558_ (.B1(net827),
    .Y(_1698_),
    .A1(_1695_),
    .A2(_1697_));
 sg13g2_o21ai_1 _5559_ (.B1(_1698_),
    .Y(_1699_),
    .A1(net820),
    .A2(_1519_));
 sg13g2_o21ai_1 _5560_ (.B1(_1484_),
    .Y(_1700_),
    .A1(_1694_),
    .A2(_1699_));
 sg13g2_nor2_1 _5561_ (.A(_1573_),
    .B(_1634_),
    .Y(_1701_));
 sg13g2_a21o_1 _5562_ (.A2(_1701_),
    .A1(_1700_),
    .B1(_1658_),
    .X(_1702_));
 sg13g2_nor2b_1 _5563_ (.A(_1480_),
    .B_N(_1482_),
    .Y(_1703_));
 sg13g2_xnor2_1 _5564_ (.Y(_1704_),
    .A(net940),
    .B(_1051_));
 sg13g2_nand2_1 _5565_ (.Y(_1705_),
    .A(_1466_),
    .B(_1704_));
 sg13g2_nor2_1 _5566_ (.A(_1054_),
    .B(_1387_),
    .Y(_1706_));
 sg13g2_xnor2_1 _5567_ (.Y(_1707_),
    .A(_1705_),
    .B(_1706_));
 sg13g2_a21oi_1 _5568_ (.A1(_1429_),
    .A2(_1707_),
    .Y(_1708_),
    .B1(net903));
 sg13g2_nand2_1 _5569_ (.Y(_1709_),
    .A(_1470_),
    .B(_1472_));
 sg13g2_a21oi_1 _5570_ (.A1(net965),
    .A2(_1709_),
    .Y(_1710_),
    .B1(net963));
 sg13g2_nor2b_1 _5571_ (.A(_1710_),
    .B_N(net903),
    .Y(_1711_));
 sg13g2_nor3_2 _5572_ (.A(_1386_),
    .B(_1708_),
    .C(_1711_),
    .Y(_1712_));
 sg13g2_nor3_1 _5573_ (.A(\vgademo.h_count[10] ),
    .B(_3126_),
    .C(_1476_),
    .Y(_1713_));
 sg13g2_nor3_1 _5574_ (.A(_3127_),
    .B(net849),
    .C(_1713_),
    .Y(_1714_));
 sg13g2_a21oi_1 _5575_ (.A1(\vgademo.plane_u[21] ),
    .A2(net849),
    .Y(_1715_),
    .B1(_1714_));
 sg13g2_xnor2_1 _5576_ (.Y(_1716_),
    .A(_1712_),
    .B(_1715_));
 sg13g2_xnor2_1 _5577_ (.Y(_1717_),
    .A(net965),
    .B(_1709_));
 sg13g2_xor2_1 _5578_ (.B(_1704_),
    .A(_1466_),
    .X(_1718_));
 sg13g2_a221oi_1 _5579_ (.B2(_1389_),
    .C1(_1391_),
    .B1(_1718_),
    .A1(net903),
    .Y(_1719_),
    .A2(_1717_));
 sg13g2_xnor2_1 _5580_ (.Y(_1720_),
    .A(\vgademo.h_count[10] ),
    .B(_1477_));
 sg13g2_nor2_1 _5581_ (.A(net849),
    .B(_1720_),
    .Y(_1721_));
 sg13g2_a21oi_2 _5582_ (.B1(_1721_),
    .Y(_1722_),
    .A2(net850),
    .A1(_0032_));
 sg13g2_nand2_1 _5583_ (.Y(_1723_),
    .A(_1719_),
    .B(_1722_));
 sg13g2_o21ai_1 _5584_ (.B1(_1723_),
    .Y(_1724_),
    .A1(_1703_),
    .A2(_1716_));
 sg13g2_nor2_1 _5585_ (.A(_1719_),
    .B(_1722_),
    .Y(_1725_));
 sg13g2_nor2_1 _5586_ (.A(_1716_),
    .B(_1725_),
    .Y(_1726_));
 sg13g2_nor2_1 _5587_ (.A(_1703_),
    .B(_1726_),
    .Y(_1727_));
 sg13g2_mux2_1 _5588_ (.A0(_1726_),
    .A1(_1727_),
    .S(_1724_),
    .X(_1728_));
 sg13g2_o21ai_1 _5589_ (.B1(_1728_),
    .Y(_1729_),
    .A1(_1692_),
    .A2(_1702_));
 sg13g2_xnor2_1 _5590_ (.Y(_1730_),
    .A(net953),
    .B(net951));
 sg13g2_a22oi_1 _5591_ (.Y(_1731_),
    .B1(_1360_),
    .B2(net954),
    .A2(\vgademo.b_cos[7] ),
    .A1(_3116_));
 sg13g2_o21ai_1 _5592_ (.B1(_1731_),
    .Y(_1732_),
    .A1(\vgademo.bayer_j[1] ),
    .A2(_1361_));
 sg13g2_a22oi_1 _5593_ (.Y(_1733_),
    .B1(_3161_),
    .B2(\vgademo.v_count[3] ),
    .A2(_3160_),
    .A1(\vgademo.v_count[2] ));
 sg13g2_a22oi_1 _5594_ (.Y(_1734_),
    .B1(_1732_),
    .B2(_1733_),
    .A2(\vgademo.b_cos[8] ),
    .A1(_3117_));
 sg13g2_nand2_1 _5595_ (.Y(_1735_),
    .A(net960),
    .B(_1734_));
 sg13g2_nand2_1 _5596_ (.Y(_1736_),
    .A(_3162_),
    .B(_1735_));
 sg13g2_nor2_1 _5597_ (.A(net960),
    .B(_1734_),
    .Y(_1737_));
 sg13g2_xnor2_1 _5598_ (.Y(_1738_),
    .A(_3128_),
    .B(_1730_));
 sg13g2_nor2_1 _5599_ (.A(_1737_),
    .B(_1738_),
    .Y(_1739_));
 sg13g2_a22oi_1 _5600_ (.Y(_1740_),
    .B1(_1736_),
    .B2(_1739_),
    .A2(_1730_),
    .A1(net959));
 sg13g2_nor2_1 _5601_ (.A(net953),
    .B(\vgademo.b_cos[11] ),
    .Y(_1741_));
 sg13g2_a21oi_2 _5602_ (.B1(_1741_),
    .Y(_1742_),
    .A2(_1654_),
    .A1(net953));
 sg13g2_xor2_1 _5603_ (.B(_1742_),
    .A(_0016_),
    .X(_1743_));
 sg13g2_a22oi_1 _5604_ (.Y(_1744_),
    .B1(_1742_),
    .B2(net958),
    .A2(_3142_),
    .A1(net957));
 sg13g2_o21ai_1 _5605_ (.B1(_1744_),
    .Y(_1745_),
    .A1(_1740_),
    .A2(_1743_));
 sg13g2_or2_1 _5606_ (.X(_1746_),
    .B(_1653_),
    .A(_3162_));
 sg13g2_nand3_1 _5607_ (.B(_0018_),
    .C(_1746_),
    .A(net957),
    .Y(_1747_));
 sg13g2_o21ai_1 _5608_ (.B1(_1747_),
    .Y(_1748_),
    .A1(_0018_),
    .A2(_1746_));
 sg13g2_a21oi_1 _5609_ (.A1(net953),
    .A2(_1735_),
    .Y(_1749_),
    .B1(_1737_));
 sg13g2_a21oi_1 _5610_ (.A1(net959),
    .A2(net951),
    .Y(_1750_),
    .B1(_1749_));
 sg13g2_xnor2_1 _5611_ (.Y(_1751_),
    .A(_0016_),
    .B(_1655_));
 sg13g2_o21ai_1 _5612_ (.B1(_1751_),
    .Y(_1752_),
    .A1(net959),
    .A2(net951));
 sg13g2_a22oi_1 _5613_ (.Y(_1753_),
    .B1(_1655_),
    .B2(net958),
    .A2(_1653_),
    .A1(net957));
 sg13g2_o21ai_1 _5614_ (.B1(_1753_),
    .Y(_1754_),
    .A1(_1750_),
    .A2(_1752_));
 sg13g2_o21ai_1 _5615_ (.B1(_0018_),
    .Y(_1755_),
    .A1(net957),
    .A2(_1653_));
 sg13g2_nor2_1 _5616_ (.A(net955),
    .B(_1755_),
    .Y(_1756_));
 sg13g2_a21oi_1 _5617_ (.A1(_1754_),
    .A2(_1756_),
    .Y(_1757_),
    .B1(_3240_));
 sg13g2_nand2_1 _5618_ (.Y(_1758_),
    .A(_0021_),
    .B(_1757_));
 sg13g2_a221oi_1 _5619_ (.B2(_1745_),
    .C1(net955),
    .B1(_1748_),
    .A1(\vgademo.v_count[8] ),
    .Y(_1759_),
    .A2(_1746_));
 sg13g2_nand2_2 _5620_ (.Y(_1760_),
    .A(_1758_),
    .B(_1759_));
 sg13g2_nor3_2 _5621_ (.A(net815),
    .B(net813),
    .C(_1760_),
    .Y(_1761_));
 sg13g2_or3_2 _5622_ (.A(net815),
    .B(net812),
    .C(_1760_),
    .X(_1762_));
 sg13g2_nand2_1 _5623_ (.Y(_1763_),
    .A(_3161_),
    .B(\vgademo.plane_du[5] ));
 sg13g2_a22oi_1 _5624_ (.Y(_1764_),
    .B1(_1364_),
    .B2(\vgademo.b_cos[6] ),
    .A2(_3175_),
    .A1(\vgademo.b_cos[7] ));
 sg13g2_o21ai_1 _5625_ (.B1(_1764_),
    .Y(_1765_),
    .A1(\vgademo.plane_du[3] ),
    .A2(_1366_));
 sg13g2_o21ai_1 _5626_ (.B1(_1765_),
    .Y(_1766_),
    .A1(\vgademo.b_cos[7] ),
    .A2(_3175_));
 sg13g2_o21ai_1 _5627_ (.B1(_1766_),
    .Y(_1767_),
    .A1(_3161_),
    .A2(\vgademo.plane_du[5] ));
 sg13g2_a22oi_1 _5628_ (.Y(_1768_),
    .B1(_1763_),
    .B2(_1767_),
    .A2(_3179_),
    .A1(net953));
 sg13g2_a221oi_1 _5629_ (.B2(net951),
    .C1(_1768_),
    .B1(\vgademo.plane_du[7] ),
    .A1(_3162_),
    .Y(_1769_),
    .A2(\vgademo.plane_du[6] ));
 sg13g2_xnor2_1 _5630_ (.Y(_1770_),
    .A(_0054_),
    .B(_1655_));
 sg13g2_o21ai_1 _5631_ (.B1(_1770_),
    .Y(_1771_),
    .A1(net951),
    .A2(\vgademo.plane_du[7] ));
 sg13g2_a22oi_1 _5632_ (.Y(_1772_),
    .B1(_1655_),
    .B2(\vgademo.plane_du[8] ),
    .A2(_1653_),
    .A1(\vgademo.plane_du[9] ));
 sg13g2_o21ai_1 _5633_ (.B1(_1772_),
    .Y(_1773_),
    .A1(_1769_),
    .A2(_1771_));
 sg13g2_o21ai_1 _5634_ (.B1(_1773_),
    .Y(_1774_),
    .A1(\vgademo.plane_du[9] ),
    .A2(_1653_));
 sg13g2_nand2_1 _5635_ (.Y(_1775_),
    .A(\vgademo.plane_du[7] ),
    .B(_1730_));
 sg13g2_a22oi_1 _5636_ (.Y(_1776_),
    .B1(_1763_),
    .B2(_1767_),
    .A2(_3179_),
    .A1(_3162_));
 sg13g2_a21oi_1 _5637_ (.A1(net953),
    .A2(\vgademo.plane_du[6] ),
    .Y(_1777_),
    .B1(_1776_));
 sg13g2_xor2_1 _5638_ (.B(_1730_),
    .A(_0053_),
    .X(_1778_));
 sg13g2_o21ai_1 _5639_ (.B1(_1775_),
    .Y(_1779_),
    .A1(_1777_),
    .A2(_1778_));
 sg13g2_xnor2_1 _5640_ (.Y(_1780_),
    .A(_0054_),
    .B(_1742_));
 sg13g2_a22oi_1 _5641_ (.Y(_1781_),
    .B1(_1779_),
    .B2(_1780_),
    .A2(_1742_),
    .A1(\vgademo.plane_du[8] ));
 sg13g2_nand2_1 _5642_ (.Y(_1782_),
    .A(\vgademo.plane_du[9] ),
    .B(_1746_));
 sg13g2_nor2_1 _5643_ (.A(_1781_),
    .B(_1782_),
    .Y(_1783_));
 sg13g2_or2_2 _5644_ (.X(_1784_),
    .B(_1783_),
    .A(_1774_));
 sg13g2_nor3_2 _5645_ (.A(net815),
    .B(net813),
    .C(net852),
    .Y(_1785_));
 sg13g2_or3_1 _5646_ (.A(net816),
    .B(net813),
    .C(net852),
    .X(_1786_));
 sg13g2_xor2_1 _5647_ (.B(\vgademo.plane_du[7] ),
    .A(net973),
    .X(_1787_));
 sg13g2_xnor2_1 _5648_ (.Y(_1788_),
    .A(net976),
    .B(\vgademo.plane_du[6] ));
 sg13g2_nand2_1 _5649_ (.Y(_1789_),
    .A(net979),
    .B(\vgademo.plane_du[5] ));
 sg13g2_or2_1 _5650_ (.X(_1790_),
    .B(\vgademo.plane_du[5] ),
    .A(net979));
 sg13g2_nor2_1 _5651_ (.A(_3129_),
    .B(_3175_),
    .Y(_1791_));
 sg13g2_nand3_1 _5652_ (.B(_1790_),
    .C(_1791_),
    .A(_1789_),
    .Y(_1792_));
 sg13g2_a21oi_1 _5653_ (.A1(_1789_),
    .A2(_1792_),
    .Y(_1793_),
    .B1(_1788_));
 sg13g2_a21oi_2 _5654_ (.B1(_1793_),
    .Y(_1794_),
    .A2(\vgademo.plane_du[6] ),
    .A1(net976));
 sg13g2_nand2b_1 _5655_ (.Y(_1795_),
    .B(_1787_),
    .A_N(_1794_));
 sg13g2_xnor2_1 _5656_ (.Y(_1796_),
    .A(_1787_),
    .B(_1794_));
 sg13g2_nand2_1 _5657_ (.Y(_1797_),
    .A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ));
 sg13g2_nor2_1 _5658_ (.A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ),
    .Y(_1798_));
 sg13g2_xor2_1 _5659_ (.B(\vgademo.plane_u[15] ),
    .A(\vgademo.a_cos[10] ),
    .X(_1799_));
 sg13g2_xnor2_1 _5660_ (.Y(_1800_),
    .A(\vgademo.a_cos[9] ),
    .B(\vgademo.plane_u[14] ));
 sg13g2_nand2_1 _5661_ (.Y(_1801_),
    .A(\vgademo.a_cos[8] ),
    .B(\vgademo.plane_u[13] ));
 sg13g2_xnor2_1 _5662_ (.Y(_1802_),
    .A(\vgademo.a_cos[8] ),
    .B(\vgademo.plane_u[13] ));
 sg13g2_nand2_1 _5663_ (.Y(_1803_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.plane_u[12] ));
 sg13g2_xnor2_1 _5664_ (.Y(_1804_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.plane_u[12] ));
 sg13g2_or2_1 _5665_ (.X(_1805_),
    .B(\vgademo.plane_u[10] ),
    .A(\vgademo.a_cos[5] ));
 sg13g2_nand3_1 _5666_ (.B(\vgademo.plane_u[9] ),
    .C(_1805_),
    .A(\vgademo.a_cos[4] ),
    .Y(_1806_));
 sg13g2_a22oi_1 _5667_ (.Y(_1807_),
    .B1(\vgademo.plane_u[11] ),
    .B2(\vgademo.a_cos[6] ),
    .A2(\vgademo.plane_u[10] ),
    .A1(\vgademo.a_cos[5] ));
 sg13g2_a22oi_1 _5668_ (.Y(_1808_),
    .B1(_1806_),
    .B2(_1807_),
    .A2(_3187_),
    .A1(_3156_));
 sg13g2_nand2b_1 _5669_ (.Y(_1809_),
    .B(_1808_),
    .A_N(_1804_));
 sg13g2_a21o_1 _5670_ (.A2(_1809_),
    .A1(_1803_),
    .B1(_1802_),
    .X(_1810_));
 sg13g2_a21oi_1 _5671_ (.A1(_1801_),
    .A2(_1810_),
    .Y(_1811_),
    .B1(_1800_));
 sg13g2_a21oi_2 _5672_ (.B1(_1811_),
    .Y(_1812_),
    .A2(\vgademo.plane_u[14] ),
    .A1(\vgademo.a_cos[9] ));
 sg13g2_o21ai_1 _5673_ (.B1(_1797_),
    .Y(_1813_),
    .A1(_1798_),
    .A2(_1812_));
 sg13g2_and2_1 _5674_ (.A(\vgademo.a_cos[11] ),
    .B(\vgademo.plane_u[16] ),
    .X(_1814_));
 sg13g2_xor2_1 _5675_ (.B(\vgademo.plane_u[16] ),
    .A(\vgademo.a_cos[11] ),
    .X(_1815_));
 sg13g2_xnor2_1 _5676_ (.Y(_1816_),
    .A(_1813_),
    .B(_1815_));
 sg13g2_inv_1 _5677_ (.Y(_1817_),
    .A(_1816_));
 sg13g2_xor2_1 _5678_ (.B(_1816_),
    .A(_1796_),
    .X(_1818_));
 sg13g2_o21ai_1 _5679_ (.B1(_1795_),
    .Y(_1819_),
    .A1(_3134_),
    .A2(_3181_));
 sg13g2_and2_1 _5680_ (.A(net970),
    .B(\vgademo.plane_du[8] ),
    .X(_1820_));
 sg13g2_xor2_1 _5681_ (.B(\vgademo.plane_du[8] ),
    .A(net970),
    .X(_1821_));
 sg13g2_xnor2_1 _5682_ (.Y(_1822_),
    .A(_1819_),
    .B(_1821_));
 sg13g2_nor2_1 _5683_ (.A(_1818_),
    .B(_1822_),
    .Y(_1823_));
 sg13g2_nor2_1 _5684_ (.A(_3133_),
    .B(_3185_),
    .Y(_1824_));
 sg13g2_xor2_1 _5685_ (.B(\vgademo.plane_du[9] ),
    .A(net967),
    .X(_1825_));
 sg13g2_a21o_1 _5686_ (.A2(_1821_),
    .A1(_1819_),
    .B1(_1820_),
    .X(_1826_));
 sg13g2_xor2_1 _5687_ (.B(_1826_),
    .A(_1825_),
    .X(_1827_));
 sg13g2_inv_1 _5688_ (.Y(_1828_),
    .A(_1827_));
 sg13g2_and2_1 _5689_ (.A(\vgademo.a_cos[12] ),
    .B(\vgademo.plane_u[17] ),
    .X(_1829_));
 sg13g2_a21o_1 _5690_ (.A2(_1815_),
    .A1(_1813_),
    .B1(_1814_),
    .X(_1830_));
 sg13g2_xor2_1 _5691_ (.B(\vgademo.plane_u[17] ),
    .A(\vgademo.a_cos[12] ),
    .X(_1831_));
 sg13g2_a21o_1 _5692_ (.A2(_1831_),
    .A1(_1830_),
    .B1(_1829_),
    .X(_1832_));
 sg13g2_xor2_1 _5693_ (.B(\vgademo.plane_u[18] ),
    .A(\vgademo.a_cos[13] ),
    .X(_1833_));
 sg13g2_xnor2_1 _5694_ (.Y(_1834_),
    .A(_1832_),
    .B(_1833_));
 sg13g2_nor2_1 _5695_ (.A(_1828_),
    .B(_1834_),
    .Y(_1835_));
 sg13g2_xnor2_1 _5696_ (.Y(_1836_),
    .A(_1827_),
    .B(_1834_));
 sg13g2_xnor2_1 _5697_ (.Y(_1837_),
    .A(_1830_),
    .B(_1831_));
 sg13g2_xor2_1 _5698_ (.B(_1837_),
    .A(_1822_),
    .X(_1838_));
 sg13g2_nand3_1 _5699_ (.B(_1817_),
    .C(_1838_),
    .A(_1796_),
    .Y(_1839_));
 sg13g2_o21ai_1 _5700_ (.B1(_1839_),
    .Y(_1840_),
    .A1(_1822_),
    .A2(_1837_));
 sg13g2_a21oi_1 _5701_ (.A1(_1836_),
    .A2(_1840_),
    .Y(_1841_),
    .B1(_1835_));
 sg13g2_a21o_1 _5702_ (.A2(\vgademo.plane_u[18] ),
    .A1(\vgademo.a_cos[13] ),
    .B1(_1832_),
    .X(_1842_));
 sg13g2_o21ai_1 _5703_ (.B1(_1842_),
    .Y(_1843_),
    .A1(\vgademo.a_cos[13] ),
    .A2(\vgademo.plane_u[18] ));
 sg13g2_a21oi_1 _5704_ (.A1(_1825_),
    .A2(_1826_),
    .Y(_1844_),
    .B1(_1824_));
 sg13g2_xor2_1 _5705_ (.B(\vgademo.a_cos[14] ),
    .A(net964),
    .X(_1845_));
 sg13g2_xor2_1 _5706_ (.B(\vgademo.plane_u[19] ),
    .A(\vgademo.plane_du[10] ),
    .X(_1846_));
 sg13g2_xnor2_1 _5707_ (.Y(_1847_),
    .A(_1845_),
    .B(_1846_));
 sg13g2_xnor2_1 _5708_ (.Y(_1848_),
    .A(_1844_),
    .B(_1847_));
 sg13g2_xnor2_1 _5709_ (.Y(_1849_),
    .A(_1843_),
    .B(_1848_));
 sg13g2_xnor2_1 _5710_ (.Y(_1850_),
    .A(_1841_),
    .B(_1849_));
 sg13g2_xnor2_1 _5711_ (.Y(_1851_),
    .A(_1836_),
    .B(_1840_));
 sg13g2_nor2_1 _5712_ (.A(net1033),
    .B(_1818_),
    .Y(_1852_));
 sg13g2_nand2b_1 _5713_ (.Y(_1853_),
    .B(net1029),
    .A_N(_1838_));
 sg13g2_a21o_1 _5714_ (.A2(_1817_),
    .A1(_1796_),
    .B1(_1838_),
    .X(_1854_));
 sg13g2_and2_1 _5715_ (.A(_3110_),
    .B(_1839_),
    .X(_1855_));
 sg13g2_a22oi_1 _5716_ (.Y(_1856_),
    .B1(_1854_),
    .B2(_1855_),
    .A2(_1853_),
    .A1(_1852_));
 sg13g2_o21ai_1 _5717_ (.B1(_1856_),
    .Y(_1857_),
    .A1(net1025),
    .A2(_1851_));
 sg13g2_inv_1 _5718_ (.Y(_1858_),
    .A(_1857_));
 sg13g2_a221oi_1 _5719_ (.B2(net1025),
    .C1(_1858_),
    .B1(_1851_),
    .A1(net1022),
    .Y(_1859_),
    .A2(_1850_));
 sg13g2_nor2_1 _5720_ (.A(net1022),
    .B(_1850_),
    .Y(_1860_));
 sg13g2_nand2_1 _5721_ (.Y(_1861_),
    .A(net1019),
    .B(net1018));
 sg13g2_nor3_2 _5722_ (.A(_1859_),
    .B(_1860_),
    .C(_1861_),
    .Y(_1862_));
 sg13g2_xor2_1 _5723_ (.B(_1836_),
    .A(net1038),
    .X(_1863_));
 sg13g2_xnor2_1 _5724_ (.Y(_1864_),
    .A(net1029),
    .B(_1796_));
 sg13g2_xnor2_1 _5725_ (.Y(_1865_),
    .A(_3108_),
    .B(_1816_));
 sg13g2_nand3_1 _5726_ (.B(_1864_),
    .C(_1865_),
    .A(net1018),
    .Y(_1866_));
 sg13g2_xor2_1 _5727_ (.B(_1838_),
    .A(net1033),
    .X(_1867_));
 sg13g2_nor3_2 _5728_ (.A(_1863_),
    .B(_1866_),
    .C(_1867_),
    .Y(_1868_));
 sg13g2_inv_1 _5729_ (.Y(_1869_),
    .A(_1868_));
 sg13g2_nor2_2 _5730_ (.A(_1862_),
    .B(net842),
    .Y(_1870_));
 sg13g2_nand2b_2 _5731_ (.Y(_1871_),
    .B(_1870_),
    .A_N(_1823_));
 sg13g2_nand3_1 _5732_ (.B(net810),
    .C(_1871_),
    .A(net847),
    .Y(_1872_));
 sg13g2_nand2_1 _5733_ (.Y(_1873_),
    .A(net1041),
    .B(net966));
 sg13g2_nand2_1 _5734_ (.Y(_1874_),
    .A(net969),
    .B(net1039));
 sg13g2_nand2_1 _5735_ (.Y(_1875_),
    .A(net966),
    .B(net1039));
 sg13g2_nand2_1 _5736_ (.Y(_1876_),
    .A(net1041),
    .B(net969));
 sg13g2_xor2_1 _5737_ (.B(_1876_),
    .A(_1875_),
    .X(_1877_));
 sg13g2_nand2_1 _5738_ (.Y(_1878_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1877_));
 sg13g2_o21ai_1 _5739_ (.B1(_1878_),
    .Y(_1879_),
    .A1(_1875_),
    .A2(_1876_));
 sg13g2_nand2_1 _5740_ (.Y(_1880_),
    .A(net964),
    .B(net1039));
 sg13g2_xor2_1 _5741_ (.B(_1880_),
    .A(_1873_),
    .X(_1881_));
 sg13g2_nand2_1 _5742_ (.Y(_1882_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1881_));
 sg13g2_xnor2_1 _5743_ (.Y(_1883_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1881_));
 sg13g2_nand2b_1 _5744_ (.Y(_1884_),
    .B(_1879_),
    .A_N(_1883_));
 sg13g2_xor2_1 _5745_ (.B(_1883_),
    .A(_1879_),
    .X(_1885_));
 sg13g2_o21ai_1 _5746_ (.B1(_1884_),
    .Y(_1886_),
    .A1(_3131_),
    .A2(_1885_));
 sg13g2_o21ai_1 _5747_ (.B1(_1882_),
    .Y(_1887_),
    .A1(_1873_),
    .A2(_1880_));
 sg13g2_nand2_1 _5748_ (.Y(_1888_),
    .A(net1041),
    .B(net962));
 sg13g2_nor2_1 _5749_ (.A(_1880_),
    .B(_1888_),
    .Y(_1889_));
 sg13g2_a22oi_1 _5750_ (.Y(_1890_),
    .B1(net1039),
    .B2(net962),
    .A2(net964),
    .A1(net1041));
 sg13g2_nor2_1 _5751_ (.A(_1889_),
    .B(_1890_),
    .Y(_1891_));
 sg13g2_xnor2_1 _5752_ (.Y(_1892_),
    .A(\vgademo.linelfsr[11] ),
    .B(_1891_));
 sg13g2_nand2b_1 _5753_ (.Y(_1893_),
    .B(_1887_),
    .A_N(_1892_));
 sg13g2_xor2_1 _5754_ (.B(_1892_),
    .A(_1887_),
    .X(_1894_));
 sg13g2_xnor2_1 _5755_ (.Y(_1895_),
    .A(_3130_),
    .B(_1894_));
 sg13g2_nand2b_1 _5756_ (.Y(_1896_),
    .B(_1886_),
    .A_N(_1895_));
 sg13g2_xor2_1 _5757_ (.B(_1895_),
    .A(_1886_),
    .X(_1897_));
 sg13g2_nand2_1 _5758_ (.Y(_1898_),
    .A(net971),
    .B(net1040));
 sg13g2_nand2_1 _5759_ (.Y(_1899_),
    .A(net1041),
    .B(net971));
 sg13g2_xor2_1 _5760_ (.B(_1899_),
    .A(_1874_),
    .X(_1900_));
 sg13g2_nand2_1 _5761_ (.Y(_1901_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1900_));
 sg13g2_o21ai_1 _5762_ (.B1(_1901_),
    .Y(_1902_),
    .A1(_1874_),
    .A2(_1899_));
 sg13g2_xnor2_1 _5763_ (.Y(_1903_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1877_));
 sg13g2_nand2b_1 _5764_ (.Y(_1904_),
    .B(_1902_),
    .A_N(_1903_));
 sg13g2_xor2_1 _5765_ (.B(_1903_),
    .A(_1902_),
    .X(_1905_));
 sg13g2_o21ai_1 _5766_ (.B1(_1904_),
    .Y(_1906_),
    .A1(net940),
    .A2(_1905_));
 sg13g2_xnor2_1 _5767_ (.Y(_1907_),
    .A(_3131_),
    .B(_1885_));
 sg13g2_inv_1 _5768_ (.Y(_1908_),
    .A(_1907_));
 sg13g2_xor2_1 _5769_ (.B(_1907_),
    .A(_1906_),
    .X(_1909_));
 sg13g2_xnor2_1 _5770_ (.Y(_1910_),
    .A(net940),
    .B(_1905_));
 sg13g2_nand2_1 _5771_ (.Y(_1911_),
    .A(net975),
    .B(net1040));
 sg13g2_nand2_1 _5772_ (.Y(_1912_),
    .A(net1042),
    .B(net975));
 sg13g2_xor2_1 _5773_ (.B(_1912_),
    .A(_1898_),
    .X(_1913_));
 sg13g2_nand2_1 _5774_ (.Y(_1914_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1913_));
 sg13g2_o21ai_1 _5775_ (.B1(_1914_),
    .Y(_1915_),
    .A1(_1898_),
    .A2(_1912_));
 sg13g2_xnor2_1 _5776_ (.Y(_1916_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1900_));
 sg13g2_nand2b_1 _5777_ (.Y(_1917_),
    .B(_1915_),
    .A_N(_1916_));
 sg13g2_xor2_1 _5778_ (.B(_1916_),
    .A(_1915_),
    .X(_1918_));
 sg13g2_o21ai_1 _5779_ (.B1(_1917_),
    .Y(_1919_),
    .A1(_3133_),
    .A2(_1918_));
 sg13g2_nand2b_1 _5780_ (.Y(_1920_),
    .B(_1910_),
    .A_N(_1919_));
 sg13g2_inv_1 _5781_ (.Y(_1921_),
    .A(_1920_));
 sg13g2_nand2b_1 _5782_ (.Y(_1922_),
    .B(_1919_),
    .A_N(_1910_));
 sg13g2_nand2_1 _5783_ (.Y(_1923_),
    .A(net1042),
    .B(net978));
 sg13g2_xor2_1 _5784_ (.B(_1923_),
    .A(_1911_),
    .X(_1924_));
 sg13g2_nand2_1 _5785_ (.Y(_1925_),
    .A(\vgademo.linelfsr[6] ),
    .B(_1924_));
 sg13g2_o21ai_1 _5786_ (.B1(_1925_),
    .Y(_1926_),
    .A1(_1911_),
    .A2(_1923_));
 sg13g2_xnor2_1 _5787_ (.Y(_1927_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1913_));
 sg13g2_nor2b_1 _5788_ (.A(_1927_),
    .B_N(_1926_),
    .Y(_1928_));
 sg13g2_nand2b_1 _5789_ (.Y(_1929_),
    .B(_1927_),
    .A_N(_1926_));
 sg13g2_nand2b_1 _5790_ (.Y(_1930_),
    .B(_1929_),
    .A_N(_1928_));
 sg13g2_a21o_1 _5791_ (.A2(_1929_),
    .A1(\vgademo.a_scrolly[7] ),
    .B1(_1928_),
    .X(_1931_));
 sg13g2_xnor2_1 _5792_ (.Y(_1932_),
    .A(_3133_),
    .B(_1918_));
 sg13g2_nor2b_1 _5793_ (.A(_1932_),
    .B_N(_1931_),
    .Y(_1933_));
 sg13g2_xnor2_1 _5794_ (.Y(_1934_),
    .A(_1931_),
    .B(_1932_));
 sg13g2_nor3_1 _5795_ (.A(_3129_),
    .B(_3197_),
    .C(_1923_),
    .Y(_1935_));
 sg13g2_a22oi_1 _5796_ (.Y(_1936_),
    .B1(net978),
    .B2(net1040),
    .A2(net980),
    .A1(net1042));
 sg13g2_nor2_1 _5797_ (.A(_1935_),
    .B(_1936_),
    .Y(_1937_));
 sg13g2_a21o_1 _5798_ (.A2(_1937_),
    .A1(\vgademo.linelfsr[5] ),
    .B1(_1935_),
    .X(_1938_));
 sg13g2_xnor2_1 _5799_ (.Y(_1939_),
    .A(\vgademo.linelfsr[6] ),
    .B(_1924_));
 sg13g2_nand2b_1 _5800_ (.Y(_1940_),
    .B(_1938_),
    .A_N(_1939_));
 sg13g2_xor2_1 _5801_ (.B(_1939_),
    .A(_1938_),
    .X(_1941_));
 sg13g2_o21ai_1 _5802_ (.B1(_1940_),
    .Y(_1942_),
    .A1(_3134_),
    .A2(_1941_));
 sg13g2_xor2_1 _5803_ (.B(_1930_),
    .A(net970),
    .X(_1943_));
 sg13g2_nor2b_1 _5804_ (.A(_1942_),
    .B_N(_1943_),
    .Y(_1944_));
 sg13g2_nand2b_1 _5805_ (.Y(_1945_),
    .B(_1942_),
    .A_N(_1943_));
 sg13g2_nand3_1 _5806_ (.B(net1039),
    .C(\vgademo.linelfsr[4] ),
    .A(net980),
    .Y(_1946_));
 sg13g2_a21o_1 _5807_ (.A2(net1039),
    .A1(net980),
    .B1(\vgademo.linelfsr[4] ),
    .X(_1947_));
 sg13g2_nand2_1 _5808_ (.Y(_1948_),
    .A(_1946_),
    .B(_1947_));
 sg13g2_o21ai_1 _5809_ (.B1(_1946_),
    .Y(_1949_),
    .A1(_3136_),
    .A2(_1948_));
 sg13g2_xnor2_1 _5810_ (.Y(_1950_),
    .A(\vgademo.linelfsr[5] ),
    .B(_1937_));
 sg13g2_nand2b_1 _5811_ (.Y(_1951_),
    .B(_1949_),
    .A_N(_1950_));
 sg13g2_xor2_1 _5812_ (.B(_1950_),
    .A(_1949_),
    .X(_1952_));
 sg13g2_o21ai_1 _5813_ (.B1(_1951_),
    .Y(_1953_),
    .A1(_3135_),
    .A2(_1952_));
 sg13g2_xnor2_1 _5814_ (.Y(_1954_),
    .A(_3134_),
    .B(_1941_));
 sg13g2_nor2b_1 _5815_ (.A(_1954_),
    .B_N(_1953_),
    .Y(_1955_));
 sg13g2_xnor2_1 _5816_ (.Y(_1956_),
    .A(_3135_),
    .B(_1952_));
 sg13g2_xnor2_1 _5817_ (.Y(_1957_),
    .A(_3136_),
    .B(_1948_));
 sg13g2_nand2_1 _5818_ (.Y(_1958_),
    .A(\vgademo.linelfsr[3] ),
    .B(net981));
 sg13g2_nor2_1 _5819_ (.A(_1957_),
    .B(_1958_),
    .Y(_1959_));
 sg13g2_nor2b_1 _5820_ (.A(_1956_),
    .B_N(_1959_),
    .Y(_1960_));
 sg13g2_xnor2_1 _5821_ (.Y(_1961_),
    .A(_1953_),
    .B(_1954_));
 sg13g2_a21oi_1 _5822_ (.A1(_1960_),
    .A2(_1961_),
    .Y(_1962_),
    .B1(_1955_));
 sg13g2_o21ai_1 _5823_ (.B1(_1945_),
    .Y(_1963_),
    .A1(_1944_),
    .A2(_1962_));
 sg13g2_a21oi_1 _5824_ (.A1(_1934_),
    .A2(_1963_),
    .Y(_1964_),
    .B1(_1933_));
 sg13g2_o21ai_1 _5825_ (.B1(_1922_),
    .Y(_1965_),
    .A1(_1921_),
    .A2(_1964_));
 sg13g2_nor2b_1 _5826_ (.A(_1909_),
    .B_N(_1965_),
    .Y(_1966_));
 sg13g2_a21oi_1 _5827_ (.A1(_1906_),
    .A2(_1908_),
    .Y(_1967_),
    .B1(_1966_));
 sg13g2_o21ai_1 _5828_ (.B1(_1896_),
    .Y(_1968_),
    .A1(_1897_),
    .A2(_1967_));
 sg13g2_o21ai_1 _5829_ (.B1(_1893_),
    .Y(_1969_),
    .A1(_3130_),
    .A2(_1894_));
 sg13g2_a21oi_1 _5830_ (.A1(\vgademo.linelfsr[11] ),
    .A2(_1891_),
    .Y(_1970_),
    .B1(_1889_));
 sg13g2_nand2_1 _5831_ (.Y(_1971_),
    .A(net961),
    .B(net1039));
 sg13g2_xor2_1 _5832_ (.B(_1971_),
    .A(\vgademo.linelfsr[12] ),
    .X(_1972_));
 sg13g2_xnor2_1 _5833_ (.Y(_1973_),
    .A(_1888_),
    .B(_1972_));
 sg13g2_xnor2_1 _5834_ (.Y(_1974_),
    .A(_1970_),
    .B(_1973_));
 sg13g2_xnor2_1 _5835_ (.Y(_1975_),
    .A(\vgademo.a_scrolly[12] ),
    .B(_1974_));
 sg13g2_xnor2_1 _5836_ (.Y(_1976_),
    .A(_1969_),
    .B(_1975_));
 sg13g2_xnor2_1 _5837_ (.Y(_1977_),
    .A(_1968_),
    .B(_1976_));
 sg13g2_xor2_1 _5838_ (.B(_1967_),
    .A(_1897_),
    .X(_1978_));
 sg13g2_inv_1 _5839_ (.Y(_1979_),
    .A(_1978_));
 sg13g2_xnor2_1 _5840_ (.Y(_1980_),
    .A(_1909_),
    .B(_1965_));
 sg13g2_inv_1 _5841_ (.Y(_1981_),
    .A(_1980_));
 sg13g2_xnor2_1 _5842_ (.Y(_1982_),
    .A(_1934_),
    .B(_1963_));
 sg13g2_nor2b_1 _5843_ (.A(_1944_),
    .B_N(_1945_),
    .Y(_1983_));
 sg13g2_xnor2_1 _5844_ (.Y(_1984_),
    .A(_1962_),
    .B(_1983_));
 sg13g2_xnor2_1 _5845_ (.Y(_1985_),
    .A(_1956_),
    .B(_1959_));
 sg13g2_xor2_1 _5846_ (.B(net980),
    .A(\vgademo.linelfsr[3] ),
    .X(_1986_));
 sg13g2_inv_1 _5847_ (.Y(_1987_),
    .A(_1986_));
 sg13g2_nor2_2 _5848_ (.A(_1957_),
    .B(_1987_),
    .Y(_1988_));
 sg13g2_and2_1 _5849_ (.A(_1985_),
    .B(_1988_),
    .X(_1989_));
 sg13g2_xor2_1 _5850_ (.B(_1961_),
    .A(_1960_),
    .X(_1990_));
 sg13g2_nand3_1 _5851_ (.B(_1989_),
    .C(_1990_),
    .A(_1984_),
    .Y(_1991_));
 sg13g2_nor2_1 _5852_ (.A(_1982_),
    .B(_1991_),
    .Y(_1992_));
 sg13g2_nand2_1 _5853_ (.Y(_1993_),
    .A(_1920_),
    .B(_1922_));
 sg13g2_xor2_1 _5854_ (.B(_1993_),
    .A(_1964_),
    .X(_1994_));
 sg13g2_inv_1 _5855_ (.Y(_1995_),
    .A(_1994_));
 sg13g2_nand2_1 _5856_ (.Y(_1996_),
    .A(_1992_),
    .B(_1994_));
 sg13g2_nor2_1 _5857_ (.A(_1981_),
    .B(_1996_),
    .Y(_1997_));
 sg13g2_nand2_1 _5858_ (.Y(_1998_),
    .A(_1978_),
    .B(_1997_));
 sg13g2_xnor2_1 _5859_ (.Y(_1999_),
    .A(_1980_),
    .B(_1996_));
 sg13g2_xnor2_1 _5860_ (.Y(_2000_),
    .A(_1985_),
    .B(_1988_));
 sg13g2_xor2_1 _5861_ (.B(_1958_),
    .A(_1957_),
    .X(_2001_));
 sg13g2_nor2_1 _5862_ (.A(_1986_),
    .B(_2001_),
    .Y(_2002_));
 sg13g2_nor2_1 _5863_ (.A(_1988_),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_nor3_1 _5864_ (.A(\vgademo.audio_snare_frames[3] ),
    .B(_1988_),
    .C(_2002_),
    .Y(_2004_));
 sg13g2_xnor2_1 _5865_ (.Y(_2005_),
    .A(\vgademo.audio_snare_frames[3] ),
    .B(_2003_));
 sg13g2_xnor2_1 _5866_ (.Y(_2006_),
    .A(net999),
    .B(_1986_));
 sg13g2_nand2_1 _5867_ (.Y(_2007_),
    .A(\vgademo.linelfsr[2] ),
    .B(net939));
 sg13g2_or2_1 _5868_ (.X(_2008_),
    .B(_2007_),
    .A(_2006_));
 sg13g2_o21ai_1 _5869_ (.B1(_2008_),
    .Y(_2009_),
    .A1(net999),
    .A2(_1986_));
 sg13g2_a21oi_1 _5870_ (.A1(_2005_),
    .A2(_2009_),
    .Y(_2010_),
    .B1(_2004_));
 sg13g2_nor2_1 _5871_ (.A(_2000_),
    .B(_2010_),
    .Y(_2011_));
 sg13g2_and3_1 _5872_ (.X(_2012_),
    .A(_1961_),
    .B(_1983_),
    .C(_2011_));
 sg13g2_nand4_1 _5873_ (.B(_1922_),
    .C(_1934_),
    .A(_1920_),
    .Y(_2013_),
    .D(_2012_));
 sg13g2_inv_1 _5874_ (.Y(_2014_),
    .A(_2013_));
 sg13g2_a21oi_1 _5875_ (.A1(_1999_),
    .A2(_2014_),
    .Y(_2015_),
    .B1(_1997_));
 sg13g2_nor2_1 _5876_ (.A(_1979_),
    .B(_2015_),
    .Y(_2016_));
 sg13g2_mux2_1 _5877_ (.A0(_2016_),
    .A1(_1998_),
    .S(_1977_),
    .X(_2017_));
 sg13g2_inv_1 _5878_ (.Y(_2018_),
    .A(_2017_));
 sg13g2_xnor2_1 _5879_ (.Y(_2019_),
    .A(_1978_),
    .B(_2015_));
 sg13g2_nor2_1 _5880_ (.A(_0039_),
    .B(_2019_),
    .Y(_2020_));
 sg13g2_xor2_1 _5881_ (.B(_1991_),
    .A(_1982_),
    .X(_2021_));
 sg13g2_xnor2_1 _5882_ (.Y(_2022_),
    .A(_2012_),
    .B(_2021_));
 sg13g2_nand2_1 _5883_ (.Y(_2023_),
    .A(net984),
    .B(_2022_));
 sg13g2_o21ai_1 _5884_ (.B1(_1990_),
    .Y(_2024_),
    .A1(_1989_),
    .A2(_2011_));
 sg13g2_xnor2_1 _5885_ (.Y(_2025_),
    .A(_0035_),
    .B(_1984_));
 sg13g2_xnor2_1 _5886_ (.Y(_2026_),
    .A(_2024_),
    .B(_2025_));
 sg13g2_or3_1 _5887_ (.A(_1989_),
    .B(_1990_),
    .C(_2011_),
    .X(_2027_));
 sg13g2_and2_1 _5888_ (.A(_2024_),
    .B(_2027_),
    .X(_2028_));
 sg13g2_xnor2_1 _5889_ (.Y(_2029_),
    .A(_2000_),
    .B(_2010_));
 sg13g2_xor2_1 _5890_ (.B(_2009_),
    .A(_2005_),
    .X(_2030_));
 sg13g2_nand2_1 _5891_ (.Y(_2031_),
    .A(\vgademo.h_count[0] ),
    .B(_2007_));
 sg13g2_o21ai_1 _5892_ (.B1(_2031_),
    .Y(_2032_),
    .A1(\vgademo.linelfsr[2] ),
    .A2(net939));
 sg13g2_nand2_1 _5893_ (.Y(_2033_),
    .A(net986),
    .B(_2006_));
 sg13g2_o21ai_1 _5894_ (.B1(_2032_),
    .Y(_2034_),
    .A1(net986),
    .A2(_2006_));
 sg13g2_nand3_1 _5895_ (.B(_2033_),
    .C(_2034_),
    .A(_2008_),
    .Y(_2035_));
 sg13g2_nand3b_1 _5896_ (.B(_2030_),
    .C(_2035_),
    .Y(_2036_),
    .A_N(_0033_));
 sg13g2_a21oi_1 _5897_ (.A1(_0033_),
    .A2(_2035_),
    .Y(_2037_),
    .B1(\vgademo.h_count[2] ));
 sg13g2_or2_1 _5898_ (.X(_2038_),
    .B(_2037_),
    .A(_2030_));
 sg13g2_nand2_1 _5899_ (.Y(_2039_),
    .A(net985),
    .B(_2029_));
 sg13g2_nand3_1 _5900_ (.B(_2038_),
    .C(_2039_),
    .A(_2036_),
    .Y(_2040_));
 sg13g2_o21ai_1 _5901_ (.B1(_2040_),
    .Y(_2041_),
    .A1(net985),
    .A2(_2029_));
 sg13g2_o21ai_1 _5902_ (.B1(_2041_),
    .Y(_2042_),
    .A1(_0044_),
    .A2(_2028_));
 sg13g2_a21oi_1 _5903_ (.A1(_0044_),
    .A2(_2028_),
    .Y(_2043_),
    .B1(_2026_));
 sg13g2_xor2_1 _5904_ (.B(_2024_),
    .A(_1984_),
    .X(_2044_));
 sg13g2_a22oi_1 _5905_ (.Y(_2045_),
    .B1(_2044_),
    .B2(\vgademo.h_count[5] ),
    .A2(_2043_),
    .A1(_2042_));
 sg13g2_xor2_1 _5906_ (.B(_2022_),
    .A(_0036_),
    .X(_2046_));
 sg13g2_o21ai_1 _5907_ (.B1(_2023_),
    .Y(_2047_),
    .A1(_2045_),
    .A2(_2046_));
 sg13g2_a21oi_1 _5908_ (.A1(_2012_),
    .A2(_2021_),
    .Y(_2048_),
    .B1(_1992_));
 sg13g2_xnor2_1 _5909_ (.Y(_2049_),
    .A(_1995_),
    .B(_2048_));
 sg13g2_o21ai_1 _5910_ (.B1(_2047_),
    .Y(_2050_),
    .A1(\vgademo.h_count[7] ),
    .A2(_2049_));
 sg13g2_xnor2_1 _5911_ (.Y(_2051_),
    .A(_1999_),
    .B(_2013_));
 sg13g2_nor2_1 _5912_ (.A(_0038_),
    .B(_2051_),
    .Y(_2052_));
 sg13g2_a21oi_1 _5913_ (.A1(\vgademo.h_count[7] ),
    .A2(_2049_),
    .Y(_2053_),
    .B1(_2052_));
 sg13g2_a21oi_1 _5914_ (.A1(_2050_),
    .A2(_2053_),
    .Y(_2054_),
    .B1(_2020_));
 sg13g2_a22oi_1 _5915_ (.Y(_2055_),
    .B1(_2051_),
    .B2(_0038_),
    .A2(_2019_),
    .A1(_0039_));
 sg13g2_nand2_1 _5916_ (.Y(_2056_),
    .A(_2054_),
    .B(_2055_));
 sg13g2_o21ai_1 _5917_ (.B1(_2056_),
    .Y(_2057_),
    .A1(_3126_),
    .A2(_2019_));
 sg13g2_xnor2_1 _5918_ (.Y(_2058_),
    .A(_3127_),
    .B(_2017_));
 sg13g2_a22oi_1 _5919_ (.Y(_2059_),
    .B1(_2057_),
    .B2(_2058_),
    .A2(_2018_),
    .A1(\vgademo.h_count[10] ));
 sg13g2_a21o_1 _5920_ (.A2(_2016_),
    .A1(_1977_),
    .B1(_2059_),
    .X(_2060_));
 sg13g2_a22oi_1 _5921_ (.Y(_2061_),
    .B1(_1986_),
    .B2(_3119_),
    .A2(_3120_),
    .A1(\vgademo.linelfsr[2] ));
 sg13g2_a21oi_1 _5922_ (.A1(net986),
    .A2(_1987_),
    .Y(_2062_),
    .B1(_2061_));
 sg13g2_xnor2_1 _5923_ (.Y(_2063_),
    .A(_0033_),
    .B(_2001_));
 sg13g2_nand2b_1 _5924_ (.Y(_2064_),
    .B(\vgademo.h_count[2] ),
    .A_N(_2001_));
 sg13g2_o21ai_1 _5925_ (.B1(_2064_),
    .Y(_2065_),
    .A1(_2062_),
    .A2(_2063_));
 sg13g2_nand2_1 _5926_ (.Y(_2066_),
    .A(net985),
    .B(_2065_));
 sg13g2_nand2_1 _5927_ (.Y(_2067_),
    .A(_1985_),
    .B(_2066_));
 sg13g2_o21ai_1 _5928_ (.B1(_2067_),
    .Y(_2068_),
    .A1(net985),
    .A2(_2065_));
 sg13g2_o21ai_1 _5929_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_0044_),
    .A2(_1990_));
 sg13g2_nand2_1 _5930_ (.Y(_2070_),
    .A(_0044_),
    .B(_1990_));
 sg13g2_nand3b_1 _5931_ (.B(_2069_),
    .C(_2070_),
    .Y(_2071_),
    .A_N(_2025_));
 sg13g2_o21ai_1 _5932_ (.B1(_2071_),
    .Y(_2072_),
    .A1(net941),
    .A2(_1984_));
 sg13g2_xnor2_1 _5933_ (.Y(_2073_),
    .A(_0036_),
    .B(_1982_));
 sg13g2_nand2_1 _5934_ (.Y(_2074_),
    .A(_2072_),
    .B(_2073_));
 sg13g2_a22oi_1 _5935_ (.Y(_2075_),
    .B1(_1995_),
    .B2(\vgademo.h_count[7] ),
    .A2(_1982_),
    .A1(net984));
 sg13g2_a22oi_1 _5936_ (.Y(_2076_),
    .B1(_2074_),
    .B2(_2075_),
    .A2(_1994_),
    .A1(_3125_));
 sg13g2_xor2_1 _5937_ (.B(_1980_),
    .A(_0038_),
    .X(_2077_));
 sg13g2_a22oi_1 _5938_ (.Y(_2078_),
    .B1(_2076_),
    .B2(_2077_),
    .A2(_1981_),
    .A1(net983));
 sg13g2_a21oi_1 _5939_ (.A1(_3126_),
    .A2(_1978_),
    .Y(_2079_),
    .B1(_2078_));
 sg13g2_a21oi_1 _5940_ (.A1(\vgademo.h_count[9] ),
    .A2(_1979_),
    .Y(_2080_),
    .B1(_2079_));
 sg13g2_o21ai_1 _5941_ (.B1(_2080_),
    .Y(_2081_),
    .A1(net982),
    .A2(_1977_));
 sg13g2_nor2_1 _5942_ (.A(\vgademo.v_count[8] ),
    .B(net964),
    .Y(_2082_));
 sg13g2_nor2_1 _5943_ (.A(net956),
    .B(net963),
    .Y(_2083_));
 sg13g2_xnor2_1 _5944_ (.Y(_2084_),
    .A(net956),
    .B(net963));
 sg13g2_nand2b_1 _5945_ (.Y(_2085_),
    .B(_2084_),
    .A_N(_2082_));
 sg13g2_nand2_1 _5946_ (.Y(_2086_),
    .A(net957),
    .B(net967));
 sg13g2_xor2_1 _5947_ (.B(net964),
    .A(\vgademo.v_count[8] ),
    .X(_2087_));
 sg13g2_or2_1 _5948_ (.X(_2088_),
    .B(_2087_),
    .A(_2086_));
 sg13g2_xnor2_1 _5949_ (.Y(_2089_),
    .A(net957),
    .B(net967));
 sg13g2_nor2_1 _5950_ (.A(net958),
    .B(net970),
    .Y(_2090_));
 sg13g2_nor2_1 _5951_ (.A(_2089_),
    .B(_2090_),
    .Y(_2091_));
 sg13g2_nor2_1 _5952_ (.A(net959),
    .B(net973),
    .Y(_2092_));
 sg13g2_xor2_1 _5953_ (.B(net970),
    .A(net958),
    .X(_2093_));
 sg13g2_nor2_1 _5954_ (.A(_2092_),
    .B(_2093_),
    .Y(_2094_));
 sg13g2_or2_1 _5955_ (.X(_2095_),
    .B(net976),
    .A(net960));
 sg13g2_xnor2_1 _5956_ (.Y(_2096_),
    .A(net959),
    .B(net973));
 sg13g2_or2_1 _5957_ (.X(_2097_),
    .B(_2096_),
    .A(_2095_));
 sg13g2_xnor2_1 _5958_ (.Y(_2098_),
    .A(net960),
    .B(net976));
 sg13g2_o21ai_1 _5959_ (.B1(_2098_),
    .Y(_2099_),
    .A1(\vgademo.v_count[3] ),
    .A2(net979));
 sg13g2_a21oi_1 _5960_ (.A1(\vgademo.v_count[3] ),
    .A2(net979),
    .Y(_2100_),
    .B1(_2098_));
 sg13g2_a21o_1 _5961_ (.A2(_3129_),
    .A1(_3116_),
    .B1(_2100_),
    .X(_2101_));
 sg13g2_nand2_1 _5962_ (.Y(_2102_),
    .A(_2097_),
    .B(_2099_));
 sg13g2_nor2b_1 _5963_ (.A(_2099_),
    .B_N(_2097_),
    .Y(_2103_));
 sg13g2_a21oi_1 _5964_ (.A1(_2095_),
    .A2(_2096_),
    .Y(_2104_),
    .B1(_2103_));
 sg13g2_o21ai_1 _5965_ (.B1(_2104_),
    .Y(_2105_),
    .A1(_2101_),
    .A2(_2102_));
 sg13g2_nand2_1 _5966_ (.Y(_2106_),
    .A(_2092_),
    .B(_2093_));
 sg13g2_nand2b_1 _5967_ (.Y(_2107_),
    .B(_2106_),
    .A_N(_2094_));
 sg13g2_a21oi_1 _5968_ (.A1(_2105_),
    .A2(_2106_),
    .Y(_2108_),
    .B1(_2094_));
 sg13g2_xnor2_1 _5969_ (.Y(_2109_),
    .A(_2089_),
    .B(_2090_));
 sg13g2_nor2_1 _5970_ (.A(_2108_),
    .B(_2109_),
    .Y(_2110_));
 sg13g2_nor2_1 _5971_ (.A(_2091_),
    .B(_2110_),
    .Y(_2111_));
 sg13g2_xnor2_1 _5972_ (.Y(_2112_),
    .A(_2086_),
    .B(_2087_));
 sg13g2_o21ai_1 _5973_ (.B1(_2088_),
    .Y(_2113_),
    .A1(_2111_),
    .A2(_2112_));
 sg13g2_xor2_1 _5974_ (.B(_2084_),
    .A(_2082_),
    .X(_2114_));
 sg13g2_nand2b_1 _5975_ (.Y(_2115_),
    .B(_2113_),
    .A_N(_2114_));
 sg13g2_xnor2_1 _5976_ (.Y(_2116_),
    .A(_3130_),
    .B(_2083_));
 sg13g2_a21oi_1 _5977_ (.A1(_2085_),
    .A2(_2115_),
    .Y(_2117_),
    .B1(_2116_));
 sg13g2_nor2_1 _5978_ (.A(_0019_),
    .B(_2083_),
    .Y(_2118_));
 sg13g2_nor2_1 _5979_ (.A(_2117_),
    .B(_2118_),
    .Y(_2119_));
 sg13g2_nand2b_1 _5980_ (.Y(_2120_),
    .B(_2119_),
    .A_N(\vgademo.a_scrolly[12] ));
 sg13g2_nor2b_1 _5981_ (.A(\vgademo.a_scrolly[13] ),
    .B_N(_2120_),
    .Y(_2121_));
 sg13g2_xnor2_1 _5982_ (.Y(_2122_),
    .A(_0066_),
    .B(_2121_));
 sg13g2_a22oi_1 _5983_ (.Y(_2123_),
    .B1(_2120_),
    .B2(\vgademo.a_scrolly[13] ),
    .A2(_2119_),
    .A1(_1055_));
 sg13g2_xor2_1 _5984_ (.B(_2107_),
    .A(_2105_),
    .X(_2124_));
 sg13g2_and3_1 _5985_ (.X(_2125_),
    .A(_2085_),
    .B(_2115_),
    .C(_2116_));
 sg13g2_o21ai_1 _5986_ (.B1(_2123_),
    .Y(_2126_),
    .A1(_2117_),
    .A2(_2125_));
 sg13g2_xnor2_1 _5987_ (.Y(_2127_),
    .A(_2111_),
    .B(_2112_));
 sg13g2_xnor2_1 _5988_ (.Y(_2128_),
    .A(_2108_),
    .B(_2109_));
 sg13g2_xnor2_1 _5989_ (.Y(_2129_),
    .A(_0067_),
    .B(_2119_));
 sg13g2_inv_1 _5990_ (.Y(_2130_),
    .A(_2129_));
 sg13g2_nand2_1 _5991_ (.Y(_2131_),
    .A(_2123_),
    .B(_2130_));
 sg13g2_xor2_1 _5992_ (.B(_2114_),
    .A(_2113_),
    .X(_2132_));
 sg13g2_nand2_1 _5993_ (.Y(_2133_),
    .A(_2123_),
    .B(_2132_));
 sg13g2_or4_1 _5994_ (.A(_2124_),
    .B(_2127_),
    .C(_2128_),
    .D(_2130_),
    .X(_2134_));
 sg13g2_nand3_1 _5995_ (.B(_2126_),
    .C(_2133_),
    .A(_2122_),
    .Y(_2135_));
 sg13g2_a21oi_2 _5996_ (.B1(_2135_),
    .Y(_2136_),
    .A2(_2134_),
    .A1(_2123_));
 sg13g2_a21oi_1 _5997_ (.A1(net982),
    .A2(_1977_),
    .Y(_2137_),
    .B1(_2136_));
 sg13g2_nand3_1 _5998_ (.B(_2081_),
    .C(_2137_),
    .A(_2060_),
    .Y(_2138_));
 sg13g2_nand4_1 _5999_ (.B(net966),
    .C(_1069_),
    .A(_3129_),
    .Y(_2139_),
    .D(_1220_));
 sg13g2_mux2_1 _6000_ (.A0(_0066_),
    .A1(_1221_),
    .S(_2139_),
    .X(_2140_));
 sg13g2_nor2_2 _6001_ (.A(_1058_),
    .B(_2140_),
    .Y(_2141_));
 sg13g2_inv_1 _6002_ (.Y(_2142_),
    .A(_2141_));
 sg13g2_o21ai_1 _6003_ (.B1(_2138_),
    .Y(_2143_),
    .A1(_3140_),
    .A2(_2142_));
 sg13g2_nand2_1 _6004_ (.Y(_2144_),
    .A(_2122_),
    .B(_2142_));
 sg13g2_nor2_1 _6005_ (.A(net847),
    .B(_2144_),
    .Y(_2145_));
 sg13g2_a22oi_1 _6006_ (.Y(_2146_),
    .B1(_2145_),
    .B2(_2131_),
    .A2(_2143_),
    .A1(_1354_));
 sg13g2_a21o_1 _6007_ (.A2(_2146_),
    .A1(_1872_),
    .B1(_1761_),
    .X(_2147_));
 sg13g2_and2_1 _6008_ (.A(_1380_),
    .B(_1502_),
    .X(_2148_));
 sg13g2_inv_1 _6009_ (.Y(_2149_),
    .A(_2148_));
 sg13g2_xnor2_1 _6010_ (.Y(_2150_),
    .A(_1380_),
    .B(_1502_));
 sg13g2_nand2_1 _6011_ (.Y(_2151_),
    .A(net858),
    .B(_2150_));
 sg13g2_nand2_1 _6012_ (.Y(_2152_),
    .A(_1379_),
    .B(_1497_));
 sg13g2_xnor2_1 _6013_ (.Y(_2153_),
    .A(_1378_),
    .B(_1498_));
 sg13g2_o21ai_1 _6014_ (.B1(_2152_),
    .Y(_2154_),
    .A1(_2149_),
    .A2(_2153_));
 sg13g2_xnor2_1 _6015_ (.Y(_2155_),
    .A(_1495_),
    .B(_1572_));
 sg13g2_xnor2_1 _6016_ (.Y(_2156_),
    .A(_2154_),
    .B(_2155_));
 sg13g2_a21oi_1 _6017_ (.A1(_1761_),
    .A2(_2156_),
    .Y(_2157_),
    .B1(_1328_));
 sg13g2_xnor2_1 _6018_ (.Y(_2158_),
    .A(_2148_),
    .B(_2153_));
 sg13g2_inv_1 _6019_ (.Y(_2159_),
    .A(_2158_));
 sg13g2_nor4_2 _6020_ (.A(net815),
    .B(net812),
    .C(_1760_),
    .Y(_2160_),
    .D(_2159_));
 sg13g2_a21o_1 _6021_ (.A2(_2160_),
    .A1(_2156_),
    .B1(_1328_),
    .X(_2161_));
 sg13g2_nand2_2 _6022_ (.Y(_2162_),
    .A(_2151_),
    .B(_2161_));
 sg13g2_a21oi_1 _6023_ (.A1(_2147_),
    .A2(_2162_),
    .Y(_2163_),
    .B1(_1332_));
 sg13g2_a21o_1 _6024_ (.A2(_2162_),
    .A1(_2147_),
    .B1(_1332_),
    .X(_2164_));
 sg13g2_and3_1 _6025_ (.X(_2165_),
    .A(_1762_),
    .B(_2126_),
    .C(_2145_));
 sg13g2_nand3_1 _6026_ (.B(_1816_),
    .C(_1869_),
    .A(_1796_),
    .Y(_2166_));
 sg13g2_a21o_2 _6027_ (.A2(net842),
    .A1(_0055_),
    .B1(_1862_),
    .X(_2167_));
 sg13g2_nor2b_2 _6028_ (.A(_2167_),
    .B_N(_2166_),
    .Y(_2168_));
 sg13g2_o21ai_1 _6029_ (.B1(net848),
    .Y(_2169_),
    .A1(_1785_),
    .A2(_2168_));
 sg13g2_and2_2 _6030_ (.A(_1354_),
    .B(_2138_),
    .X(_2170_));
 sg13g2_or2_1 _6031_ (.X(_2171_),
    .B(_2170_),
    .A(_1761_));
 sg13g2_nand2_1 _6032_ (.Y(_2172_),
    .A(_0075_),
    .B(_2141_));
 sg13g2_a21oi_2 _6033_ (.B1(_1761_),
    .Y(_2173_),
    .A2(_2172_),
    .A1(_2170_));
 sg13g2_a21oi_1 _6034_ (.A1(_2169_),
    .A2(_2173_),
    .Y(_2174_),
    .B1(_2165_));
 sg13g2_a221oi_1 _6035_ (.B2(_2173_),
    .C1(_2165_),
    .B1(_2169_),
    .A1(_2151_),
    .Y(_2175_),
    .A2(_2161_));
 sg13g2_nand2_1 _6036_ (.Y(_2176_),
    .A(_2162_),
    .B(_2174_));
 sg13g2_xnor2_1 _6037_ (.Y(_2177_),
    .A(\vgademo.h_count[0] ),
    .B(net980));
 sg13g2_xnor2_1 _6038_ (.Y(_2178_),
    .A(_3115_),
    .B(_2177_));
 sg13g2_xnor2_1 _6039_ (.Y(_2179_),
    .A(\vgademo.bayer_j[0] ),
    .B(net936));
 sg13g2_o21ai_1 _6040_ (.B1(_2163_),
    .Y(_2180_),
    .A1(_2176_),
    .A2(_2179_));
 sg13g2_o21ai_1 _6041_ (.B1(_2164_),
    .Y(_2181_),
    .A1(_2175_),
    .A2(_2178_));
 sg13g2_nand2_1 _6042_ (.Y(_2182_),
    .A(_2180_),
    .B(_2181_));
 sg13g2_nor4_2 _6043_ (.A(net814),
    .B(net813),
    .C(_1760_),
    .Y(_2183_),
    .D(_2156_));
 sg13g2_nand2_1 _6044_ (.Y(_2184_),
    .A(_2159_),
    .B(_2183_));
 sg13g2_a221oi_1 _6045_ (.B2(_2159_),
    .C1(_1328_),
    .B1(_2183_),
    .A1(_2156_),
    .Y(_2185_),
    .A2(_2160_));
 sg13g2_nor2_1 _6046_ (.A(_1328_),
    .B(_2150_),
    .Y(_2186_));
 sg13g2_or2_1 _6047_ (.X(_2187_),
    .B(_2186_),
    .A(_2185_));
 sg13g2_nor3_1 _6048_ (.A(_1796_),
    .B(_1816_),
    .C(net842),
    .Y(_2188_));
 sg13g2_nor2_2 _6049_ (.A(_1818_),
    .B(net842),
    .Y(_2189_));
 sg13g2_inv_1 _6050_ (.Y(_2190_),
    .A(_2189_));
 sg13g2_and3_1 _6051_ (.X(_2191_),
    .A(_1788_),
    .B(_1789_),
    .C(_1792_));
 sg13g2_nor3_1 _6052_ (.A(_1793_),
    .B(_2190_),
    .C(_2191_),
    .Y(_2192_));
 sg13g2_a21o_2 _6053_ (.A2(net842),
    .A1(_0057_),
    .B1(_1862_),
    .X(_2193_));
 sg13g2_nor2_1 _6054_ (.A(_2192_),
    .B(_2193_),
    .Y(_2194_));
 sg13g2_nor4_1 _6055_ (.A(net814),
    .B(net812),
    .C(net852),
    .D(_1871_),
    .Y(_2195_));
 sg13g2_a221oi_1 _6056_ (.B2(_2194_),
    .C1(_2195_),
    .B1(net811),
    .A1(net855),
    .Y(_2196_),
    .A2(net853));
 sg13g2_nand2_1 _6057_ (.Y(_2197_),
    .A(_0056_),
    .B(_2141_));
 sg13g2_a21oi_2 _6058_ (.B1(net847),
    .Y(_2198_),
    .A2(_2197_),
    .A1(_2138_));
 sg13g2_a21o_1 _6059_ (.A2(_2145_),
    .A1(_2133_),
    .B1(_2198_),
    .X(_2199_));
 sg13g2_o21ai_1 _6060_ (.B1(_1762_),
    .Y(_2200_),
    .A1(_2196_),
    .A2(_2199_));
 sg13g2_nand2_1 _6061_ (.Y(_2201_),
    .A(_2187_),
    .B(_2200_));
 sg13g2_a21oi_1 _6062_ (.A1(_2187_),
    .A2(_2200_),
    .Y(_2202_),
    .B1(net936));
 sg13g2_nand3_1 _6063_ (.B(_2187_),
    .C(_2200_),
    .A(net936),
    .Y(_2203_));
 sg13g2_nor2b_1 _6064_ (.A(_2202_),
    .B_N(_2203_),
    .Y(_2204_));
 sg13g2_a21oi_1 _6065_ (.A1(_2176_),
    .A2(_2203_),
    .Y(_2205_),
    .B1(_2202_));
 sg13g2_xnor2_1 _6066_ (.Y(_2206_),
    .A(_2175_),
    .B(_2179_));
 sg13g2_xnor2_1 _6067_ (.Y(_2207_),
    .A(_2163_),
    .B(_2206_));
 sg13g2_nand2_1 _6068_ (.Y(_2208_),
    .A(_2205_),
    .B(_2207_));
 sg13g2_o21ai_1 _6069_ (.B1(_2170_),
    .Y(_2209_),
    .A1(_3139_),
    .A2(_2142_));
 sg13g2_nand2_1 _6070_ (.Y(_2210_),
    .A(_1762_),
    .B(_2209_));
 sg13g2_a21oi_1 _6071_ (.A1(_2123_),
    .A2(_2127_),
    .Y(_2211_),
    .B1(_2144_));
 sg13g2_o21ai_1 _6072_ (.B1(_1762_),
    .Y(_2212_),
    .A1(_2209_),
    .A2(_2211_));
 sg13g2_nor4_1 _6073_ (.A(net814),
    .B(net812),
    .C(net852),
    .D(_2168_),
    .Y(_2213_));
 sg13g2_a21o_1 _6074_ (.A2(_1790_),
    .A1(_1789_),
    .B1(_1791_),
    .X(_2214_));
 sg13g2_nand3_1 _6075_ (.B(_2189_),
    .C(_2214_),
    .A(_1792_),
    .Y(_2215_));
 sg13g2_a21o_2 _6076_ (.A2(net842),
    .A1(_0062_),
    .B1(_1862_),
    .X(_2216_));
 sg13g2_nor2b_1 _6077_ (.A(_2216_),
    .B_N(_2215_),
    .Y(_2217_));
 sg13g2_inv_1 _6078_ (.Y(_2218_),
    .A(_2217_));
 sg13g2_a221oi_1 _6079_ (.B2(_2218_),
    .C1(_2213_),
    .B1(net810),
    .A1(net855),
    .Y(_2219_),
    .A2(net853));
 sg13g2_o21ai_1 _6080_ (.B1(_2157_),
    .Y(_2220_),
    .A1(_2212_),
    .A2(_2219_));
 sg13g2_o21ai_1 _6081_ (.B1(_2170_),
    .Y(_2221_),
    .A1(_3138_),
    .A2(_2142_));
 sg13g2_nand2_1 _6082_ (.Y(_2222_),
    .A(_1762_),
    .B(_2221_));
 sg13g2_a21oi_1 _6083_ (.A1(_2123_),
    .A2(_2128_),
    .Y(_2223_),
    .B1(_2144_));
 sg13g2_o21ai_1 _6084_ (.B1(_1762_),
    .Y(_2224_),
    .A1(_2221_),
    .A2(_2223_));
 sg13g2_nor4_1 _6085_ (.A(net814),
    .B(net812),
    .C(net852),
    .D(_2194_),
    .Y(_2225_));
 sg13g2_nor2_1 _6086_ (.A(net981),
    .B(\vgademo.plane_du[4] ),
    .Y(_2226_));
 sg13g2_or3_1 _6087_ (.A(_1791_),
    .B(_2190_),
    .C(_2226_),
    .X(_2227_));
 sg13g2_a21oi_2 _6088_ (.B1(_1862_),
    .Y(_2228_),
    .A2(net842),
    .A1(_0059_));
 sg13g2_nand2_1 _6089_ (.Y(_2229_),
    .A(_2227_),
    .B(_2228_));
 sg13g2_a221oi_1 _6090_ (.B2(_2229_),
    .C1(_2225_),
    .B1(net810),
    .A1(net855),
    .Y(_2230_),
    .A2(net853));
 sg13g2_o21ai_1 _6091_ (.B1(net858),
    .Y(_2231_),
    .A1(_2224_),
    .A2(_2230_));
 sg13g2_xor2_1 _6092_ (.B(net981),
    .A(\vgademo.h_count[2] ),
    .X(_2232_));
 sg13g2_nand2_1 _6093_ (.Y(_2233_),
    .A(_2231_),
    .B(_2232_));
 sg13g2_nor2_1 _6094_ (.A(_2231_),
    .B(_2232_),
    .Y(_2234_));
 sg13g2_a21oi_1 _6095_ (.A1(_2164_),
    .A2(_2233_),
    .Y(_2235_),
    .B1(_2234_));
 sg13g2_xor2_1 _6096_ (.B(net981),
    .A(\vgademo.h_count[1] ),
    .X(_2236_));
 sg13g2_a21oi_2 _6097_ (.B1(_1862_),
    .Y(_2237_),
    .A2(net842),
    .A1(_0058_));
 sg13g2_o21ai_1 _6098_ (.B1(_2237_),
    .Y(_2238_),
    .A1(_3173_),
    .A2(_2190_));
 sg13g2_nor4_1 _6099_ (.A(net814),
    .B(net812),
    .C(net852),
    .D(_2217_),
    .Y(_2239_));
 sg13g2_a221oi_1 _6100_ (.B2(_2238_),
    .C1(_2239_),
    .B1(net811),
    .A1(net855),
    .Y(_2240_),
    .A2(net853));
 sg13g2_a21o_1 _6101_ (.A2(_2124_),
    .A1(_2123_),
    .B1(_2144_),
    .X(_2241_));
 sg13g2_a21o_1 _6102_ (.A2(_2241_),
    .A1(_2170_),
    .B1(_1761_),
    .X(_2242_));
 sg13g2_o21ai_1 _6103_ (.B1(net858),
    .Y(_2243_),
    .A1(_2240_),
    .A2(_2242_));
 sg13g2_and2_1 _6104_ (.A(net935),
    .B(_2243_),
    .X(_2244_));
 sg13g2_or2_1 _6105_ (.X(_2245_),
    .B(_2243_),
    .A(net935));
 sg13g2_xnor2_1 _6106_ (.Y(_2246_),
    .A(net935),
    .B(_2243_));
 sg13g2_xnor2_1 _6107_ (.Y(_2247_),
    .A(_2231_),
    .B(_2246_));
 sg13g2_o21ai_1 _6108_ (.B1(_2247_),
    .Y(_2248_),
    .A1(_2220_),
    .A2(_2235_));
 sg13g2_a21o_1 _6109_ (.A2(_2245_),
    .A1(_2231_),
    .B1(_2244_),
    .X(_2249_));
 sg13g2_xnor2_1 _6110_ (.Y(_2250_),
    .A(\vgademo.bayer_j[1] ),
    .B(net935));
 sg13g2_inv_1 _6111_ (.Y(_2251_),
    .A(_2250_));
 sg13g2_and2_1 _6112_ (.A(_2220_),
    .B(_2251_),
    .X(_2252_));
 sg13g2_xnor2_1 _6113_ (.Y(_2253_),
    .A(_2220_),
    .B(_2250_));
 sg13g2_xor2_1 _6114_ (.B(_2253_),
    .A(_2201_),
    .X(_2254_));
 sg13g2_a22oi_1 _6115_ (.Y(_2255_),
    .B1(_2249_),
    .B2(_2254_),
    .A2(_2235_),
    .A1(_2220_));
 sg13g2_xnor2_1 _6116_ (.Y(_2256_),
    .A(_2176_),
    .B(_2204_));
 sg13g2_a21oi_1 _6117_ (.A1(_2201_),
    .A2(_2253_),
    .Y(_2257_),
    .B1(_2252_));
 sg13g2_nor2_1 _6118_ (.A(_2249_),
    .B(_2254_),
    .Y(_2258_));
 sg13g2_a221oi_1 _6119_ (.B2(_2257_),
    .C1(_2258_),
    .B1(_2256_),
    .A1(_2248_),
    .Y(_2259_),
    .A2(_2255_));
 sg13g2_or2_1 _6120_ (.X(_2260_),
    .B(_2207_),
    .A(_2205_));
 sg13g2_o21ai_1 _6121_ (.B1(_2260_),
    .Y(_2261_),
    .A1(_2256_),
    .A2(_2257_));
 sg13g2_o21ai_1 _6122_ (.B1(_2208_),
    .Y(_2262_),
    .A1(_2259_),
    .A2(_2261_));
 sg13g2_nor2_1 _6123_ (.A(_2182_),
    .B(_2262_),
    .Y(_2263_));
 sg13g2_nor4_1 _6124_ (.A(\vgademo.h_count[3] ),
    .B(\vgademo.h_count[2] ),
    .C(\vgademo.h_count[4] ),
    .D(\vgademo.h_count[5] ),
    .Y(_2264_));
 sg13g2_o21ai_1 _6125_ (.B1(_0577_),
    .Y(_2265_),
    .A1(_3210_),
    .A2(_2264_));
 sg13g2_nand2_2 _6126_ (.Y(_2266_),
    .A(_3127_),
    .B(_2265_));
 sg13g2_nor2_1 _6127_ (.A(\vgademo.v_count[2] ),
    .B(\vgademo.v_count[3] ),
    .Y(_2267_));
 sg13g2_nand4_1 _6128_ (.B(_3240_),
    .C(_3244_),
    .A(_3239_),
    .Y(_2268_),
    .D(_2267_));
 sg13g2_a21oi_1 _6129_ (.A1(\vgademo.v_count[8] ),
    .A2(_3242_),
    .Y(_2269_),
    .B1(net956));
 sg13g2_nand3_1 _6130_ (.B(_2268_),
    .C(_2269_),
    .A(_2266_),
    .Y(_2270_));
 sg13g2_a21oi_1 _6131_ (.A1(_2182_),
    .A2(_2262_),
    .Y(_2271_),
    .B1(_2270_));
 sg13g2_nor2b_1 _6132_ (.A(_2263_),
    .B_N(_2271_),
    .Y(_0256_));
 sg13g2_o21ai_1 _6133_ (.B1(_2180_),
    .Y(_2272_),
    .A1(_2182_),
    .A2(_2262_));
 sg13g2_nor2b_1 _6134_ (.A(_2270_),
    .B_N(_2272_),
    .Y(_0257_));
 sg13g2_nand2_1 _6135_ (.Y(_2273_),
    .A(\vgademo.a_sin[6] ),
    .B(net918));
 sg13g2_xnor2_1 _6136_ (.Y(_0258_),
    .A(net252),
    .B(_2273_));
 sg13g2_nor2_1 _6137_ (.A(net304),
    .B(net917),
    .Y(_2274_));
 sg13g2_nor2b_1 _6138_ (.A(\vgademo.a_sin[7] ),
    .B_N(\vgademo.a_cos[1] ),
    .Y(_2275_));
 sg13g2_xor2_1 _6139_ (.B(net304),
    .A(\vgademo.a_sin[7] ),
    .X(_2276_));
 sg13g2_nor2b_1 _6140_ (.A(net252),
    .B_N(\vgademo.a_sin[6] ),
    .Y(_2277_));
 sg13g2_nor2_1 _6141_ (.A(_2276_),
    .B(_2277_),
    .Y(_2278_));
 sg13g2_xnor2_1 _6142_ (.Y(_2279_),
    .A(_2276_),
    .B(_2277_));
 sg13g2_a21oi_1 _6143_ (.A1(net917),
    .A2(_2279_),
    .Y(_0259_),
    .B1(_2274_));
 sg13g2_nand2_1 _6144_ (.Y(_2280_),
    .A(_3167_),
    .B(net319));
 sg13g2_xnor2_1 _6145_ (.Y(_2281_),
    .A(\vgademo.a_sin[8] ),
    .B(\vgademo.a_cos[2] ));
 sg13g2_nor3_1 _6146_ (.A(_2275_),
    .B(_2278_),
    .C(_2281_),
    .Y(_2282_));
 sg13g2_o21ai_1 _6147_ (.B1(_2281_),
    .Y(_2283_),
    .A1(_2275_),
    .A2(_2278_));
 sg13g2_nor2b_1 _6148_ (.A(_2282_),
    .B_N(_2283_),
    .Y(_2284_));
 sg13g2_mux2_1 _6149_ (.A0(net319),
    .A1(_2284_),
    .S(net917),
    .X(_0260_));
 sg13g2_nand2_1 _6150_ (.Y(_2285_),
    .A(net372),
    .B(net912));
 sg13g2_nor2b_1 _6151_ (.A(\vgademo.a_sin[9] ),
    .B_N(\vgademo.a_cos[3] ),
    .Y(_2286_));
 sg13g2_xor2_1 _6152_ (.B(\vgademo.a_sin[9] ),
    .A(\vgademo.a_cos[3] ),
    .X(_2287_));
 sg13g2_nand3_1 _6153_ (.B(_2283_),
    .C(_2287_),
    .A(_2280_),
    .Y(_2288_));
 sg13g2_a21oi_2 _6154_ (.B1(_2287_),
    .Y(_2289_),
    .A2(_2283_),
    .A1(_2280_));
 sg13g2_nand2_1 _6155_ (.Y(_2290_),
    .A(net917),
    .B(_2288_));
 sg13g2_o21ai_1 _6156_ (.B1(_2285_),
    .Y(_0261_),
    .A1(_2289_),
    .A2(_2290_));
 sg13g2_xnor2_1 _6157_ (.Y(_2291_),
    .A(\vgademo.a_cos[4] ),
    .B(\vgademo.a_sin[10] ));
 sg13g2_o21ai_1 _6158_ (.B1(_2291_),
    .Y(_2292_),
    .A1(_2286_),
    .A2(_2289_));
 sg13g2_or3_1 _6159_ (.A(_2286_),
    .B(_2289_),
    .C(_2291_),
    .X(_2293_));
 sg13g2_a21oi_1 _6160_ (.A1(_2292_),
    .A2(_2293_),
    .Y(_2294_),
    .B1(net913));
 sg13g2_a21oi_1 _6161_ (.A1(_3154_),
    .A2(net913),
    .Y(_0262_),
    .B1(_2294_));
 sg13g2_o21ai_1 _6162_ (.B1(_2292_),
    .Y(_2295_),
    .A1(_3154_),
    .A2(\vgademo.a_sin[10] ));
 sg13g2_nand2b_1 _6163_ (.Y(_2296_),
    .B(\vgademo.a_sin[11] ),
    .A_N(\vgademo.a_cos[5] ));
 sg13g2_nor2b_1 _6164_ (.A(\vgademo.a_sin[11] ),
    .B_N(\vgademo.a_cos[5] ),
    .Y(_2297_));
 sg13g2_xnor2_1 _6165_ (.Y(_2298_),
    .A(\vgademo.a_cos[5] ),
    .B(\vgademo.a_sin[11] ));
 sg13g2_o21ai_1 _6166_ (.B1(net919),
    .Y(_2299_),
    .A1(_2295_),
    .A2(_2298_));
 sg13g2_a21oi_1 _6167_ (.A1(_2295_),
    .A2(_2298_),
    .Y(_2300_),
    .B1(_2299_));
 sg13g2_a21o_1 _6168_ (.A2(net913),
    .A1(net527),
    .B1(_2300_),
    .X(_0263_));
 sg13g2_xor2_1 _6169_ (.B(\vgademo.a_sin[12] ),
    .A(\vgademo.a_cos[6] ),
    .X(_2301_));
 sg13g2_a21oi_1 _6170_ (.A1(_2295_),
    .A2(_2296_),
    .Y(_2302_),
    .B1(_2297_));
 sg13g2_nor2_1 _6171_ (.A(_2301_),
    .B(_2302_),
    .Y(_2303_));
 sg13g2_xor2_1 _6172_ (.B(_2302_),
    .A(_2301_),
    .X(_2304_));
 sg13g2_and2_1 _6173_ (.A(net917),
    .B(_2304_),
    .X(_2305_));
 sg13g2_a21o_1 _6174_ (.A2(net912),
    .A1(net494),
    .B1(_2305_),
    .X(_0264_));
 sg13g2_a21oi_1 _6175_ (.A1(\vgademo.a_cos[6] ),
    .A2(_3170_),
    .Y(_2306_),
    .B1(_2303_));
 sg13g2_xnor2_1 _6176_ (.Y(_2307_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.a_sin[13] ));
 sg13g2_nand2b_1 _6177_ (.Y(_2308_),
    .B(_2307_),
    .A_N(_2306_));
 sg13g2_xnor2_1 _6178_ (.Y(_2309_),
    .A(_2306_),
    .B(_2307_));
 sg13g2_nor2_1 _6179_ (.A(net911),
    .B(_2309_),
    .Y(_2310_));
 sg13g2_a21oi_1 _6180_ (.A1(_3159_),
    .A2(net910),
    .Y(_0265_),
    .B1(_2310_));
 sg13g2_xnor2_1 _6181_ (.Y(_2311_),
    .A(\vgademo.a_cos[8] ),
    .B(\vgademo.a_sin[14] ));
 sg13g2_o21ai_1 _6182_ (.B1(_2308_),
    .Y(_2312_),
    .A1(_3159_),
    .A2(\vgademo.a_sin[13] ));
 sg13g2_and2_1 _6183_ (.A(_2311_),
    .B(_2312_),
    .X(_2313_));
 sg13g2_xor2_1 _6184_ (.B(_2312_),
    .A(_2311_),
    .X(_2314_));
 sg13g2_mux2_1 _6185_ (.A0(net559),
    .A1(_2314_),
    .S(net918),
    .X(_0266_));
 sg13g2_nor2_1 _6186_ (.A(net525),
    .B(net916),
    .Y(_2315_));
 sg13g2_xnor2_1 _6187_ (.Y(_2316_),
    .A(\vgademo.a_cos[9] ),
    .B(\vgademo.a_sin[14] ));
 sg13g2_a21oi_1 _6188_ (.A1(\vgademo.a_cos[8] ),
    .A2(_3171_),
    .Y(_2317_),
    .B1(_2313_));
 sg13g2_xor2_1 _6189_ (.B(_2317_),
    .A(_2316_),
    .X(_2318_));
 sg13g2_a21oi_1 _6190_ (.A1(net916),
    .A2(_2318_),
    .Y(_0267_),
    .B1(_2315_));
 sg13g2_nor2_1 _6191_ (.A(\vgademo.a_cos[10] ),
    .B(_3171_),
    .Y(_2319_));
 sg13g2_nand2_1 _6192_ (.Y(_2320_),
    .A(\vgademo.a_cos[10] ),
    .B(_3171_));
 sg13g2_nor2b_1 _6193_ (.A(_2319_),
    .B_N(_2320_),
    .Y(_2321_));
 sg13g2_and2_1 _6194_ (.A(_2313_),
    .B(_2316_),
    .X(_2322_));
 sg13g2_o21ai_1 _6195_ (.B1(_3171_),
    .Y(_2323_),
    .A1(\vgademo.a_cos[8] ),
    .A2(\vgademo.a_cos[9] ));
 sg13g2_nor2b_1 _6196_ (.A(_2322_),
    .B_N(_2323_),
    .Y(_2324_));
 sg13g2_xnor2_1 _6197_ (.Y(_2325_),
    .A(_2321_),
    .B(_2324_));
 sg13g2_mux2_1 _6198_ (.A0(net483),
    .A1(_2325_),
    .S(net919),
    .X(_0268_));
 sg13g2_nor2_1 _6199_ (.A(net438),
    .B(net916),
    .Y(_2326_));
 sg13g2_o21ai_1 _6200_ (.B1(_2320_),
    .Y(_2327_),
    .A1(_2319_),
    .A2(_2324_));
 sg13g2_xnor2_1 _6201_ (.Y(_2328_),
    .A(\vgademo.a_cos[11] ),
    .B(\vgademo.a_sin[14] ));
 sg13g2_xnor2_1 _6202_ (.Y(_2329_),
    .A(_2327_),
    .B(_2328_));
 sg13g2_a21oi_1 _6203_ (.A1(net916),
    .A2(_2329_),
    .Y(_0269_),
    .B1(_2326_));
 sg13g2_nor2b_1 _6204_ (.A(\vgademo.a_sin[14] ),
    .B_N(\vgademo.a_cos[12] ),
    .Y(_2330_));
 sg13g2_nand2b_1 _6205_ (.Y(_2331_),
    .B(\vgademo.a_sin[14] ),
    .A_N(\vgademo.a_cos[12] ));
 sg13g2_nand2b_1 _6206_ (.Y(_2332_),
    .B(_2331_),
    .A_N(_2330_));
 sg13g2_nand3_1 _6207_ (.B(_2322_),
    .C(_2328_),
    .A(_2321_),
    .Y(_2333_));
 sg13g2_o21ai_1 _6208_ (.B1(_3171_),
    .Y(_2334_),
    .A1(\vgademo.a_cos[10] ),
    .A2(\vgademo.a_cos[11] ));
 sg13g2_nand3_1 _6209_ (.B(_2333_),
    .C(_2334_),
    .A(_2323_),
    .Y(_2335_));
 sg13g2_xnor2_1 _6210_ (.Y(_2336_),
    .A(_2332_),
    .B(_2335_));
 sg13g2_mux2_1 _6211_ (.A0(net356),
    .A1(_2336_),
    .S(net916),
    .X(_0270_));
 sg13g2_nor2_1 _6212_ (.A(net215),
    .B(net916),
    .Y(_2337_));
 sg13g2_a21oi_1 _6213_ (.A1(_2331_),
    .A2(_2335_),
    .Y(_2338_),
    .B1(_2330_));
 sg13g2_nor2_1 _6214_ (.A(\vgademo.a_cos[13] ),
    .B(_3171_),
    .Y(_2339_));
 sg13g2_nand2_1 _6215_ (.Y(_2340_),
    .A(\vgademo.a_cos[13] ),
    .B(_3171_));
 sg13g2_nor2b_1 _6216_ (.A(_2339_),
    .B_N(_2340_),
    .Y(_2341_));
 sg13g2_xnor2_1 _6217_ (.Y(_2342_),
    .A(_2338_),
    .B(_2341_));
 sg13g2_a21oi_1 _6218_ (.A1(net916),
    .A2(_2342_),
    .Y(_0271_),
    .B1(_2337_));
 sg13g2_nand2_1 _6219_ (.Y(_2343_),
    .A(net464),
    .B(net914));
 sg13g2_o21ai_1 _6220_ (.B1(_2340_),
    .Y(_2344_),
    .A1(_2338_),
    .A2(_2339_));
 sg13g2_xnor2_1 _6221_ (.Y(_2345_),
    .A(\vgademo.a_cos[14] ),
    .B(\vgademo.a_sin[14] ));
 sg13g2_xnor2_1 _6222_ (.Y(_2346_),
    .A(_2344_),
    .B(_2345_));
 sg13g2_inv_1 _6223_ (.Y(_2347_),
    .A(net823));
 sg13g2_o21ai_1 _6224_ (.B1(_2343_),
    .Y(_0272_),
    .A1(net914),
    .A2(net823));
 sg13g2_xor2_1 _6225_ (.B(_2305_),
    .A(net218),
    .X(_0273_));
 sg13g2_nand2_1 _6226_ (.Y(_2348_),
    .A(net218),
    .B(_2304_));
 sg13g2_xnor2_1 _6227_ (.Y(_2349_),
    .A(\vgademo.a_sin[1] ),
    .B(_2309_));
 sg13g2_nor2_1 _6228_ (.A(_2348_),
    .B(_2349_),
    .Y(_2350_));
 sg13g2_nand2_1 _6229_ (.Y(_2351_),
    .A(net294),
    .B(net911));
 sg13g2_a21o_1 _6230_ (.A2(_2349_),
    .A1(_2348_),
    .B1(net910),
    .X(_2352_));
 sg13g2_o21ai_1 _6231_ (.B1(_2351_),
    .Y(_0274_),
    .A1(_2350_),
    .A2(_2352_));
 sg13g2_and2_1 _6232_ (.A(\vgademo.a_sin[2] ),
    .B(_2314_),
    .X(_2353_));
 sg13g2_xnor2_1 _6233_ (.Y(_2354_),
    .A(\vgademo.a_sin[2] ),
    .B(_2314_));
 sg13g2_a21oi_1 _6234_ (.A1(\vgademo.a_sin[1] ),
    .A2(_2309_),
    .Y(_2355_),
    .B1(_2350_));
 sg13g2_nor2_1 _6235_ (.A(_2354_),
    .B(_2355_),
    .Y(_2356_));
 sg13g2_nand2_1 _6236_ (.Y(_2357_),
    .A(net300),
    .B(net910));
 sg13g2_a21o_1 _6237_ (.A2(_2355_),
    .A1(_2354_),
    .B1(net910),
    .X(_2358_));
 sg13g2_o21ai_1 _6238_ (.B1(_2357_),
    .Y(_0275_),
    .A1(_2356_),
    .A2(_2358_));
 sg13g2_or2_1 _6239_ (.X(_2359_),
    .B(_2318_),
    .A(_3164_));
 sg13g2_xnor2_1 _6240_ (.Y(_2360_),
    .A(\vgademo.a_sin[3] ),
    .B(_2318_));
 sg13g2_o21ai_1 _6241_ (.B1(_2360_),
    .Y(_2361_),
    .A1(_2353_),
    .A2(_2356_));
 sg13g2_or3_1 _6242_ (.A(_2353_),
    .B(_2356_),
    .C(_2360_),
    .X(_2362_));
 sg13g2_a21oi_1 _6243_ (.A1(_2361_),
    .A2(_2362_),
    .Y(_2363_),
    .B1(net910));
 sg13g2_a21oi_1 _6244_ (.A1(_3164_),
    .A2(net910),
    .Y(_0276_),
    .B1(_2363_));
 sg13g2_and2_1 _6245_ (.A(\vgademo.a_sin[4] ),
    .B(_2325_),
    .X(_2364_));
 sg13g2_xnor2_1 _6246_ (.Y(_2365_),
    .A(\vgademo.a_sin[4] ),
    .B(_2325_));
 sg13g2_a21oi_1 _6247_ (.A1(_2359_),
    .A2(_2361_),
    .Y(_2366_),
    .B1(_2365_));
 sg13g2_nand3_1 _6248_ (.B(_2361_),
    .C(_2365_),
    .A(_2359_),
    .Y(_2367_));
 sg13g2_nand2_1 _6249_ (.Y(_2368_),
    .A(net366),
    .B(net914));
 sg13g2_nand2_1 _6250_ (.Y(_2369_),
    .A(net916),
    .B(_2367_));
 sg13g2_o21ai_1 _6251_ (.B1(_2368_),
    .Y(_0277_),
    .A1(_2366_),
    .A2(_2369_));
 sg13g2_nand2b_1 _6252_ (.Y(_2370_),
    .B(\vgademo.a_sin[5] ),
    .A_N(_2329_));
 sg13g2_xnor2_1 _6253_ (.Y(_2371_),
    .A(\vgademo.a_sin[5] ),
    .B(_2329_));
 sg13g2_o21ai_1 _6254_ (.B1(_2371_),
    .Y(_2372_),
    .A1(_2364_),
    .A2(_2366_));
 sg13g2_or3_1 _6255_ (.A(_2364_),
    .B(_2366_),
    .C(_2371_),
    .X(_2373_));
 sg13g2_a21oi_1 _6256_ (.A1(_2372_),
    .A2(_2373_),
    .Y(_2374_),
    .B1(net914));
 sg13g2_a21oi_1 _6257_ (.A1(_3165_),
    .A2(net914),
    .Y(_0278_),
    .B1(_2374_));
 sg13g2_and2_1 _6258_ (.A(\vgademo.a_sin[6] ),
    .B(_2336_),
    .X(_2375_));
 sg13g2_xnor2_1 _6259_ (.Y(_2376_),
    .A(\vgademo.a_sin[6] ),
    .B(_2336_));
 sg13g2_a21oi_1 _6260_ (.A1(_2370_),
    .A2(_2372_),
    .Y(_2377_),
    .B1(_2376_));
 sg13g2_nand3_1 _6261_ (.B(_2372_),
    .C(_2376_),
    .A(_2370_),
    .Y(_2378_));
 sg13g2_nand2_1 _6262_ (.Y(_2379_),
    .A(net479),
    .B(net910));
 sg13g2_nand2_1 _6263_ (.Y(_2380_),
    .A(net918),
    .B(_2378_));
 sg13g2_o21ai_1 _6264_ (.B1(_2379_),
    .Y(_0279_),
    .A1(_2377_),
    .A2(_2380_));
 sg13g2_nand2_1 _6265_ (.Y(_2381_),
    .A(net448),
    .B(_2342_));
 sg13g2_xnor2_1 _6266_ (.Y(_2382_),
    .A(_3166_),
    .B(_2342_));
 sg13g2_o21ai_1 _6267_ (.B1(_2382_),
    .Y(_2383_),
    .A1(_2375_),
    .A2(_2377_));
 sg13g2_or3_1 _6268_ (.A(_2375_),
    .B(_2377_),
    .C(_2382_),
    .X(_2384_));
 sg13g2_a21oi_1 _6269_ (.A1(_2383_),
    .A2(_2384_),
    .Y(_2385_),
    .B1(net911));
 sg13g2_a21oi_1 _6270_ (.A1(_3166_),
    .A2(net910),
    .Y(_0280_),
    .B1(_2385_));
 sg13g2_xnor2_1 _6271_ (.Y(_2386_),
    .A(_3167_),
    .B(net823));
 sg13g2_a21oi_1 _6272_ (.A1(_2381_),
    .A2(_2383_),
    .Y(_2387_),
    .B1(_2386_));
 sg13g2_nand3_1 _6273_ (.B(_2383_),
    .C(_2386_),
    .A(_2381_),
    .Y(_2388_));
 sg13g2_nand3b_1 _6274_ (.B(_2388_),
    .C(net917),
    .Y(_2389_),
    .A_N(_2387_));
 sg13g2_o21ai_1 _6275_ (.B1(_2389_),
    .Y(_0281_),
    .A1(_3167_),
    .A2(net917));
 sg13g2_nand2_1 _6276_ (.Y(_2390_),
    .A(net466),
    .B(net912));
 sg13g2_xnor2_1 _6277_ (.Y(_2391_),
    .A(\vgademo.a_sin[9] ),
    .B(net823));
 sg13g2_a21oi_1 _6278_ (.A1(\vgademo.a_sin[8] ),
    .A2(_2347_),
    .Y(_2392_),
    .B1(_2387_));
 sg13g2_xor2_1 _6279_ (.B(_2392_),
    .A(_2391_),
    .X(_2393_));
 sg13g2_o21ai_1 _6280_ (.B1(_2390_),
    .Y(_0282_),
    .A1(net912),
    .A2(_2393_));
 sg13g2_xnor2_1 _6281_ (.Y(_2394_),
    .A(\vgademo.a_sin[10] ),
    .B(net822));
 sg13g2_a21oi_2 _6282_ (.B1(net822),
    .Y(_2395_),
    .A2(_3168_),
    .A1(_3167_));
 sg13g2_and2_1 _6283_ (.A(_2387_),
    .B(_2391_),
    .X(_2396_));
 sg13g2_o21ai_1 _6284_ (.B1(_2394_),
    .Y(_2397_),
    .A1(_2395_),
    .A2(_2396_));
 sg13g2_or3_1 _6285_ (.A(_2394_),
    .B(_2395_),
    .C(_2396_),
    .X(_2398_));
 sg13g2_a21oi_1 _6286_ (.A1(_2397_),
    .A2(_2398_),
    .Y(_2399_),
    .B1(net912));
 sg13g2_a21oi_1 _6287_ (.A1(_3169_),
    .A2(net912),
    .Y(_0283_),
    .B1(_2399_));
 sg13g2_nand2_1 _6288_ (.Y(_2400_),
    .A(net488),
    .B(net912));
 sg13g2_xnor2_1 _6289_ (.Y(_2401_),
    .A(\vgademo.a_sin[11] ),
    .B(net822));
 sg13g2_o21ai_1 _6290_ (.B1(_2397_),
    .Y(_2402_),
    .A1(_3169_),
    .A2(net822));
 sg13g2_xnor2_1 _6291_ (.Y(_2403_),
    .A(_2401_),
    .B(_2402_));
 sg13g2_o21ai_1 _6292_ (.B1(_2400_),
    .Y(_0284_),
    .A1(net912),
    .A2(_2403_));
 sg13g2_nor2_1 _6293_ (.A(net486),
    .B(net918),
    .Y(_2404_));
 sg13g2_nand3_1 _6294_ (.B(_2396_),
    .C(_2401_),
    .A(_2394_),
    .Y(_2405_));
 sg13g2_o21ai_1 _6295_ (.B1(_2347_),
    .Y(_2406_),
    .A1(\vgademo.a_sin[10] ),
    .A2(\vgademo.a_sin[11] ));
 sg13g2_nand2_1 _6296_ (.Y(_2407_),
    .A(_2405_),
    .B(_2406_));
 sg13g2_nor2_2 _6297_ (.A(_2395_),
    .B(_2407_),
    .Y(_2408_));
 sg13g2_xnor2_1 _6298_ (.Y(_2409_),
    .A(_3170_),
    .B(net822));
 sg13g2_xnor2_1 _6299_ (.Y(_2410_),
    .A(_2408_),
    .B(_2409_));
 sg13g2_a21oi_1 _6300_ (.A1(net917),
    .A2(_2410_),
    .Y(_0285_),
    .B1(_2404_));
 sg13g2_o21ai_1 _6301_ (.B1(_2408_),
    .Y(_2411_),
    .A1(net486),
    .A2(net822));
 sg13g2_a21o_1 _6302_ (.A2(net822),
    .A1(net490),
    .B1(_2408_),
    .X(_2412_));
 sg13g2_nand3_1 _6303_ (.B(_2411_),
    .C(_2412_),
    .A(_0591_),
    .Y(_2413_));
 sg13g2_xnor2_1 _6304_ (.Y(_0286_),
    .A(net467),
    .B(_2413_));
 sg13g2_xor2_1 _6305_ (.B(net822),
    .A(net589),
    .X(_2414_));
 sg13g2_nor2_1 _6306_ (.A(_2413_),
    .B(_2414_),
    .Y(_2415_));
 sg13g2_xnor2_1 _6307_ (.Y(_0287_),
    .A(_3171_),
    .B(_2415_));
 sg13g2_and4_2 _6308_ (.A(\vgademo.h_count[10] ),
    .B(net1051),
    .C(_0576_),
    .D(_0577_),
    .X(_2416_));
 sg13g2_mux2_1 _6309_ (.A0(net315),
    .A1(_0498_),
    .S(net891),
    .X(_0288_));
 sg13g2_mux2_1 _6310_ (.A0(net348),
    .A1(_0513_),
    .S(net891),
    .X(_0289_));
 sg13g2_mux2_1 _6311_ (.A0(net354),
    .A1(_0527_),
    .S(net891),
    .X(_0290_));
 sg13g2_mux2_1 _6312_ (.A0(net505),
    .A1(_0541_),
    .S(net891),
    .X(_0291_));
 sg13g2_mux2_1 _6313_ (.A0(net485),
    .A1(_0554_),
    .S(net891),
    .X(_0292_));
 sg13g2_mux2_1 _6314_ (.A0(net352),
    .A1(_0560_),
    .S(net891),
    .X(_0293_));
 sg13g2_nor2_1 _6315_ (.A(net417),
    .B(net891),
    .Y(_2417_));
 sg13g2_a21oi_1 _6316_ (.A1(_0559_),
    .A2(net891),
    .Y(_0294_),
    .B1(_2417_));
 sg13g2_o21ai_1 _6317_ (.B1(net925),
    .Y(_2418_),
    .A1(\vgademo.b_sin[7] ),
    .A2(net900));
 sg13g2_nand2b_1 _6318_ (.Y(_2419_),
    .B(\vgademo.b_sin[7] ),
    .A_N(net285));
 sg13g2_nor2_1 _6319_ (.A(net900),
    .B(net923),
    .Y(_2420_));
 sg13g2_nand2_1 _6320_ (.Y(_2421_),
    .A(net894),
    .B(_0581_));
 sg13g2_a22oi_1 _6321_ (.Y(_2422_),
    .B1(_2418_),
    .B2(net285),
    .A2(net887),
    .A1(\vgademo.a_cos[3] ));
 sg13g2_o21ai_1 _6322_ (.B1(net286),
    .Y(_0295_),
    .A1(_2419_),
    .A2(_2421_));
 sg13g2_nor2b_1 _6323_ (.A(\vgademo.b_sin[8] ),
    .B_N(\vgademo.b_cos[1] ),
    .Y(_2423_));
 sg13g2_xnor2_1 _6324_ (.Y(_2424_),
    .A(net335),
    .B(\vgademo.b_sin[8] ));
 sg13g2_xnor2_1 _6325_ (.Y(_2425_),
    .A(_2419_),
    .B(_2424_));
 sg13g2_nor2_1 _6326_ (.A(net335),
    .B(net925),
    .Y(_2426_));
 sg13g2_a221oi_1 _6327_ (.B2(_2425_),
    .C1(_2426_),
    .B1(_2420_),
    .A1(_3154_),
    .Y(_0296_),
    .A2(net887));
 sg13g2_nand2b_1 _6328_ (.Y(_2427_),
    .B(net887),
    .A_N(\vgademo.a_cos[5] ));
 sg13g2_a21oi_1 _6329_ (.A1(_2419_),
    .A2(_2424_),
    .Y(_2428_),
    .B1(_2423_));
 sg13g2_xnor2_1 _6330_ (.Y(_2429_),
    .A(net431),
    .B(\vgademo.b_sin[9] ));
 sg13g2_nor2b_1 _6331_ (.A(_2428_),
    .B_N(_2429_),
    .Y(_2430_));
 sg13g2_xor2_1 _6332_ (.B(_2429_),
    .A(_2428_),
    .X(_2431_));
 sg13g2_o21ai_1 _6333_ (.B1(_2427_),
    .Y(_2432_),
    .A1(net431),
    .A2(_0581_));
 sg13g2_a21oi_1 _6334_ (.A1(_2420_),
    .A2(_2431_),
    .Y(_0297_),
    .B1(net432));
 sg13g2_nor2b_1 _6335_ (.A(\vgademo.b_sin[10] ),
    .B_N(\vgademo.b_cos[3] ),
    .Y(_2433_));
 sg13g2_xnor2_1 _6336_ (.Y(_2434_),
    .A(\vgademo.b_cos[3] ),
    .B(\vgademo.b_sin[10] ));
 sg13g2_a21oi_1 _6337_ (.A1(\vgademo.b_cos[2] ),
    .A2(_3155_),
    .Y(_2435_),
    .B1(_2430_));
 sg13g2_nor2b_1 _6338_ (.A(_2435_),
    .B_N(_2434_),
    .Y(_2436_));
 sg13g2_xor2_1 _6339_ (.B(_2435_),
    .A(_2434_),
    .X(_2437_));
 sg13g2_nor2_1 _6340_ (.A(net344),
    .B(net925),
    .Y(_2438_));
 sg13g2_a221oi_1 _6341_ (.B2(_2437_),
    .C1(_2438_),
    .B1(net883),
    .A1(_3156_),
    .Y(_0298_),
    .A2(net886));
 sg13g2_xnor2_1 _6342_ (.Y(_2439_),
    .A(\vgademo.b_cos[4] ),
    .B(net947));
 sg13g2_o21ai_1 _6343_ (.B1(_2439_),
    .Y(_2440_),
    .A1(_2433_),
    .A2(_2436_));
 sg13g2_or3_1 _6344_ (.A(_2433_),
    .B(_2436_),
    .C(_2439_),
    .X(_2441_));
 sg13g2_nand3_1 _6345_ (.B(_2440_),
    .C(_2441_),
    .A(net893),
    .Y(_2442_));
 sg13g2_a21oi_1 _6346_ (.A1(\vgademo.a_cos[7] ),
    .A2(net900),
    .Y(_2443_),
    .B1(net922));
 sg13g2_a22oi_1 _6347_ (.Y(_0299_),
    .B1(_2442_),
    .B2(_2443_),
    .A2(net922),
    .A1(_3157_));
 sg13g2_xor2_1 _6348_ (.B(\vgademo.b_cos[5] ),
    .A(net947),
    .X(_2444_));
 sg13g2_o21ai_1 _6349_ (.B1(_2440_),
    .Y(_2445_),
    .A1(_3157_),
    .A2(net947));
 sg13g2_nand2_1 _6350_ (.Y(_2446_),
    .A(\vgademo.a_cos[8] ),
    .B(net925));
 sg13g2_xor2_1 _6351_ (.B(_2445_),
    .A(_2444_),
    .X(_2447_));
 sg13g2_a22oi_1 _6352_ (.Y(_2448_),
    .B1(_2447_),
    .B2(net893),
    .A2(_2446_),
    .A1(net882));
 sg13g2_a21o_1 _6353_ (.A2(net921),
    .A1(net546),
    .B1(_2448_),
    .X(_0300_));
 sg13g2_xor2_1 _6354_ (.B(net954),
    .A(net946),
    .X(_2449_));
 sg13g2_o21ai_1 _6355_ (.B1(_3158_),
    .Y(_2450_),
    .A1(\vgademo.b_cos[4] ),
    .A2(\vgademo.b_cos[5] ));
 sg13g2_or2_1 _6356_ (.X(_2451_),
    .B(_2444_),
    .A(_2440_));
 sg13g2_a21oi_1 _6357_ (.A1(_2450_),
    .A2(_2451_),
    .Y(_2452_),
    .B1(_2449_));
 sg13g2_nand3_1 _6358_ (.B(_2450_),
    .C(_2451_),
    .A(_2449_),
    .Y(_2453_));
 sg13g2_nand2_1 _6359_ (.Y(_2454_),
    .A(net883),
    .B(_2453_));
 sg13g2_a22oi_1 _6360_ (.Y(_2455_),
    .B1(net886),
    .B2(net525),
    .A2(net922),
    .A1(net954));
 sg13g2_o21ai_1 _6361_ (.B1(_2455_),
    .Y(_0301_),
    .A1(_2452_),
    .A2(_2454_));
 sg13g2_xor2_1 _6362_ (.B(\vgademo.b_cos[7] ),
    .A(net946),
    .X(_2456_));
 sg13g2_a21oi_1 _6363_ (.A1(_3158_),
    .A2(net954),
    .Y(_2457_),
    .B1(_2452_));
 sg13g2_xor2_1 _6364_ (.B(_2457_),
    .A(_2456_),
    .X(_2458_));
 sg13g2_nand2_1 _6365_ (.Y(_2459_),
    .A(net483),
    .B(net885));
 sg13g2_a22oi_1 _6366_ (.Y(_2460_),
    .B1(net883),
    .B2(_2458_),
    .A2(net921),
    .A1(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6367_ (.Y(_0302_),
    .A(_2459_),
    .B(_2460_));
 sg13g2_xor2_1 _6368_ (.B(\vgademo.b_cos[8] ),
    .A(net946),
    .X(_2461_));
 sg13g2_nor3_1 _6369_ (.A(_2449_),
    .B(_2451_),
    .C(_2456_),
    .Y(_2462_));
 sg13g2_o21ai_1 _6370_ (.B1(_3158_),
    .Y(_2463_),
    .A1(net954),
    .A2(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6371_ (.Y(_2464_),
    .A(_2450_),
    .B(_2463_));
 sg13g2_nor2_1 _6372_ (.A(_2462_),
    .B(_2464_),
    .Y(_2465_));
 sg13g2_nor2_1 _6373_ (.A(_2461_),
    .B(_2465_),
    .Y(_2466_));
 sg13g2_xor2_1 _6374_ (.B(_2465_),
    .A(_2461_),
    .X(_2467_));
 sg13g2_nand2_1 _6375_ (.Y(_2468_),
    .A(net438),
    .B(net885));
 sg13g2_a22oi_1 _6376_ (.Y(_2469_),
    .B1(net883),
    .B2(_2467_),
    .A2(net921),
    .A1(\vgademo.b_cos[8] ));
 sg13g2_nand2_1 _6377_ (.Y(_0303_),
    .A(_2468_),
    .B(_2469_));
 sg13g2_xnor2_1 _6378_ (.Y(_2470_),
    .A(net946),
    .B(net953));
 sg13g2_a21oi_1 _6379_ (.A1(_3158_),
    .A2(\vgademo.b_cos[8] ),
    .Y(_2471_),
    .B1(_2466_));
 sg13g2_xnor2_1 _6380_ (.Y(_2472_),
    .A(_2470_),
    .B(_2471_));
 sg13g2_nand2_1 _6381_ (.Y(_2473_),
    .A(net356),
    .B(net885));
 sg13g2_a22oi_1 _6382_ (.Y(_2474_),
    .B1(net883),
    .B2(_2472_),
    .A2(net921),
    .A1(net953));
 sg13g2_nand2_1 _6383_ (.Y(_0304_),
    .A(_2473_),
    .B(_2474_));
 sg13g2_a21oi_1 _6384_ (.A1(_3161_),
    .A2(_3162_),
    .Y(_2475_),
    .B1(net946));
 sg13g2_a21oi_1 _6385_ (.A1(_2466_),
    .A2(_2470_),
    .Y(_2476_),
    .B1(_2475_));
 sg13g2_xnor2_1 _6386_ (.Y(_2477_),
    .A(net946),
    .B(net952));
 sg13g2_nor2b_1 _6387_ (.A(_2476_),
    .B_N(_2477_),
    .Y(_2478_));
 sg13g2_xnor2_1 _6388_ (.Y(_2479_),
    .A(_2476_),
    .B(_2477_));
 sg13g2_nand2_1 _6389_ (.Y(_2480_),
    .A(net410),
    .B(net885));
 sg13g2_a22oi_1 _6390_ (.Y(_2481_),
    .B1(net883),
    .B2(_2479_),
    .A2(net921),
    .A1(net952));
 sg13g2_nand2_1 _6391_ (.Y(_0305_),
    .A(_2480_),
    .B(_2481_));
 sg13g2_a21oi_2 _6392_ (.B1(_2478_),
    .Y(_2482_),
    .A2(net952),
    .A1(_3158_));
 sg13g2_xnor2_1 _6393_ (.Y(_2483_),
    .A(net947),
    .B(\vgademo.b_cos[11] ));
 sg13g2_xnor2_1 _6394_ (.Y(_2484_),
    .A(_2482_),
    .B(_2483_));
 sg13g2_nand2_1 _6395_ (.Y(_2485_),
    .A(net464),
    .B(net885));
 sg13g2_a22oi_1 _6396_ (.Y(_2486_),
    .B1(net883),
    .B2(net841),
    .A2(net922),
    .A1(net472));
 sg13g2_nand2_1 _6397_ (.Y(_0306_),
    .A(_2485_),
    .B(_2486_));
 sg13g2_mux2_1 _6398_ (.A0(net349),
    .A1(_0226_),
    .S(_0654_),
    .X(_0307_));
 sg13g2_a21oi_1 _6399_ (.A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ),
    .Y(_2487_),
    .B1(net948));
 sg13g2_o21ai_1 _6400_ (.B1(_2487_),
    .Y(_2488_),
    .A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ));
 sg13g2_o21ai_1 _6401_ (.B1(_2488_),
    .Y(_2489_),
    .A1(_3102_),
    .A2(_0070_));
 sg13g2_nand2_1 _6402_ (.Y(_2490_),
    .A(\vgademo.plane_dx_div.r[16] ),
    .B(_2489_));
 sg13g2_xnor2_1 _6403_ (.Y(_2491_),
    .A(\vgademo.plane_dx_div.r[16] ),
    .B(_2489_));
 sg13g2_a21oi_1 _6404_ (.A1(net908),
    .A2(_2491_),
    .Y(_2492_),
    .B1(_1101_));
 sg13g2_mux2_1 _6405_ (.A0(_2492_),
    .A1(_1100_),
    .S(_1112_),
    .X(_2493_));
 sg13g2_o21ai_1 _6406_ (.B1(_2493_),
    .Y(_2494_),
    .A1(net395),
    .A2(_0654_));
 sg13g2_inv_1 _6407_ (.Y(_0308_),
    .A(_2494_));
 sg13g2_nor2_1 _6408_ (.A(net333),
    .B(_0654_),
    .Y(_2495_));
 sg13g2_o21ai_1 _6409_ (.B1(\vgademo.plane_dx_div.d[18] ),
    .Y(_2496_),
    .A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ));
 sg13g2_or3_2 _6410_ (.A(\vgademo.plane_dx_div.d[16] ),
    .B(\vgademo.plane_dx_div.d[17] ),
    .C(\vgademo.plane_dx_div.d[18] ),
    .X(_2497_));
 sg13g2_a21oi_1 _6411_ (.A1(_2496_),
    .A2(_2497_),
    .Y(_2498_),
    .B1(net948));
 sg13g2_a21oi_1 _6412_ (.A1(net948),
    .A2(_0073_),
    .Y(_2499_),
    .B1(_2498_));
 sg13g2_nand2_1 _6413_ (.Y(_2500_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2499_));
 sg13g2_xnor2_1 _6414_ (.Y(_2501_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2499_));
 sg13g2_xnor2_1 _6415_ (.Y(_2502_),
    .A(_2490_),
    .B(_2501_));
 sg13g2_nand2_1 _6416_ (.Y(_2503_),
    .A(_1100_),
    .B(_1111_));
 sg13g2_nand2b_1 _6417_ (.Y(_2504_),
    .B(_2503_),
    .A_N(_1125_));
 sg13g2_xor2_1 _6418_ (.B(_2503_),
    .A(_1125_),
    .X(_2505_));
 sg13g2_a221oi_1 _6419_ (.B2(_0650_),
    .C1(_2495_),
    .B1(_2505_),
    .A1(net908),
    .Y(_0309_),
    .A2(_2502_));
 sg13g2_nor2_1 _6420_ (.A(net340),
    .B(_0654_),
    .Y(_2506_));
 sg13g2_a21oi_1 _6421_ (.A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2497_),
    .Y(_2507_),
    .B1(net948));
 sg13g2_o21ai_1 _6422_ (.B1(_2507_),
    .Y(_2508_),
    .A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2497_));
 sg13g2_o21ai_1 _6423_ (.B1(_2508_),
    .Y(_2509_),
    .A1(_3102_),
    .A2(_0076_));
 sg13g2_and2_1 _6424_ (.A(\vgademo.plane_dx_div.r[18] ),
    .B(_2509_),
    .X(_2510_));
 sg13g2_xor2_1 _6425_ (.B(_2509_),
    .A(\vgademo.plane_dx_div.r[18] ),
    .X(_2511_));
 sg13g2_o21ai_1 _6426_ (.B1(_2500_),
    .Y(_2512_),
    .A1(_2490_),
    .A2(_2501_));
 sg13g2_xnor2_1 _6427_ (.Y(_2513_),
    .A(_2511_),
    .B(_2512_));
 sg13g2_nand2b_1 _6428_ (.Y(_2514_),
    .B(_1140_),
    .A_N(_2504_));
 sg13g2_xor2_1 _6429_ (.B(_2504_),
    .A(_1140_),
    .X(_2515_));
 sg13g2_a221oi_1 _6430_ (.B2(_0650_),
    .C1(_2506_),
    .B1(_2515_),
    .A1(net908),
    .Y(_0310_),
    .A2(_2513_));
 sg13g2_nor2_1 _6431_ (.A(net277),
    .B(_0654_),
    .Y(_2516_));
 sg13g2_o21ai_1 _6432_ (.B1(\vgademo.plane_dx_div.d[20] ),
    .Y(_2517_),
    .A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2497_));
 sg13g2_or3_2 _6433_ (.A(\vgademo.plane_dx_div.d[19] ),
    .B(\vgademo.plane_dx_div.d[20] ),
    .C(_2497_),
    .X(_2518_));
 sg13g2_a21oi_1 _6434_ (.A1(_2517_),
    .A2(_2518_),
    .Y(_2519_),
    .B1(net948));
 sg13g2_a21oi_1 _6435_ (.A1(net948),
    .A2(_0079_),
    .Y(_2520_),
    .B1(_2519_));
 sg13g2_nand2_1 _6436_ (.Y(_2521_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .B(_2520_));
 sg13g2_xnor2_1 _6437_ (.Y(_2522_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .B(_2520_));
 sg13g2_a21oi_1 _6438_ (.A1(_2511_),
    .A2(_2512_),
    .Y(_2523_),
    .B1(_2510_));
 sg13g2_xnor2_1 _6439_ (.Y(_2524_),
    .A(_2522_),
    .B(_2523_));
 sg13g2_nor2_1 _6440_ (.A(_1155_),
    .B(_2514_),
    .Y(_2525_));
 sg13g2_xnor2_1 _6441_ (.Y(_2526_),
    .A(_1155_),
    .B(_2514_));
 sg13g2_a221oi_1 _6442_ (.B2(net929),
    .C1(_2516_),
    .B1(_2526_),
    .A1(net908),
    .Y(_0311_),
    .A2(_2524_));
 sg13g2_nor2_1 _6443_ (.A(net313),
    .B(_0654_),
    .Y(_2527_));
 sg13g2_xor2_1 _6444_ (.B(_2518_),
    .A(\vgademo.plane_dx_div.d[21] ),
    .X(_2528_));
 sg13g2_nor2_1 _6445_ (.A(net949),
    .B(_2528_),
    .Y(_2529_));
 sg13g2_and2_1 _6446_ (.A(net949),
    .B(_0081_),
    .X(_2530_));
 sg13g2_nor3_1 _6447_ (.A(_3141_),
    .B(_2529_),
    .C(_2530_),
    .Y(_2531_));
 sg13g2_o21ai_1 _6448_ (.B1(_3141_),
    .Y(_2532_),
    .A1(_2529_),
    .A2(_2530_));
 sg13g2_nor2b_1 _6449_ (.A(_2531_),
    .B_N(_2532_),
    .Y(_2533_));
 sg13g2_o21ai_1 _6450_ (.B1(_2521_),
    .Y(_2534_),
    .A1(_2522_),
    .A2(_2523_));
 sg13g2_xnor2_1 _6451_ (.Y(_2535_),
    .A(_2533_),
    .B(_2534_));
 sg13g2_nand2_1 _6452_ (.Y(_2536_),
    .A(_1173_),
    .B(_2525_));
 sg13g2_xnor2_1 _6453_ (.Y(_2537_),
    .A(_1173_),
    .B(_2525_));
 sg13g2_a221oi_1 _6454_ (.B2(net929),
    .C1(_2527_),
    .B1(_2537_),
    .A1(net908),
    .Y(_0312_),
    .A2(_2535_));
 sg13g2_nand2b_1 _6455_ (.Y(_2538_),
    .B(_1191_),
    .A_N(_2536_));
 sg13g2_xor2_1 _6456_ (.B(_2536_),
    .A(_1191_),
    .X(_2539_));
 sg13g2_a21oi_1 _6457_ (.A1(_2532_),
    .A2(_2534_),
    .Y(_2540_),
    .B1(_2531_));
 sg13g2_nand2b_1 _6458_ (.Y(_2541_),
    .B(net948),
    .A_N(_0013_));
 sg13g2_o21ai_1 _6459_ (.B1(\vgademo.plane_dx_div.d[22] ),
    .Y(_2542_),
    .A1(\vgademo.plane_dx_div.d[21] ),
    .A2(_2518_));
 sg13g2_nor3_1 _6460_ (.A(\vgademo.plane_dx_div.d[21] ),
    .B(\vgademo.plane_dx_div.d[22] ),
    .C(_2518_),
    .Y(_2543_));
 sg13g2_nand2_1 _6461_ (.Y(_2544_),
    .A(_3102_),
    .B(_2542_));
 sg13g2_o21ai_1 _6462_ (.B1(_2541_),
    .Y(_2545_),
    .A1(_2543_),
    .A2(_2544_));
 sg13g2_or2_1 _6463_ (.X(_2546_),
    .B(_2545_),
    .A(\vgademo.plane_dx_div.r[21] ));
 sg13g2_nand2_1 _6464_ (.Y(_2547_),
    .A(net313),
    .B(_2545_));
 sg13g2_nand2_1 _6465_ (.Y(_2548_),
    .A(_2546_),
    .B(_2547_));
 sg13g2_nand2_1 _6466_ (.Y(_2549_),
    .A(_2540_),
    .B(_2547_));
 sg13g2_xnor2_1 _6467_ (.Y(_2550_),
    .A(_2540_),
    .B(_2548_));
 sg13g2_nor2_1 _6468_ (.A(net351),
    .B(_0654_),
    .Y(_2551_));
 sg13g2_a221oi_1 _6469_ (.B2(net908),
    .C1(_2551_),
    .B1(_2550_),
    .A1(net929),
    .Y(_0313_),
    .A2(_2539_));
 sg13g2_nand2b_1 _6470_ (.Y(_2552_),
    .B(\vgademo.plane_dx_div.d[23] ),
    .A_N(_2543_));
 sg13g2_nand2b_1 _6471_ (.Y(_2553_),
    .B(_2543_),
    .A_N(\vgademo.plane_dx_div.d[23] ));
 sg13g2_nand3_1 _6472_ (.B(_2552_),
    .C(_2553_),
    .A(_3102_),
    .Y(_2554_));
 sg13g2_o21ai_1 _6473_ (.B1(_2554_),
    .Y(_2555_),
    .A1(_3102_),
    .A2(_0017_));
 sg13g2_and2_1 _6474_ (.A(\vgademo.plane_dx_div.r[22] ),
    .B(_2555_),
    .X(_2556_));
 sg13g2_xor2_1 _6475_ (.B(_2555_),
    .A(\vgademo.plane_dx_div.r[22] ),
    .X(_2557_));
 sg13g2_a21oi_1 _6476_ (.A1(_2546_),
    .A2(_2549_),
    .Y(_2558_),
    .B1(_2557_));
 sg13g2_and3_1 _6477_ (.X(_2559_),
    .A(_2546_),
    .B(_2549_),
    .C(_2557_));
 sg13g2_nor2_1 _6478_ (.A(_2558_),
    .B(_2559_),
    .Y(_2560_));
 sg13g2_nand2_1 _6479_ (.Y(_2561_),
    .A(_1207_),
    .B(_2538_));
 sg13g2_nor2_1 _6480_ (.A(_1207_),
    .B(_2538_),
    .Y(_2562_));
 sg13g2_nor2_1 _6481_ (.A(net926),
    .B(_2562_),
    .Y(_2563_));
 sg13g2_a221oi_1 _6482_ (.B2(_2563_),
    .C1(net905),
    .B1(_2561_),
    .A1(net926),
    .Y(_2564_),
    .A2(_2560_));
 sg13g2_a21oi_1 _6483_ (.A1(_3144_),
    .A2(net905),
    .Y(_0314_),
    .B1(_2564_));
 sg13g2_nand2_1 _6484_ (.Y(_2565_),
    .A(\vgademo.plane_dx_div.d[24] ),
    .B(_2553_));
 sg13g2_nor2_1 _6485_ (.A(\vgademo.plane_dx_div.d[24] ),
    .B(_2553_),
    .Y(_2566_));
 sg13g2_nor2_1 _6486_ (.A(net949),
    .B(_2566_),
    .Y(_2567_));
 sg13g2_a22oi_1 _6487_ (.Y(_2568_),
    .B1(_2565_),
    .B2(_2567_),
    .A2(_3143_),
    .A1(net949));
 sg13g2_xnor2_1 _6488_ (.Y(_2569_),
    .A(\vgademo.plane_dx_div.r[23] ),
    .B(_2568_));
 sg13g2_nor3_1 _6489_ (.A(_2556_),
    .B(_2559_),
    .C(_2569_),
    .Y(_2570_));
 sg13g2_o21ai_1 _6490_ (.B1(_2569_),
    .Y(_2571_),
    .A1(_2556_),
    .A2(_2559_));
 sg13g2_nor2_1 _6491_ (.A(net927),
    .B(_2570_),
    .Y(_2572_));
 sg13g2_a21oi_1 _6492_ (.A1(_2571_),
    .A2(_2572_),
    .Y(_2573_),
    .B1(net905));
 sg13g2_o21ai_1 _6493_ (.B1(_1216_),
    .Y(_2574_),
    .A1(_1207_),
    .A2(_2538_));
 sg13g2_nor2_1 _6494_ (.A(_1217_),
    .B(_2563_),
    .Y(_2575_));
 sg13g2_o21ai_1 _6495_ (.B1(_2574_),
    .Y(_2576_),
    .A1(_1217_),
    .A2(_2563_));
 sg13g2_a22oi_1 _6496_ (.Y(_0315_),
    .B1(_2573_),
    .B2(_2576_),
    .A2(net905),
    .A1(_3145_));
 sg13g2_o21ai_1 _6497_ (.B1(_2571_),
    .Y(_2577_),
    .A1(_3144_),
    .A2(_2568_));
 sg13g2_xnor2_1 _6498_ (.Y(_2578_),
    .A(\vgademo.plane_dx_div.r[24] ),
    .B(_2567_));
 sg13g2_xnor2_1 _6499_ (.Y(_2579_),
    .A(_2577_),
    .B(_2578_));
 sg13g2_a21oi_1 _6500_ (.A1(net926),
    .A2(_2579_),
    .Y(_2580_),
    .B1(net905));
 sg13g2_a22oi_1 _6501_ (.Y(_0316_),
    .B1(_2575_),
    .B2(_2580_),
    .A2(net905),
    .A1(_3102_));
 sg13g2_and2_1 _6502_ (.A(_2150_),
    .B(_2159_),
    .X(_2581_));
 sg13g2_inv_1 _6503_ (.Y(_2582_),
    .A(_2581_));
 sg13g2_and2_1 _6504_ (.A(_2183_),
    .B(_2582_),
    .X(_2583_));
 sg13g2_o21ai_1 _6505_ (.B1(_1870_),
    .Y(_2584_),
    .A1(_1818_),
    .A2(_1828_));
 sg13g2_and2_1 _6506_ (.A(net847),
    .B(_2584_),
    .X(_2585_));
 sg13g2_a221oi_1 _6507_ (.B2(net810),
    .C1(_1761_),
    .B1(_2585_),
    .A1(_1354_),
    .Y(_2586_),
    .A2(_2143_));
 sg13g2_nor2_1 _6508_ (.A(_2583_),
    .B(_2586_),
    .Y(_2587_));
 sg13g2_o21ai_1 _6509_ (.B1(net858),
    .Y(_2588_),
    .A1(_2583_),
    .A2(_2586_));
 sg13g2_and2_1 _6510_ (.A(_1331_),
    .B(_2588_),
    .X(_2589_));
 sg13g2_a21oi_2 _6511_ (.B1(_2167_),
    .Y(_2590_),
    .A2(_1869_),
    .A1(_1823_));
 sg13g2_o21ai_1 _6512_ (.B1(net847),
    .Y(_2591_),
    .A1(_1785_),
    .A2(_2590_));
 sg13g2_a221oi_1 _6513_ (.B2(_2173_),
    .C1(_2161_),
    .B1(_2591_),
    .A1(_2183_),
    .Y(_2592_),
    .A2(_2582_));
 sg13g2_nand2_1 _6514_ (.Y(_2593_),
    .A(_2178_),
    .B(_2592_));
 sg13g2_nand2_1 _6515_ (.Y(_2594_),
    .A(_2589_),
    .B(_2593_));
 sg13g2_nor2_1 _6516_ (.A(_2178_),
    .B(_2592_),
    .Y(_2595_));
 sg13g2_nor2_1 _6517_ (.A(_2589_),
    .B(_2595_),
    .Y(_2596_));
 sg13g2_a21oi_1 _6518_ (.A1(_2589_),
    .A2(_2593_),
    .Y(_2597_),
    .B1(_2596_));
 sg13g2_nor2b_1 _6519_ (.A(_2193_),
    .B_N(_2166_),
    .Y(_2598_));
 sg13g2_nor4_1 _6520_ (.A(net814),
    .B(net812),
    .C(net852),
    .D(_2584_),
    .Y(_2599_));
 sg13g2_a221oi_1 _6521_ (.B2(_2598_),
    .C1(_2599_),
    .B1(net810),
    .A1(net855),
    .Y(_2600_),
    .A2(net853));
 sg13g2_o21ai_1 _6522_ (.B1(_1762_),
    .Y(_2601_),
    .A1(_2198_),
    .A2(_2600_));
 sg13g2_nand2_2 _6523_ (.Y(_2602_),
    .A(_2185_),
    .B(_2601_));
 sg13g2_nand2b_1 _6524_ (.Y(_2603_),
    .B(_2602_),
    .A_N(net936));
 sg13g2_xor2_1 _6525_ (.B(_2602_),
    .A(net936),
    .X(_2604_));
 sg13g2_o21ai_1 _6526_ (.B1(_2603_),
    .Y(_2605_),
    .A1(_2592_),
    .A2(_2604_));
 sg13g2_xnor2_1 _6527_ (.Y(_2606_),
    .A(_2178_),
    .B(_2592_));
 sg13g2_xnor2_1 _6528_ (.Y(_2607_),
    .A(_2589_),
    .B(_2606_));
 sg13g2_or2_1 _6529_ (.X(_2608_),
    .B(_2607_),
    .A(_2605_));
 sg13g2_nor2_1 _6530_ (.A(_2192_),
    .B(_2216_),
    .Y(_2609_));
 sg13g2_nor4_1 _6531_ (.A(net814),
    .B(net812),
    .C(net852),
    .D(_2609_),
    .Y(_2610_));
 sg13g2_nand2_1 _6532_ (.Y(_2611_),
    .A(_2227_),
    .B(_2237_));
 sg13g2_a221oi_1 _6533_ (.B2(_2611_),
    .C1(_2610_),
    .B1(net811),
    .A1(net855),
    .Y(_2612_),
    .A2(net853));
 sg13g2_o21ai_1 _6534_ (.B1(_1329_),
    .Y(_2613_),
    .A1(_2171_),
    .A2(_2612_));
 sg13g2_nand2_1 _6535_ (.Y(_2614_),
    .A(net935),
    .B(_2613_));
 sg13g2_and2_1 _6536_ (.A(_2215_),
    .B(_2228_),
    .X(_2615_));
 sg13g2_mux2_1 _6537_ (.A0(_2598_),
    .A1(_2615_),
    .S(net810),
    .X(_2616_));
 sg13g2_a21oi_1 _6538_ (.A1(net847),
    .A2(_2616_),
    .Y(_2617_),
    .B1(_2222_));
 sg13g2_nor2_2 _6539_ (.A(_1328_),
    .B(_2617_),
    .Y(_2618_));
 sg13g2_nor2_1 _6540_ (.A(net935),
    .B(_2613_),
    .Y(_2619_));
 sg13g2_xor2_1 _6541_ (.B(_2613_),
    .A(net935),
    .X(_2620_));
 sg13g2_o21ai_1 _6542_ (.B1(_2614_),
    .Y(_2621_),
    .A1(_2618_),
    .A2(_2619_));
 sg13g2_mux2_1 _6543_ (.A0(_2590_),
    .A1(_2609_),
    .S(net810),
    .X(_2622_));
 sg13g2_a21oi_2 _6544_ (.B1(_2210_),
    .Y(_2623_),
    .A2(_2622_),
    .A1(net847));
 sg13g2_and2_1 _6545_ (.A(_2183_),
    .B(_2581_),
    .X(_2624_));
 sg13g2_a21o_1 _6546_ (.A2(_2161_),
    .A1(_2151_),
    .B1(_2624_),
    .X(_2625_));
 sg13g2_or2_1 _6547_ (.X(_2626_),
    .B(_2625_),
    .A(_2623_));
 sg13g2_o21ai_1 _6548_ (.B1(_2251_),
    .Y(_2627_),
    .A1(_2623_),
    .A2(_2625_));
 sg13g2_or3_1 _6549_ (.A(_2251_),
    .B(_2623_),
    .C(_2625_),
    .X(_2628_));
 sg13g2_nand3_1 _6550_ (.B(_2627_),
    .C(_2628_),
    .A(_2602_),
    .Y(_2629_));
 sg13g2_a21o_1 _6551_ (.A2(_2628_),
    .A1(_2627_),
    .B1(_2602_),
    .X(_2630_));
 sg13g2_and2_1 _6552_ (.A(_2629_),
    .B(_2630_),
    .X(_2631_));
 sg13g2_nand2_1 _6553_ (.Y(_2632_),
    .A(_2232_),
    .B(_2587_));
 sg13g2_a21oi_1 _6554_ (.A1(_1331_),
    .A2(_2588_),
    .Y(_2633_),
    .B1(_2232_));
 sg13g2_o21ai_1 _6555_ (.B1(_2632_),
    .Y(_2634_),
    .A1(_2618_),
    .A2(_2633_));
 sg13g2_or2_1 _6556_ (.X(_2635_),
    .B(_2634_),
    .A(_2626_));
 sg13g2_xnor2_1 _6557_ (.Y(_2636_),
    .A(_2618_),
    .B(_2620_));
 sg13g2_a21o_1 _6558_ (.A2(_2634_),
    .A1(_2626_),
    .B1(_2636_),
    .X(_2637_));
 sg13g2_a22oi_1 _6559_ (.Y(_2638_),
    .B1(_2635_),
    .B2(_2637_),
    .A2(_2631_),
    .A1(_2621_));
 sg13g2_xor2_1 _6560_ (.B(_2604_),
    .A(_2592_),
    .X(_2639_));
 sg13g2_xnor2_1 _6561_ (.Y(_2640_),
    .A(_2592_),
    .B(_2604_));
 sg13g2_and2_1 _6562_ (.A(_2627_),
    .B(_2629_),
    .X(_2641_));
 sg13g2_nand2_1 _6563_ (.Y(_2642_),
    .A(_2627_),
    .B(_2629_));
 sg13g2_a21oi_1 _6564_ (.A1(_2629_),
    .A2(_2630_),
    .Y(_2643_),
    .B1(_2621_));
 sg13g2_a21o_1 _6565_ (.A2(_2641_),
    .A1(_2640_),
    .B1(_2643_),
    .X(_2644_));
 sg13g2_a22oi_1 _6566_ (.Y(_2645_),
    .B1(_2639_),
    .B2(_2642_),
    .A2(_2607_),
    .A1(_2605_));
 sg13g2_o21ai_1 _6567_ (.B1(_2645_),
    .Y(_2646_),
    .A1(_2638_),
    .A2(_2644_));
 sg13g2_a21oi_1 _6568_ (.A1(_2608_),
    .A2(_2646_),
    .Y(_2647_),
    .B1(_2597_));
 sg13g2_and3_1 _6569_ (.X(_2648_),
    .A(_2597_),
    .B(_2608_),
    .C(_2646_));
 sg13g2_nand3_1 _6570_ (.B(_2608_),
    .C(_2646_),
    .A(_2597_),
    .Y(_2649_));
 sg13g2_nor3_1 _6571_ (.A(_2270_),
    .B(_2647_),
    .C(_2648_),
    .Y(_0317_));
 sg13g2_a21oi_1 _6572_ (.A1(_2594_),
    .A2(_2649_),
    .Y(_0318_),
    .B1(_2270_));
 sg13g2_nand2_1 _6573_ (.Y(_2650_),
    .A(\vgademo.b_sin[0] ),
    .B(_2458_));
 sg13g2_xnor2_1 _6574_ (.Y(_2651_),
    .A(net414),
    .B(_2458_));
 sg13g2_a22oi_1 _6575_ (.Y(_2652_),
    .B1(net886),
    .B2(net385),
    .A2(net921),
    .A1(net414));
 sg13g2_o21ai_1 _6576_ (.B1(_2652_),
    .Y(_0319_),
    .A1(net882),
    .A2(_2651_));
 sg13g2_xnor2_1 _6577_ (.Y(_2653_),
    .A(net378),
    .B(_2467_));
 sg13g2_or2_1 _6578_ (.X(_2654_),
    .B(_2653_),
    .A(_2650_));
 sg13g2_inv_1 _6579_ (.Y(_2655_),
    .A(_2654_));
 sg13g2_a21o_1 _6580_ (.A2(_2653_),
    .A1(_2650_),
    .B1(net882),
    .X(_2656_));
 sg13g2_a22oi_1 _6581_ (.Y(_2657_),
    .B1(net885),
    .B2(net366),
    .A2(net921),
    .A1(net378));
 sg13g2_o21ai_1 _6582_ (.B1(_2657_),
    .Y(_0320_),
    .A1(_2655_),
    .A2(_2656_));
 sg13g2_a21oi_1 _6583_ (.A1(net378),
    .A2(_2467_),
    .Y(_2658_),
    .B1(_2655_));
 sg13g2_xnor2_1 _6584_ (.Y(_2659_),
    .A(net380),
    .B(_2472_));
 sg13g2_nor2_1 _6585_ (.A(_2658_),
    .B(_2659_),
    .Y(_2660_));
 sg13g2_a21o_1 _6586_ (.A2(_2659_),
    .A1(_2658_),
    .B1(net882),
    .X(_2661_));
 sg13g2_a22oi_1 _6587_ (.Y(_2662_),
    .B1(net885),
    .B2(net365),
    .A2(net921),
    .A1(net380));
 sg13g2_o21ai_1 _6588_ (.B1(_2662_),
    .Y(_0321_),
    .A1(_2660_),
    .A2(_2661_));
 sg13g2_a21oi_1 _6589_ (.A1(\vgademo.b_sin[2] ),
    .A2(_2472_),
    .Y(_2663_),
    .B1(_2660_));
 sg13g2_nand2_1 _6590_ (.Y(_2664_),
    .A(net405),
    .B(_2479_));
 sg13g2_xnor2_1 _6591_ (.Y(_2665_),
    .A(net405),
    .B(_2479_));
 sg13g2_or2_1 _6592_ (.X(_2666_),
    .B(_2665_),
    .A(_2663_));
 sg13g2_a21oi_1 _6593_ (.A1(_2663_),
    .A2(_2665_),
    .Y(_2667_),
    .B1(net882));
 sg13g2_nand2_1 _6594_ (.Y(_2668_),
    .A(_2666_),
    .B(_2667_));
 sg13g2_a22oi_1 _6595_ (.Y(_2669_),
    .B1(net886),
    .B2(\vgademo.a_sin[6] ),
    .A2(net922),
    .A1(net405));
 sg13g2_nand2_1 _6596_ (.Y(_0322_),
    .A(_2668_),
    .B(net406));
 sg13g2_nand2_1 _6597_ (.Y(_2670_),
    .A(\vgademo.b_sin[4] ),
    .B(net839));
 sg13g2_xnor2_1 _6598_ (.Y(_2671_),
    .A(\vgademo.b_sin[4] ),
    .B(net841));
 sg13g2_a21o_1 _6599_ (.A2(_2666_),
    .A1(_2664_),
    .B1(_2671_),
    .X(_2672_));
 sg13g2_nand3_1 _6600_ (.B(_2666_),
    .C(_2671_),
    .A(_2664_),
    .Y(_2673_));
 sg13g2_nand3_1 _6601_ (.B(_2672_),
    .C(_2673_),
    .A(net883),
    .Y(_2674_));
 sg13g2_a22oi_1 _6602_ (.Y(_2675_),
    .B1(net886),
    .B2(net448),
    .A2(net923),
    .A1(\vgademo.b_sin[4] ));
 sg13g2_nand2_1 _6603_ (.Y(_0323_),
    .A(_2674_),
    .B(net449));
 sg13g2_nand2_1 _6604_ (.Y(_2676_),
    .A(net298),
    .B(net924));
 sg13g2_xor2_1 _6605_ (.B(net840),
    .A(net298),
    .X(_2677_));
 sg13g2_and2_1 _6606_ (.A(_2670_),
    .B(_2672_),
    .X(_2678_));
 sg13g2_o21ai_1 _6607_ (.B1(net894),
    .Y(_2679_),
    .A1(_2677_),
    .A2(_2678_));
 sg13g2_a21oi_1 _6608_ (.A1(_2677_),
    .A2(_2678_),
    .Y(_2680_),
    .B1(_2679_));
 sg13g2_o21ai_1 _6609_ (.B1(net925),
    .Y(_2681_),
    .A1(\vgademo.a_sin[8] ),
    .A2(net894));
 sg13g2_o21ai_1 _6610_ (.B1(_2676_),
    .Y(_0324_),
    .A1(_2680_),
    .A2(_2681_));
 sg13g2_xnor2_1 _6611_ (.Y(_2682_),
    .A(\vgademo.b_sin[6] ),
    .B(net840));
 sg13g2_o21ai_1 _6612_ (.B1(net840),
    .Y(_2683_),
    .A1(\vgademo.b_sin[4] ),
    .A2(\vgademo.b_sin[5] ));
 sg13g2_nor2b_1 _6613_ (.A(_2672_),
    .B_N(_2677_),
    .Y(_2684_));
 sg13g2_nor2b_1 _6614_ (.A(_2684_),
    .B_N(_2683_),
    .Y(_2685_));
 sg13g2_nor2_1 _6615_ (.A(_2682_),
    .B(_2685_),
    .Y(_2686_));
 sg13g2_a21o_1 _6616_ (.A2(_2685_),
    .A1(_2682_),
    .B1(net882),
    .X(_2687_));
 sg13g2_a22oi_1 _6617_ (.Y(_2688_),
    .B1(net886),
    .B2(\vgademo.a_sin[9] ),
    .A2(net923),
    .A1(net418));
 sg13g2_o21ai_1 _6618_ (.B1(net419),
    .Y(_0325_),
    .A1(_2686_),
    .A2(_2687_));
 sg13g2_nand2_1 _6619_ (.Y(_2689_),
    .A(net358),
    .B(net923));
 sg13g2_xnor2_1 _6620_ (.Y(_2690_),
    .A(\vgademo.b_sin[7] ),
    .B(net840));
 sg13g2_a21oi_1 _6621_ (.A1(\vgademo.b_sin[6] ),
    .A2(net839),
    .Y(_2691_),
    .B1(_2686_));
 sg13g2_inv_1 _6622_ (.Y(_2692_),
    .A(_2691_));
 sg13g2_o21ai_1 _6623_ (.B1(net894),
    .Y(_2693_),
    .A1(_2690_),
    .A2(_2692_));
 sg13g2_a21oi_1 _6624_ (.A1(_2690_),
    .A2(_2692_),
    .Y(_2694_),
    .B1(_2693_));
 sg13g2_o21ai_1 _6625_ (.B1(net925),
    .Y(_2695_),
    .A1(\vgademo.a_sin[10] ),
    .A2(net894));
 sg13g2_o21ai_1 _6626_ (.B1(_2689_),
    .Y(_0326_),
    .A1(_2694_),
    .A2(_2695_));
 sg13g2_nand2_1 _6627_ (.Y(_2696_),
    .A(\vgademo.b_sin[8] ),
    .B(net839));
 sg13g2_xnor2_1 _6628_ (.Y(_2697_),
    .A(\vgademo.b_sin[8] ),
    .B(net839));
 sg13g2_nor2_1 _6629_ (.A(_2682_),
    .B(_2690_),
    .Y(_2698_));
 sg13g2_o21ai_1 _6630_ (.B1(net839),
    .Y(_2699_),
    .A1(\vgademo.b_sin[7] ),
    .A2(\vgademo.b_sin[6] ));
 sg13g2_nand2_1 _6631_ (.Y(_2700_),
    .A(_2683_),
    .B(_2699_));
 sg13g2_a21oi_1 _6632_ (.A1(_2684_),
    .A2(_2698_),
    .Y(_2701_),
    .B1(_2700_));
 sg13g2_or2_1 _6633_ (.X(_2702_),
    .B(_2701_),
    .A(_2697_));
 sg13g2_a21oi_1 _6634_ (.A1(_2697_),
    .A2(_2701_),
    .Y(_2703_),
    .B1(net882));
 sg13g2_nand2_1 _6635_ (.Y(_2704_),
    .A(_2702_),
    .B(_2703_));
 sg13g2_a22oi_1 _6636_ (.Y(_2705_),
    .B1(net886),
    .B2(net488),
    .A2(net923),
    .A1(net489));
 sg13g2_nand2_1 _6637_ (.Y(_0327_),
    .A(_2704_),
    .B(_2705_));
 sg13g2_nand2_1 _6638_ (.Y(_2706_),
    .A(net436),
    .B(net923));
 sg13g2_o21ai_1 _6639_ (.B1(net925),
    .Y(_2707_),
    .A1(\vgademo.a_sin[12] ),
    .A2(net893));
 sg13g2_nand2_1 _6640_ (.Y(_2708_),
    .A(_2696_),
    .B(_2702_));
 sg13g2_xnor2_1 _6641_ (.Y(_2709_),
    .A(\vgademo.b_sin[9] ),
    .B(net839));
 sg13g2_o21ai_1 _6642_ (.B1(net893),
    .Y(_2710_),
    .A1(_2708_),
    .A2(_2709_));
 sg13g2_a21oi_1 _6643_ (.A1(_2708_),
    .A2(_2709_),
    .Y(_2711_),
    .B1(_2710_));
 sg13g2_o21ai_1 _6644_ (.B1(_2706_),
    .Y(_0328_),
    .A1(_2707_),
    .A2(_2711_));
 sg13g2_nand2_1 _6645_ (.Y(_2712_),
    .A(\vgademo.b_sin[10] ),
    .B(net841));
 sg13g2_xnor2_1 _6646_ (.Y(_2713_),
    .A(\vgademo.b_sin[10] ),
    .B(net841));
 sg13g2_a21o_1 _6647_ (.A2(net839),
    .A1(\vgademo.b_sin[9] ),
    .B1(_2708_),
    .X(_2714_));
 sg13g2_o21ai_1 _6648_ (.B1(_2714_),
    .Y(_2715_),
    .A1(\vgademo.b_sin[9] ),
    .A2(net839));
 sg13g2_or2_1 _6649_ (.X(_2716_),
    .B(_2715_),
    .A(_2713_));
 sg13g2_a21oi_1 _6650_ (.A1(_2713_),
    .A2(_2715_),
    .Y(_2717_),
    .B1(net882));
 sg13g2_nand2_1 _6651_ (.Y(_2718_),
    .A(_2716_),
    .B(_2717_));
 sg13g2_a22oi_1 _6652_ (.Y(_2719_),
    .B1(net887),
    .B2(net467),
    .A2(net923),
    .A1(\vgademo.b_sin[10] ));
 sg13g2_nand2_1 _6653_ (.Y(_0329_),
    .A(_2718_),
    .B(net468));
 sg13g2_nand2_1 _6654_ (.Y(_2720_),
    .A(net946),
    .B(net922));
 sg13g2_nand2_1 _6655_ (.Y(_2721_),
    .A(_2712_),
    .B(_2716_));
 sg13g2_xnor2_1 _6656_ (.Y(_2722_),
    .A(\vgademo.b_cos[11] ),
    .B(_2482_));
 sg13g2_o21ai_1 _6657_ (.B1(net893),
    .Y(_2723_),
    .A1(_2721_),
    .A2(_2722_));
 sg13g2_a21oi_1 _6658_ (.A1(_2721_),
    .A2(_2722_),
    .Y(_2724_),
    .B1(_2723_));
 sg13g2_o21ai_1 _6659_ (.B1(net925),
    .Y(_2725_),
    .A1(\vgademo.a_sin[14] ),
    .A2(net893));
 sg13g2_o21ai_1 _6660_ (.B1(_2720_),
    .Y(_0330_),
    .A1(_2724_),
    .A2(_2725_));
 sg13g2_o21ai_1 _6661_ (.B1(net1067),
    .Y(_2726_),
    .A1(net901),
    .A2(_2266_));
 sg13g2_inv_1 _6662_ (.Y(_2727_),
    .A(net876));
 sg13g2_nand2_1 _6663_ (.Y(_2728_),
    .A(net219),
    .B(\vgademo.plane_du[0] ));
 sg13g2_nand2_1 _6664_ (.Y(_2729_),
    .A(net283),
    .B(net310));
 sg13g2_xor2_1 _6665_ (.B(\vgademo.plane_du[1] ),
    .A(\vgademo.plane_u[1] ),
    .X(_2730_));
 sg13g2_nand2b_1 _6666_ (.Y(_2731_),
    .B(_2730_),
    .A_N(_2728_));
 sg13g2_xor2_1 _6667_ (.B(_2730_),
    .A(_2728_),
    .X(_2732_));
 sg13g2_nor2_1 _6668_ (.A(net900),
    .B(_2732_),
    .Y(_2733_));
 sg13g2_a21oi_1 _6669_ (.A1(\vgademo.plane_dx[0] ),
    .A2(net899),
    .Y(_2734_),
    .B1(_2733_));
 sg13g2_nand2_1 _6670_ (.Y(_2735_),
    .A(net283),
    .B(net880));
 sg13g2_o21ai_1 _6671_ (.B1(_2735_),
    .Y(_0331_),
    .A1(net880),
    .A2(_2734_));
 sg13g2_nand2_1 _6672_ (.Y(_2736_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_xnor2_1 _6673_ (.Y(_2737_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_nand3_1 _6674_ (.B(_2731_),
    .C(_2737_),
    .A(_2729_),
    .Y(_2738_));
 sg13g2_a21o_1 _6675_ (.A2(_2731_),
    .A1(_2729_),
    .B1(_2737_),
    .X(_2739_));
 sg13g2_nand3_1 _6676_ (.B(_2738_),
    .C(_2739_),
    .A(net895),
    .Y(_2740_));
 sg13g2_nand2_1 _6677_ (.Y(_2741_),
    .A(_3098_),
    .B(net950));
 sg13g2_xnor2_1 _6678_ (.Y(_2742_),
    .A(\vgademo.plane_dx[1] ),
    .B(net950));
 sg13g2_a21oi_1 _6679_ (.A1(net899),
    .A2(_2742_),
    .Y(_2743_),
    .B1(net880));
 sg13g2_a22oi_1 _6680_ (.Y(_0332_),
    .B1(_2740_),
    .B2(_2743_),
    .A2(net876),
    .A1(_3172_));
 sg13g2_nand2_1 _6681_ (.Y(_2744_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_xnor2_1 _6682_ (.Y(_2745_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_nand3_1 _6683_ (.B(_2739_),
    .C(_2745_),
    .A(_2736_),
    .Y(_2746_));
 sg13g2_a21o_1 _6684_ (.A2(_2739_),
    .A1(_2736_),
    .B1(_2745_),
    .X(_2747_));
 sg13g2_nor2_1 _6685_ (.A(\vgademo.plane_dx[2] ),
    .B(_2741_),
    .Y(_2748_));
 sg13g2_xnor2_1 _6686_ (.Y(_2749_),
    .A(\vgademo.plane_dx[2] ),
    .B(_2741_));
 sg13g2_a21oi_1 _6687_ (.A1(_2746_),
    .A2(_2747_),
    .Y(_2750_),
    .B1(net901));
 sg13g2_a21oi_1 _6688_ (.A1(net899),
    .A2(_2749_),
    .Y(_2751_),
    .B1(_2750_));
 sg13g2_mux2_1 _6689_ (.A0(net377),
    .A1(_2751_),
    .S(_2727_),
    .X(_0333_));
 sg13g2_xnor2_1 _6690_ (.Y(_2752_),
    .A(\vgademo.plane_u[4] ),
    .B(\vgademo.plane_du[4] ));
 sg13g2_nand3_1 _6691_ (.B(_2747_),
    .C(_2752_),
    .A(_2744_),
    .Y(_2753_));
 sg13g2_a21o_1 _6692_ (.A2(_2747_),
    .A1(_2744_),
    .B1(_2752_),
    .X(_2754_));
 sg13g2_and2_1 _6693_ (.A(_0580_),
    .B(_2753_),
    .X(_2755_));
 sg13g2_nor2_1 _6694_ (.A(\vgademo.plane_dx[3] ),
    .B(_2748_),
    .Y(_2756_));
 sg13g2_xnor2_1 _6695_ (.Y(_2757_),
    .A(\vgademo.plane_dx[3] ),
    .B(_2748_));
 sg13g2_a221oi_1 _6696_ (.B2(net901),
    .C1(net876),
    .B1(_2757_),
    .A1(_2754_),
    .Y(_2758_),
    .A2(_2755_));
 sg13g2_a21oi_1 _6697_ (.A1(_3174_),
    .A2(net876),
    .Y(_0334_),
    .B1(_2758_));
 sg13g2_o21ai_1 _6698_ (.B1(_2754_),
    .Y(_2759_),
    .A1(_3174_),
    .A2(_3175_));
 sg13g2_or2_1 _6699_ (.X(_2760_),
    .B(\vgademo.plane_du[5] ),
    .A(\vgademo.plane_u[5] ));
 sg13g2_nand2_1 _6700_ (.Y(_2761_),
    .A(net337),
    .B(\vgademo.plane_du[5] ));
 sg13g2_nand2_1 _6701_ (.Y(_2762_),
    .A(_2760_),
    .B(_2761_));
 sg13g2_nand2b_1 _6702_ (.Y(_2763_),
    .B(\vgademo.plane_dx[0] ),
    .A_N(_0023_));
 sg13g2_xnor2_1 _6703_ (.Y(_2764_),
    .A(\vgademo.plane_dx[0] ),
    .B(net1015));
 sg13g2_nand2_1 _6704_ (.Y(_2765_),
    .A(_0022_),
    .B(_2764_));
 sg13g2_xnor2_1 _6705_ (.Y(_2766_),
    .A(_0022_),
    .B(_2764_));
 sg13g2_o21ai_1 _6706_ (.B1(net899),
    .Y(_2767_),
    .A1(_2756_),
    .A2(_2766_));
 sg13g2_a21oi_1 _6707_ (.A1(_2756_),
    .A2(_2766_),
    .Y(_2768_),
    .B1(_2767_));
 sg13g2_nor2_1 _6708_ (.A(net876),
    .B(_2768_),
    .Y(_2769_));
 sg13g2_xnor2_1 _6709_ (.Y(_2770_),
    .A(_2759_),
    .B(_2762_));
 sg13g2_nand2_1 _6710_ (.Y(_2771_),
    .A(net892),
    .B(_2770_));
 sg13g2_a22oi_1 _6711_ (.Y(_0335_),
    .B1(_2769_),
    .B2(_2771_),
    .A2(net876),
    .A1(_3176_));
 sg13g2_nand2_1 _6712_ (.Y(_2772_),
    .A(net353),
    .B(\vgademo.plane_du[6] ));
 sg13g2_xnor2_1 _6713_ (.Y(_2773_),
    .A(\vgademo.plane_u[6] ),
    .B(\vgademo.plane_du[6] ));
 sg13g2_nand2_1 _6714_ (.Y(_2774_),
    .A(_2759_),
    .B(_2760_));
 sg13g2_nand3_1 _6715_ (.B(_2773_),
    .C(_2774_),
    .A(_2761_),
    .Y(_2775_));
 sg13g2_a21o_1 _6716_ (.A2(_2774_),
    .A1(_2761_),
    .B1(_2773_),
    .X(_2776_));
 sg13g2_nand3_1 _6717_ (.B(_2775_),
    .C(_2776_),
    .A(net892),
    .Y(_2777_));
 sg13g2_nand2_1 _6718_ (.Y(_2778_),
    .A(net1013),
    .B(\vgademo.plane_dx[1] ));
 sg13g2_xor2_1 _6719_ (.B(\vgademo.plane_dx[1] ),
    .A(net1013),
    .X(_2779_));
 sg13g2_nand2b_1 _6720_ (.Y(_2780_),
    .B(_2779_),
    .A_N(_2763_));
 sg13g2_xnor2_1 _6721_ (.Y(_2781_),
    .A(_2763_),
    .B(_2779_));
 sg13g2_xnor2_1 _6722_ (.Y(_2782_),
    .A(net950),
    .B(_2781_));
 sg13g2_nor2b_1 _6723_ (.A(_2764_),
    .B_N(_2782_),
    .Y(_2783_));
 sg13g2_xnor2_1 _6724_ (.Y(_2784_),
    .A(_2764_),
    .B(_2782_));
 sg13g2_o21ai_1 _6725_ (.B1(_2765_),
    .Y(_2785_),
    .A1(_2756_),
    .A2(_2766_));
 sg13g2_and2_1 _6726_ (.A(_2784_),
    .B(_2785_),
    .X(_2786_));
 sg13g2_o21ai_1 _6727_ (.B1(net899),
    .Y(_2787_),
    .A1(_2784_),
    .A2(_2785_));
 sg13g2_nor2_1 _6728_ (.A(_2786_),
    .B(_2787_),
    .Y(_2788_));
 sg13g2_nor2_1 _6729_ (.A(net877),
    .B(_2788_),
    .Y(_2789_));
 sg13g2_a22oi_1 _6730_ (.Y(_0336_),
    .B1(_2777_),
    .B2(_2789_),
    .A2(net877),
    .A1(_3178_));
 sg13g2_nand2_1 _6731_ (.Y(_2790_),
    .A(\vgademo.plane_u[7] ),
    .B(\vgademo.plane_du[7] ));
 sg13g2_xnor2_1 _6732_ (.Y(_2791_),
    .A(\vgademo.plane_u[7] ),
    .B(\vgademo.plane_du[7] ));
 sg13g2_nand3_1 _6733_ (.B(_2776_),
    .C(_2791_),
    .A(_2772_),
    .Y(_2792_));
 sg13g2_a21o_1 _6734_ (.A2(_2776_),
    .A1(_2772_),
    .B1(_2791_),
    .X(_2793_));
 sg13g2_nand3_1 _6735_ (.B(_2792_),
    .C(_2793_),
    .A(net892),
    .Y(_2794_));
 sg13g2_nor2_1 _6736_ (.A(_2783_),
    .B(_2786_),
    .Y(_2795_));
 sg13g2_nand2_1 _6737_ (.Y(_2796_),
    .A(\vgademo.plane_dx[0] ),
    .B(_2781_));
 sg13g2_xnor2_1 _6738_ (.Y(_2797_),
    .A(\vgademo.plane_dx_div.q[5] ),
    .B(\vgademo.plane_dx[2] ));
 sg13g2_a21oi_1 _6739_ (.A1(_2778_),
    .A2(_2780_),
    .Y(_2798_),
    .B1(_2797_));
 sg13g2_nand3_1 _6740_ (.B(_2780_),
    .C(_2797_),
    .A(_2778_),
    .Y(_2799_));
 sg13g2_nor2b_1 _6741_ (.A(_2798_),
    .B_N(_2799_),
    .Y(_2800_));
 sg13g2_xnor2_1 _6742_ (.Y(_2801_),
    .A(_0024_),
    .B(_2800_));
 sg13g2_nand2b_1 _6743_ (.Y(_2802_),
    .B(_2796_),
    .A_N(_2801_));
 sg13g2_xor2_1 _6744_ (.B(_2801_),
    .A(_2796_),
    .X(_2803_));
 sg13g2_xor2_1 _6745_ (.B(_2803_),
    .A(_2782_),
    .X(_2804_));
 sg13g2_nor2b_1 _6746_ (.A(_2804_),
    .B_N(_2795_),
    .Y(_2805_));
 sg13g2_nor2b_1 _6747_ (.A(_2795_),
    .B_N(_2804_),
    .Y(_2806_));
 sg13g2_inv_1 _6748_ (.Y(_2807_),
    .A(_2806_));
 sg13g2_nor3_1 _6749_ (.A(net895),
    .B(_2805_),
    .C(_2806_),
    .Y(_2808_));
 sg13g2_nor2_1 _6750_ (.A(net876),
    .B(_2808_),
    .Y(_2809_));
 sg13g2_a22oi_1 _6751_ (.Y(_0337_),
    .B1(_2794_),
    .B2(_2809_),
    .A2(net876),
    .A1(_3180_));
 sg13g2_xnor2_1 _6752_ (.Y(_2810_),
    .A(\vgademo.plane_u[8] ),
    .B(\vgademo.plane_du[8] ));
 sg13g2_a21oi_1 _6753_ (.A1(_2790_),
    .A2(_2793_),
    .Y(_2811_),
    .B1(_2810_));
 sg13g2_nand3_1 _6754_ (.B(_2793_),
    .C(_2810_),
    .A(_2790_),
    .Y(_2812_));
 sg13g2_nor2_1 _6755_ (.A(net899),
    .B(_2811_),
    .Y(_2813_));
 sg13g2_o21ai_1 _6756_ (.B1(_2807_),
    .Y(_2814_),
    .A1(_2782_),
    .A2(_2803_));
 sg13g2_nand2_1 _6757_ (.Y(_2815_),
    .A(\vgademo.plane_dx[1] ),
    .B(_2800_));
 sg13g2_a21oi_1 _6758_ (.A1(net1012),
    .A2(_3183_),
    .Y(_2816_),
    .B1(_2798_));
 sg13g2_xor2_1 _6759_ (.B(\vgademo.plane_dx[3] ),
    .A(net1011),
    .X(_2817_));
 sg13g2_nand2b_1 _6760_ (.Y(_2818_),
    .B(_2817_),
    .A_N(_2816_));
 sg13g2_xnor2_1 _6761_ (.Y(_2819_),
    .A(_2816_),
    .B(_2817_));
 sg13g2_xnor2_1 _6762_ (.Y(_2820_),
    .A(_0025_),
    .B(_2819_));
 sg13g2_nand2b_1 _6763_ (.Y(_2821_),
    .B(_2815_),
    .A_N(_2820_));
 sg13g2_xor2_1 _6764_ (.B(_2820_),
    .A(_2815_),
    .X(_2822_));
 sg13g2_xor2_1 _6765_ (.B(_2822_),
    .A(_2802_),
    .X(_2823_));
 sg13g2_nor2_1 _6766_ (.A(_2814_),
    .B(_2823_),
    .Y(_2824_));
 sg13g2_nand2_1 _6767_ (.Y(_2825_),
    .A(_2814_),
    .B(_2823_));
 sg13g2_nor2_1 _6768_ (.A(net895),
    .B(_2824_),
    .Y(_2826_));
 sg13g2_a221oi_1 _6769_ (.B2(_2826_),
    .C1(net877),
    .B1(_2825_),
    .A1(_2812_),
    .Y(_2827_),
    .A2(_2813_));
 sg13g2_a21oi_1 _6770_ (.A1(_3182_),
    .A2(net877),
    .Y(_0338_),
    .B1(_2827_));
 sg13g2_a21oi_2 _6771_ (.B1(_2811_),
    .Y(_2828_),
    .A2(\vgademo.plane_du[8] ),
    .A1(\vgademo.plane_u[8] ));
 sg13g2_nand2_1 _6772_ (.Y(_2829_),
    .A(_3184_),
    .B(_3185_));
 sg13g2_xor2_1 _6773_ (.B(\vgademo.plane_du[9] ),
    .A(\vgademo.plane_u[9] ),
    .X(_2830_));
 sg13g2_xnor2_1 _6774_ (.Y(_2831_),
    .A(_2828_),
    .B(_2830_));
 sg13g2_o21ai_1 _6775_ (.B1(_2825_),
    .Y(_2832_),
    .A1(_2802_),
    .A2(_2822_));
 sg13g2_xor2_1 _6776_ (.B(net950),
    .A(\vgademo.plane_dx[3] ),
    .X(_2833_));
 sg13g2_nor2_1 _6777_ (.A(net1015),
    .B(_0026_),
    .Y(_2834_));
 sg13g2_nand2_1 _6778_ (.Y(_2835_),
    .A(net1015),
    .B(_0026_));
 sg13g2_nand2b_1 _6779_ (.Y(_2836_),
    .B(_2835_),
    .A_N(_2834_));
 sg13g2_o21ai_1 _6780_ (.B1(_2818_),
    .Y(_2837_),
    .A1(_3096_),
    .A2(_0022_));
 sg13g2_xnor2_1 _6781_ (.Y(_2838_),
    .A(_2836_),
    .B(_2837_));
 sg13g2_nor2_1 _6782_ (.A(_2833_),
    .B(_2838_),
    .Y(_2839_));
 sg13g2_xnor2_1 _6783_ (.Y(_2840_),
    .A(_2833_),
    .B(_2838_));
 sg13g2_nand2_1 _6784_ (.Y(_2841_),
    .A(\vgademo.plane_dx[2] ),
    .B(_2819_));
 sg13g2_nand2b_1 _6785_ (.Y(_2842_),
    .B(_2841_),
    .A_N(_2840_));
 sg13g2_xor2_1 _6786_ (.B(_2841_),
    .A(_2840_),
    .X(_2843_));
 sg13g2_nor2_1 _6787_ (.A(_2821_),
    .B(_2843_),
    .Y(_2844_));
 sg13g2_xor2_1 _6788_ (.B(_2843_),
    .A(_2821_),
    .X(_2845_));
 sg13g2_nor2_1 _6789_ (.A(_2832_),
    .B(_2845_),
    .Y(_2846_));
 sg13g2_nand2_1 _6790_ (.Y(_2847_),
    .A(_2832_),
    .B(_2845_));
 sg13g2_nor2_1 _6791_ (.A(net896),
    .B(_2846_),
    .Y(_2848_));
 sg13g2_a221oi_1 _6792_ (.B2(_2848_),
    .C1(net879),
    .B1(_2847_),
    .A1(net896),
    .Y(_2849_),
    .A2(_2831_));
 sg13g2_a21oi_1 _6793_ (.A1(_3184_),
    .A2(net878),
    .Y(_0339_),
    .B1(_2849_));
 sg13g2_nand2_1 _6794_ (.Y(_2850_),
    .A(\vgademo.plane_u[10] ),
    .B(\vgademo.plane_du[10] ));
 sg13g2_xor2_1 _6795_ (.B(\vgademo.plane_du[10] ),
    .A(\vgademo.plane_u[10] ),
    .X(_2851_));
 sg13g2_o21ai_1 _6796_ (.B1(_2828_),
    .Y(_2852_),
    .A1(_3184_),
    .A2(_3185_));
 sg13g2_a21oi_1 _6797_ (.A1(_2829_),
    .A2(_2852_),
    .Y(_2853_),
    .B1(_2851_));
 sg13g2_nand3_1 _6798_ (.B(_2851_),
    .C(_2852_),
    .A(_2829_),
    .Y(_2854_));
 sg13g2_nor2_1 _6799_ (.A(net900),
    .B(_2853_),
    .Y(_2855_));
 sg13g2_a21oi_1 _6800_ (.A1(_2832_),
    .A2(_2845_),
    .Y(_2856_),
    .B1(_2844_));
 sg13g2_xor2_1 _6801_ (.B(net1015),
    .A(\vgademo.plane_dx[1] ),
    .X(_2857_));
 sg13g2_a21oi_1 _6802_ (.A1(_2835_),
    .A2(_2837_),
    .Y(_2858_),
    .B1(_2834_));
 sg13g2_nand2_1 _6803_ (.Y(_2859_),
    .A(net1009),
    .B(net1013));
 sg13g2_nor2_1 _6804_ (.A(net1009),
    .B(net1013),
    .Y(_2860_));
 sg13g2_xor2_1 _6805_ (.B(net1013),
    .A(net1009),
    .X(_2861_));
 sg13g2_xnor2_1 _6806_ (.Y(_2862_),
    .A(_2858_),
    .B(_2861_));
 sg13g2_nor2_1 _6807_ (.A(_2857_),
    .B(_2862_),
    .Y(_2863_));
 sg13g2_xor2_1 _6808_ (.B(_2862_),
    .A(_2857_),
    .X(_2864_));
 sg13g2_a21oi_1 _6809_ (.A1(_3097_),
    .A2(net950),
    .Y(_2865_),
    .B1(_2839_));
 sg13g2_nand2b_1 _6810_ (.Y(_2866_),
    .B(_2864_),
    .A_N(_2865_));
 sg13g2_xor2_1 _6811_ (.B(_2865_),
    .A(_2864_),
    .X(_2867_));
 sg13g2_nor2_1 _6812_ (.A(_2842_),
    .B(_2867_),
    .Y(_2868_));
 sg13g2_xnor2_1 _6813_ (.Y(_2869_),
    .A(_2842_),
    .B(_2867_));
 sg13g2_or2_1 _6814_ (.X(_2870_),
    .B(_2869_),
    .A(_2856_));
 sg13g2_a21oi_1 _6815_ (.A1(_2856_),
    .A2(_2869_),
    .Y(_2871_),
    .B1(net896));
 sg13g2_a221oi_1 _6816_ (.B2(_2871_),
    .C1(net878),
    .B1(_2870_),
    .A1(_2854_),
    .Y(_2872_),
    .A2(_2855_));
 sg13g2_a21oi_1 _6817_ (.A1(_3186_),
    .A2(net878),
    .Y(_0340_),
    .B1(_2872_));
 sg13g2_a21oi_2 _6818_ (.B1(_0027_),
    .Y(_2873_),
    .A2(_2854_),
    .A1(_2850_));
 sg13g2_nand3_1 _6819_ (.B(_2850_),
    .C(_2854_),
    .A(_0027_),
    .Y(_2874_));
 sg13g2_nor2_1 _6820_ (.A(net900),
    .B(_2873_),
    .Y(_2875_));
 sg13g2_nor2b_1 _6821_ (.A(_2868_),
    .B_N(_2870_),
    .Y(_2876_));
 sg13g2_xnor2_1 _6822_ (.Y(_2877_),
    .A(\vgademo.plane_dx_div.q[9] ),
    .B(net1012));
 sg13g2_o21ai_1 _6823_ (.B1(_2859_),
    .Y(_2878_),
    .A1(_2858_),
    .A2(_2860_));
 sg13g2_nor2b_1 _6824_ (.A(_2877_),
    .B_N(_2878_),
    .Y(_2879_));
 sg13g2_xor2_1 _6825_ (.B(_2878_),
    .A(_2877_),
    .X(_2880_));
 sg13g2_xor2_1 _6826_ (.B(\vgademo.plane_dx[2] ),
    .A(net1014),
    .X(_2881_));
 sg13g2_nand2_1 _6827_ (.Y(_2882_),
    .A(_2880_),
    .B(_2881_));
 sg13g2_xnor2_1 _6828_ (.Y(_2883_),
    .A(_2880_),
    .B(_2881_));
 sg13g2_a21oi_2 _6829_ (.B1(_2863_),
    .Y(_2884_),
    .A2(_0024_),
    .A1(net1015));
 sg13g2_nor2_1 _6830_ (.A(_2883_),
    .B(_2884_),
    .Y(_2885_));
 sg13g2_xnor2_1 _6831_ (.Y(_2886_),
    .A(_2883_),
    .B(_2884_));
 sg13g2_xnor2_1 _6832_ (.Y(_2887_),
    .A(_2866_),
    .B(_2886_));
 sg13g2_nor2_1 _6833_ (.A(_2876_),
    .B(_2887_),
    .Y(_2888_));
 sg13g2_inv_1 _6834_ (.Y(_2889_),
    .A(_2888_));
 sg13g2_a21oi_1 _6835_ (.A1(_2876_),
    .A2(_2887_),
    .Y(_2890_),
    .B1(net896));
 sg13g2_a221oi_1 _6836_ (.B2(_2890_),
    .C1(net878),
    .B1(_2889_),
    .A1(_2874_),
    .Y(_2891_),
    .A2(_2875_));
 sg13g2_a21oi_1 _6837_ (.A1(_3187_),
    .A2(net879),
    .Y(_0341_),
    .B1(_2891_));
 sg13g2_xnor2_1 _6838_ (.Y(_2892_),
    .A(_0028_),
    .B(_2873_));
 sg13g2_o21ai_1 _6839_ (.B1(_2889_),
    .Y(_2893_),
    .A1(_2866_),
    .A2(_2886_));
 sg13g2_a21oi_1 _6840_ (.A1(net1007),
    .A2(net1012),
    .Y(_2894_),
    .B1(_2879_));
 sg13g2_nand2b_1 _6841_ (.Y(_2895_),
    .B(net1011),
    .A_N(_2894_));
 sg13g2_xnor2_1 _6842_ (.Y(_2896_),
    .A(net1011),
    .B(_2894_));
 sg13g2_xor2_1 _6843_ (.B(\vgademo.plane_dx[3] ),
    .A(net1012),
    .X(_2897_));
 sg13g2_nand2b_1 _6844_ (.Y(_2898_),
    .B(_2897_),
    .A_N(_2896_));
 sg13g2_xnor2_1 _6845_ (.Y(_2899_),
    .A(_2896_),
    .B(_2897_));
 sg13g2_o21ai_1 _6846_ (.B1(_2882_),
    .Y(_2900_),
    .A1(net1013),
    .A2(_3183_));
 sg13g2_nand2_1 _6847_ (.Y(_2901_),
    .A(_2899_),
    .B(_2900_));
 sg13g2_inv_1 _6848_ (.Y(_2902_),
    .A(_2901_));
 sg13g2_xor2_1 _6849_ (.B(_2900_),
    .A(_2899_),
    .X(_2903_));
 sg13g2_xnor2_1 _6850_ (.Y(_2904_),
    .A(_2885_),
    .B(_2903_));
 sg13g2_nand2b_1 _6851_ (.Y(_2905_),
    .B(_2904_),
    .A_N(_2893_));
 sg13g2_nor2b_1 _6852_ (.A(_2904_),
    .B_N(_2893_),
    .Y(_2906_));
 sg13g2_nor2_1 _6853_ (.A(net896),
    .B(_2906_),
    .Y(_2907_));
 sg13g2_a221oi_1 _6854_ (.B2(_2907_),
    .C1(net879),
    .B1(_2905_),
    .A1(net896),
    .Y(_2908_),
    .A2(_2892_));
 sg13g2_a21oi_1 _6855_ (.A1(_3188_),
    .A2(net879),
    .Y(_0342_),
    .B1(_2908_));
 sg13g2_a21oi_1 _6856_ (.A1(_2885_),
    .A2(_2903_),
    .Y(_2909_),
    .B1(_2906_));
 sg13g2_nand2_1 _6857_ (.Y(_2910_),
    .A(_3096_),
    .B(net1015));
 sg13g2_xor2_1 _6858_ (.B(net1015),
    .A(net1011),
    .X(_2911_));
 sg13g2_nor2_1 _6859_ (.A(net1010),
    .B(_2895_),
    .Y(_2912_));
 sg13g2_xor2_1 _6860_ (.B(_2895_),
    .A(net1010),
    .X(_2913_));
 sg13g2_xor2_1 _6861_ (.B(_2913_),
    .A(_2911_),
    .X(_2914_));
 sg13g2_o21ai_1 _6862_ (.B1(_2898_),
    .Y(_2915_),
    .A1(net1012),
    .A2(_3177_));
 sg13g2_nand2_1 _6863_ (.Y(_2916_),
    .A(_2914_),
    .B(_2915_));
 sg13g2_xor2_1 _6864_ (.B(_2915_),
    .A(_2914_),
    .X(_2917_));
 sg13g2_xnor2_1 _6865_ (.Y(_2918_),
    .A(_2901_),
    .B(_2917_));
 sg13g2_nand2b_1 _6866_ (.Y(_2919_),
    .B(_2909_),
    .A_N(_2918_));
 sg13g2_nor2b_1 _6867_ (.A(_2909_),
    .B_N(_2918_),
    .Y(_2920_));
 sg13g2_nor2_1 _6868_ (.A(net895),
    .B(_2920_),
    .Y(_2921_));
 sg13g2_a21oi_1 _6869_ (.A1(net360),
    .A2(_2873_),
    .Y(_2922_),
    .B1(net381));
 sg13g2_nand3_1 _6870_ (.B(\vgademo.plane_u[13] ),
    .C(_2873_),
    .A(\vgademo.plane_u[12] ),
    .Y(_2923_));
 sg13g2_nor2b_1 _6871_ (.A(_2922_),
    .B_N(_2923_),
    .Y(_2924_));
 sg13g2_a221oi_1 _6872_ (.B2(net895),
    .C1(net878),
    .B1(_2924_),
    .A1(_2919_),
    .Y(_2925_),
    .A2(_2921_));
 sg13g2_a21oi_1 _6873_ (.A1(_3189_),
    .A2(net878),
    .Y(_0343_),
    .B1(_2925_));
 sg13g2_a21oi_1 _6874_ (.A1(_2902_),
    .A2(_2917_),
    .Y(_2926_),
    .B1(_2920_));
 sg13g2_nor2b_1 _6875_ (.A(net1014),
    .B_N(net1010),
    .Y(_2927_));
 sg13g2_xnor2_1 _6876_ (.Y(_2928_),
    .A(net1014),
    .B(net1010));
 sg13g2_and2_1 _6877_ (.A(net1009),
    .B(_2912_),
    .X(_2929_));
 sg13g2_xnor2_1 _6878_ (.Y(_2930_),
    .A(net1008),
    .B(_2912_));
 sg13g2_xor2_1 _6879_ (.B(_2930_),
    .A(_2928_),
    .X(_2931_));
 sg13g2_o21ai_1 _6880_ (.B1(_2910_),
    .Y(_2932_),
    .A1(_2911_),
    .A2(_2913_));
 sg13g2_nand2_1 _6881_ (.Y(_2933_),
    .A(_2931_),
    .B(_2932_));
 sg13g2_xnor2_1 _6882_ (.Y(_2934_),
    .A(_2931_),
    .B(_2932_));
 sg13g2_nor2_1 _6883_ (.A(_2916_),
    .B(_2934_),
    .Y(_2935_));
 sg13g2_xor2_1 _6884_ (.B(_2934_),
    .A(_2916_),
    .X(_2936_));
 sg13g2_nor2b_1 _6885_ (.A(_2926_),
    .B_N(_2936_),
    .Y(_2937_));
 sg13g2_xor2_1 _6886_ (.B(_2936_),
    .A(_2926_),
    .X(_2938_));
 sg13g2_xnor2_1 _6887_ (.Y(_2939_),
    .A(_3190_),
    .B(_2923_));
 sg13g2_nand2_1 _6888_ (.Y(_2940_),
    .A(net893),
    .B(_2939_));
 sg13g2_a21oi_1 _6889_ (.A1(net899),
    .A2(_2938_),
    .Y(_2941_),
    .B1(net878));
 sg13g2_a22oi_1 _6890_ (.Y(_2942_),
    .B1(_2940_),
    .B2(_2941_),
    .A2(net878),
    .A1(net390));
 sg13g2_inv_1 _6891_ (.Y(_0344_),
    .A(_2942_));
 sg13g2_nor2_1 _6892_ (.A(net1008),
    .B(net1012),
    .Y(_2943_));
 sg13g2_xor2_1 _6893_ (.B(net1012),
    .A(net1008),
    .X(_2944_));
 sg13g2_xnor2_1 _6894_ (.Y(_2945_),
    .A(net1007),
    .B(_2929_));
 sg13g2_xnor2_1 _6895_ (.Y(_2946_),
    .A(_2944_),
    .B(_2945_));
 sg13g2_a21oi_1 _6896_ (.A1(_2928_),
    .A2(_2930_),
    .Y(_2947_),
    .B1(_2927_));
 sg13g2_nor2_1 _6897_ (.A(_2946_),
    .B(_2947_),
    .Y(_2948_));
 sg13g2_xor2_1 _6898_ (.B(_2947_),
    .A(_2946_),
    .X(_2949_));
 sg13g2_nand2b_1 _6899_ (.Y(_2950_),
    .B(_2949_),
    .A_N(_2933_));
 sg13g2_xnor2_1 _6900_ (.Y(_2951_),
    .A(_2933_),
    .B(_2949_));
 sg13g2_or3_1 _6901_ (.A(_2935_),
    .B(_2937_),
    .C(_2951_),
    .X(_2952_));
 sg13g2_o21ai_1 _6902_ (.B1(_2951_),
    .Y(_2953_),
    .A1(_2935_),
    .A2(_2937_));
 sg13g2_nand3_1 _6903_ (.B(_2952_),
    .C(_2953_),
    .A(net899),
    .Y(_2954_));
 sg13g2_nor2_1 _6904_ (.A(_0029_),
    .B(_2923_),
    .Y(_2955_));
 sg13g2_xnor2_1 _6905_ (.Y(_2956_),
    .A(_3191_),
    .B(_2955_));
 sg13g2_a21oi_1 _6906_ (.A1(net895),
    .A2(_2956_),
    .Y(_2957_),
    .B1(net875));
 sg13g2_a22oi_1 _6907_ (.Y(_0345_),
    .B1(_2954_),
    .B2(_2957_),
    .A2(net875),
    .A1(_3191_));
 sg13g2_nand2_2 _6908_ (.Y(_2958_),
    .A(net1007),
    .B(net1011));
 sg13g2_or2_1 _6909_ (.X(_2959_),
    .B(net1011),
    .A(net1007));
 sg13g2_a21oi_1 _6910_ (.A1(_2958_),
    .A2(_2959_),
    .Y(_2960_),
    .B1(_2929_));
 sg13g2_a21oi_1 _6911_ (.A1(_2944_),
    .A2(_2945_),
    .Y(_2961_),
    .B1(_2943_));
 sg13g2_nor2b_1 _6912_ (.A(_2961_),
    .B_N(_2960_),
    .Y(_2962_));
 sg13g2_xnor2_1 _6913_ (.Y(_2963_),
    .A(_2960_),
    .B(_2961_));
 sg13g2_nand2_1 _6914_ (.Y(_2964_),
    .A(_2948_),
    .B(_2963_));
 sg13g2_xnor2_1 _6915_ (.Y(_2965_),
    .A(_2948_),
    .B(_2963_));
 sg13g2_a21o_1 _6916_ (.A2(_2953_),
    .A1(_2950_),
    .B1(_2965_),
    .X(_2966_));
 sg13g2_nand3_1 _6917_ (.B(_2953_),
    .C(_2965_),
    .A(_2950_),
    .Y(_2967_));
 sg13g2_nor3_2 _6918_ (.A(_3190_),
    .B(_3191_),
    .C(_2923_),
    .Y(_2968_));
 sg13g2_a21o_1 _6919_ (.A2(_2967_),
    .A1(_2966_),
    .B1(net895),
    .X(_2969_));
 sg13g2_xor2_1 _6920_ (.B(_2968_),
    .A(_0030_),
    .X(_2970_));
 sg13g2_a21oi_1 _6921_ (.A1(net892),
    .A2(_2970_),
    .Y(_2971_),
    .B1(net875));
 sg13g2_a22oi_1 _6922_ (.Y(_2972_),
    .B1(_2969_),
    .B2(_2971_),
    .A2(net875),
    .A1(net425));
 sg13g2_inv_1 _6923_ (.Y(_0346_),
    .A(net426));
 sg13g2_nand3_1 _6924_ (.B(\vgademo.plane_u[17] ),
    .C(_2968_),
    .A(\vgademo.plane_u[16] ),
    .Y(_2973_));
 sg13g2_inv_1 _6925_ (.Y(_2974_),
    .A(_2973_));
 sg13g2_a21oi_1 _6926_ (.A1(\vgademo.plane_u[16] ),
    .A2(_2968_),
    .Y(_2975_),
    .B1(\vgademo.plane_u[17] ));
 sg13g2_nor2_1 _6927_ (.A(net901),
    .B(_2975_),
    .Y(_2976_));
 sg13g2_nand2_1 _6928_ (.Y(_2977_),
    .A(net1010),
    .B(_2958_));
 sg13g2_xor2_1 _6929_ (.B(_2958_),
    .A(net1010),
    .X(_2978_));
 sg13g2_xnor2_1 _6930_ (.Y(_2979_),
    .A(_2962_),
    .B(_2978_));
 sg13g2_and3_1 _6931_ (.X(_2980_),
    .A(_2964_),
    .B(_2966_),
    .C(_2979_));
 sg13g2_a21oi_1 _6932_ (.A1(_2964_),
    .A2(_2966_),
    .Y(_2981_),
    .B1(_2979_));
 sg13g2_nor2_1 _6933_ (.A(_2980_),
    .B(_2981_),
    .Y(_2982_));
 sg13g2_a221oi_1 _6934_ (.B2(net901),
    .C1(net874),
    .B1(_2982_),
    .A1(_2973_),
    .Y(_2983_),
    .A2(_2976_));
 sg13g2_a21oi_1 _6935_ (.A1(_3192_),
    .A2(net874),
    .Y(_0347_),
    .B1(_2983_));
 sg13g2_nand3_1 _6936_ (.B(net1010),
    .C(_2958_),
    .A(net1008),
    .Y(_2984_));
 sg13g2_xor2_1 _6937_ (.B(_2977_),
    .A(net1008),
    .X(_2985_));
 sg13g2_a21oi_2 _6938_ (.B1(_2981_),
    .Y(_2986_),
    .A2(_2978_),
    .A1(_2962_));
 sg13g2_xnor2_1 _6939_ (.Y(_2987_),
    .A(_2985_),
    .B(_2986_));
 sg13g2_xor2_1 _6940_ (.B(_2973_),
    .A(\vgademo.plane_u[18] ),
    .X(_2988_));
 sg13g2_nand2_1 _6941_ (.Y(_2989_),
    .A(net892),
    .B(_2988_));
 sg13g2_a21oi_1 _6942_ (.A1(net901),
    .A2(_2987_),
    .Y(_2990_),
    .B1(net875));
 sg13g2_a22oi_1 _6943_ (.Y(_2991_),
    .B1(_2989_),
    .B2(_2990_),
    .A2(net874),
    .A1(net506));
 sg13g2_inv_1 _6944_ (.Y(_0348_),
    .A(_2991_));
 sg13g2_o21ai_1 _6945_ (.B1(_2984_),
    .Y(_2992_),
    .A1(_2985_),
    .A2(_2986_));
 sg13g2_nand2_1 _6946_ (.Y(_2993_),
    .A(net1007),
    .B(net1008));
 sg13g2_xor2_1 _6947_ (.B(net1008),
    .A(net1007),
    .X(_2994_));
 sg13g2_nor2_1 _6948_ (.A(_0031_),
    .B(_2973_),
    .Y(_2995_));
 sg13g2_xnor2_1 _6949_ (.Y(_2996_),
    .A(_2992_),
    .B(_2994_));
 sg13g2_nand2_1 _6950_ (.Y(_2997_),
    .A(net901),
    .B(_2996_));
 sg13g2_xnor2_1 _6951_ (.Y(_2998_),
    .A(_3193_),
    .B(_2995_));
 sg13g2_a21oi_1 _6952_ (.A1(net892),
    .A2(_2998_),
    .Y(_2999_),
    .B1(net874));
 sg13g2_a22oi_1 _6953_ (.Y(_0349_),
    .B1(_2997_),
    .B2(_2999_),
    .A2(net874),
    .A1(_3193_));
 sg13g2_nor4_1 _6954_ (.A(net1007),
    .B(net1008),
    .C(_2977_),
    .D(_2986_),
    .Y(_3000_));
 sg13g2_nor2_1 _6955_ (.A(net892),
    .B(_3000_),
    .Y(_3001_));
 sg13g2_o21ai_1 _6956_ (.B1(_3001_),
    .Y(_3002_),
    .A1(_2992_),
    .A2(_2993_));
 sg13g2_nand3_1 _6957_ (.B(\vgademo.plane_u[19] ),
    .C(_2974_),
    .A(\vgademo.plane_u[18] ),
    .Y(_3003_));
 sg13g2_xnor2_1 _6958_ (.Y(_3004_),
    .A(net328),
    .B(_3003_));
 sg13g2_a21oi_1 _6959_ (.A1(net892),
    .A2(_3004_),
    .Y(_3005_),
    .B1(net874));
 sg13g2_a22oi_1 _6960_ (.Y(_0350_),
    .B1(_3002_),
    .B2(_3005_),
    .A2(net874),
    .A1(_3194_));
 sg13g2_nor2_1 _6961_ (.A(_0032_),
    .B(_3003_),
    .Y(_3006_));
 sg13g2_a21oi_1 _6962_ (.A1(net399),
    .A2(_3006_),
    .Y(_3007_),
    .B1(net901));
 sg13g2_o21ai_1 _6963_ (.B1(_3007_),
    .Y(_3008_),
    .A1(net399),
    .A2(_3006_));
 sg13g2_nor2_1 _6964_ (.A(net875),
    .B(_3001_),
    .Y(_3009_));
 sg13g2_a22oi_1 _6965_ (.Y(_0351_),
    .B1(_3008_),
    .B2(_3009_),
    .A2(net874),
    .A1(_3195_));
 sg13g2_xor2_1 _6966_ (.B(_1808_),
    .A(_1804_),
    .X(_3010_));
 sg13g2_o21ai_1 _6967_ (.B1(_2237_),
    .Y(_3011_),
    .A1(_2190_),
    .A2(_3010_));
 sg13g2_nand3_1 _6968_ (.B(_1801_),
    .C(_1810_),
    .A(_1800_),
    .Y(_3012_));
 sg13g2_nor2b_2 _6969_ (.A(_1811_),
    .B_N(_3012_),
    .Y(_3013_));
 sg13g2_a21oi_2 _6970_ (.B1(_2216_),
    .Y(_3014_),
    .A2(_3013_),
    .A1(_2189_));
 sg13g2_nor4_1 _6971_ (.A(net816),
    .B(net813),
    .C(_1784_),
    .D(_3014_),
    .Y(_3015_));
 sg13g2_a221oi_1 _6972_ (.B2(_3011_),
    .C1(_3015_),
    .B1(net811),
    .A1(net855),
    .Y(_3016_),
    .A2(net853));
 sg13g2_o21ai_1 _6973_ (.B1(_1329_),
    .Y(_3017_),
    .A1(_2171_),
    .A2(_3016_));
 sg13g2_and2_1 _6974_ (.A(net935),
    .B(_3017_),
    .X(_3018_));
 sg13g2_xnor2_1 _6975_ (.Y(_3019_),
    .A(_1799_),
    .B(_1812_));
 sg13g2_a21oi_2 _6976_ (.B1(_2193_),
    .Y(_3020_),
    .A2(_3019_),
    .A1(_2189_));
 sg13g2_nor4_1 _6977_ (.A(net816),
    .B(net813),
    .C(_1784_),
    .D(_3020_),
    .Y(_3021_));
 sg13g2_nand3_1 _6978_ (.B(_1803_),
    .C(_1809_),
    .A(_1802_),
    .Y(_3022_));
 sg13g2_nand2_2 _6979_ (.Y(_3023_),
    .A(_1810_),
    .B(_3022_));
 sg13g2_o21ai_1 _6980_ (.B1(_2228_),
    .Y(_3024_),
    .A1(_2190_),
    .A2(_3023_));
 sg13g2_a221oi_1 _6981_ (.B2(_3024_),
    .C1(_3021_),
    .B1(net811),
    .A1(net855),
    .Y(_3025_),
    .A2(net854));
 sg13g2_o21ai_1 _6982_ (.B1(_1329_),
    .Y(_3026_),
    .A1(_2222_),
    .A2(_3025_));
 sg13g2_xor2_1 _6983_ (.B(_3017_),
    .A(_2236_),
    .X(_3027_));
 sg13g2_a21o_1 _6984_ (.A2(_3027_),
    .A1(_3026_),
    .B1(_3018_),
    .X(_3028_));
 sg13g2_o21ai_1 _6985_ (.B1(_1870_),
    .Y(_3029_),
    .A1(_1818_),
    .A2(_1837_));
 sg13g2_nor4_1 _6986_ (.A(net814),
    .B(net813),
    .C(_1784_),
    .D(_3029_),
    .Y(_3030_));
 sg13g2_a221oi_1 _6987_ (.B2(_3020_),
    .C1(_3030_),
    .B1(net811),
    .A1(net856),
    .Y(_3031_),
    .A2(net853));
 sg13g2_or2_1 _6988_ (.X(_3032_),
    .B(_2198_),
    .A(_1761_));
 sg13g2_o21ai_1 _6989_ (.B1(_2184_),
    .Y(_3033_),
    .A1(_3031_),
    .A2(_3032_));
 sg13g2_nand2_2 _6990_ (.Y(_3034_),
    .A(net858),
    .B(_3033_));
 sg13g2_or2_1 _6991_ (.X(_3035_),
    .B(_2188_),
    .A(_2167_));
 sg13g2_inv_1 _6992_ (.Y(_3036_),
    .A(_3035_));
 sg13g2_mux2_1 _6993_ (.A0(_3014_),
    .A1(_3036_),
    .S(_1785_),
    .X(_3037_));
 sg13g2_a21o_1 _6994_ (.A2(_3037_),
    .A1(net847),
    .B1(_2210_),
    .X(_3038_));
 sg13g2_a21oi_2 _6995_ (.B1(_1332_),
    .Y(_3039_),
    .A2(_3038_),
    .A1(_2162_));
 sg13g2_and2_1 _6996_ (.A(_2251_),
    .B(_3039_),
    .X(_3040_));
 sg13g2_xnor2_1 _6997_ (.Y(_3041_),
    .A(_2250_),
    .B(_3039_));
 sg13g2_xor2_1 _6998_ (.B(_3041_),
    .A(_3034_),
    .X(_3042_));
 sg13g2_and2_1 _6999_ (.A(net848),
    .B(_3029_),
    .X(_3043_));
 sg13g2_a221oi_1 _7000_ (.B2(net810),
    .C1(_1761_),
    .B1(_3043_),
    .A1(_1354_),
    .Y(_3044_),
    .A2(_2143_));
 sg13g2_and2_1 _7001_ (.A(_2158_),
    .B(_2183_),
    .X(_3045_));
 sg13g2_nor2_1 _7002_ (.A(_3044_),
    .B(_3045_),
    .Y(_3046_));
 sg13g2_o21ai_1 _7003_ (.B1(net858),
    .Y(_3047_),
    .A1(_3044_),
    .A2(_3045_));
 sg13g2_and2_1 _7004_ (.A(_1331_),
    .B(_3047_),
    .X(_3048_));
 sg13g2_a21o_1 _7005_ (.A2(_3047_),
    .A1(_1331_),
    .B1(_2232_),
    .X(_3049_));
 sg13g2_a21o_1 _7006_ (.A2(_3046_),
    .A1(_2232_),
    .B1(_3026_),
    .X(_3050_));
 sg13g2_nand3_1 _7007_ (.B(_3049_),
    .C(_3050_),
    .A(_3039_),
    .Y(_3051_));
 sg13g2_xnor2_1 _7008_ (.Y(_3052_),
    .A(_3026_),
    .B(_3027_));
 sg13g2_a21oi_1 _7009_ (.A1(_3049_),
    .A2(_3050_),
    .Y(_3053_),
    .B1(_3039_));
 sg13g2_a21oi_1 _7010_ (.A1(_3051_),
    .A2(_3052_),
    .Y(_3054_),
    .B1(_3053_));
 sg13g2_o21ai_1 _7011_ (.B1(_3054_),
    .Y(_3055_),
    .A1(_3028_),
    .A2(_3042_));
 sg13g2_o21ai_1 _7012_ (.B1(net848),
    .Y(_3056_),
    .A1(_1785_),
    .A2(_3036_));
 sg13g2_or2_1 _7013_ (.X(_3057_),
    .B(_2160_),
    .A(_1328_));
 sg13g2_a221oi_1 _7014_ (.B2(_2173_),
    .C1(_3057_),
    .B1(_3056_),
    .A1(_2150_),
    .Y(_3058_),
    .A2(_2183_));
 sg13g2_or2_1 _7015_ (.X(_3059_),
    .B(_3058_),
    .A(_1332_));
 sg13g2_a21o_1 _7016_ (.A2(_3033_),
    .A1(net858),
    .B1(net936),
    .X(_3060_));
 sg13g2_and3_1 _7017_ (.X(_3061_),
    .A(net858),
    .B(net936),
    .C(_3033_));
 sg13g2_xnor2_1 _7018_ (.Y(_3062_),
    .A(net936),
    .B(_3034_));
 sg13g2_xnor2_1 _7019_ (.Y(_3063_),
    .A(_3059_),
    .B(_3062_));
 sg13g2_a21o_1 _7020_ (.A2(_3041_),
    .A1(_3034_),
    .B1(_3040_),
    .X(_3064_));
 sg13g2_a22oi_1 _7021_ (.Y(_3065_),
    .B1(_3063_),
    .B2(_3064_),
    .A2(_3042_),
    .A1(_3028_));
 sg13g2_o21ai_1 _7022_ (.B1(_3060_),
    .Y(_3066_),
    .A1(_3059_),
    .A2(_3061_));
 sg13g2_or3_1 _7023_ (.A(_1332_),
    .B(_2178_),
    .C(_3058_),
    .X(_3067_));
 sg13g2_o21ai_1 _7024_ (.B1(_2178_),
    .Y(_3068_),
    .A1(_1332_),
    .A2(_3058_));
 sg13g2_nand3_1 _7025_ (.B(_3067_),
    .C(_3068_),
    .A(_3048_),
    .Y(_3069_));
 sg13g2_a21o_1 _7026_ (.A2(_3068_),
    .A1(_3067_),
    .B1(_3048_),
    .X(_3070_));
 sg13g2_a21o_1 _7027_ (.A2(_3070_),
    .A1(_3069_),
    .B1(_3066_),
    .X(_3071_));
 sg13g2_o21ai_1 _7028_ (.B1(_3071_),
    .Y(_3072_),
    .A1(_3063_),
    .A2(_3064_));
 sg13g2_a21oi_1 _7029_ (.A1(_3055_),
    .A2(_3065_),
    .Y(_3073_),
    .B1(_3072_));
 sg13g2_a21o_1 _7030_ (.A2(_3065_),
    .A1(_3055_),
    .B1(_3072_),
    .X(_3074_));
 sg13g2_and3_1 _7031_ (.X(_3075_),
    .A(_3066_),
    .B(_3069_),
    .C(_3070_));
 sg13g2_inv_1 _7032_ (.Y(_3076_),
    .A(_3075_));
 sg13g2_nand2_1 _7033_ (.Y(_3077_),
    .A(_3048_),
    .B(_3068_));
 sg13g2_nand2b_1 _7034_ (.Y(_3078_),
    .B(_3067_),
    .A_N(_3048_));
 sg13g2_and2_1 _7035_ (.A(_3077_),
    .B(_3078_),
    .X(_3079_));
 sg13g2_inv_1 _7036_ (.Y(_3080_),
    .A(_3079_));
 sg13g2_nor3_1 _7037_ (.A(_3073_),
    .B(_3075_),
    .C(_3079_),
    .Y(_3081_));
 sg13g2_a21oi_1 _7038_ (.A1(_3074_),
    .A2(_3076_),
    .Y(_3082_),
    .B1(_3080_));
 sg13g2_o21ai_1 _7039_ (.B1(_3079_),
    .Y(_3083_),
    .A1(_3073_),
    .A2(_3075_));
 sg13g2_nor3_1 _7040_ (.A(_2270_),
    .B(_3081_),
    .C(_3082_),
    .Y(_0352_));
 sg13g2_a21oi_1 _7041_ (.A1(_3077_),
    .A2(_3083_),
    .Y(_0353_),
    .B1(_2270_));
 sg13g2_nor2_1 _7042_ (.A(net316),
    .B(net890),
    .Y(_3084_));
 sg13g2_a21oi_1 _7043_ (.A1(_3099_),
    .A2(net890),
    .Y(_0354_),
    .B1(_3084_));
 sg13g2_nor2_1 _7044_ (.A(net310),
    .B(net888),
    .Y(_3085_));
 sg13g2_a21oi_1 _7045_ (.A1(_3098_),
    .A2(net888),
    .Y(_0355_),
    .B1(_3085_));
 sg13g2_mux2_1 _7046_ (.A0(net473),
    .A1(\vgademo.plane_dx[2] ),
    .S(net888),
    .X(_0356_));
 sg13g2_nor2_1 _7047_ (.A(net457),
    .B(net888),
    .Y(_3086_));
 sg13g2_a21oi_1 _7048_ (.A1(_3097_),
    .A2(net888),
    .Y(_0357_),
    .B1(_3086_));
 sg13g2_nor2_1 _7049_ (.A(\vgademo.plane_du[4] ),
    .B(net890),
    .Y(_3087_));
 sg13g2_a21oi_1 _7050_ (.A1(net1015),
    .A2(net890),
    .Y(_0358_),
    .B1(_3087_));
 sg13g2_mux2_1 _7051_ (.A0(net562),
    .A1(net1014),
    .S(net888),
    .X(_0359_));
 sg13g2_nand2_1 _7052_ (.Y(_3088_),
    .A(net1012),
    .B(net889));
 sg13g2_o21ai_1 _7053_ (.B1(_3088_),
    .Y(_0360_),
    .A1(_3179_),
    .A2(net889));
 sg13g2_nor2_1 _7054_ (.A(net579),
    .B(net888),
    .Y(_3089_));
 sg13g2_a21oi_1 _7055_ (.A1(_3096_),
    .A2(net888),
    .Y(_0361_),
    .B1(_3089_));
 sg13g2_nor2_1 _7056_ (.A(\vgademo.plane_du[8] ),
    .B(net889),
    .Y(_3090_));
 sg13g2_a21oi_1 _7057_ (.A1(net1010),
    .A2(net889),
    .Y(_0362_),
    .B1(_3090_));
 sg13g2_nand2_1 _7058_ (.Y(_3091_),
    .A(net1009),
    .B(net889));
 sg13g2_o21ai_1 _7059_ (.B1(_3091_),
    .Y(_0363_),
    .A1(_3185_),
    .A2(net889));
 sg13g2_mux2_1 _7060_ (.A0(\vgademo.plane_du[10] ),
    .A1(net481),
    .S(net889),
    .X(_0364_));
 sg13g2_a21oi_1 _7061_ (.A1(\vgademo.plane_du[0] ),
    .A2(_2727_),
    .Y(_3092_),
    .B1(net219));
 sg13g2_a21oi_1 _7062_ (.A1(net895),
    .A2(_2728_),
    .Y(_3093_),
    .B1(net880));
 sg13g2_nor2_1 _7063_ (.A(net220),
    .B(_3093_),
    .Y(_0365_));
 sg13g2_dfrbp_1 _7064_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net25),
    .D(_0112_),
    .Q_N(_3561_),
    .Q(\vgademo.linelfsr[0] ));
 sg13g2_dfrbp_1 _7065_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net161),
    .D(net548),
    .Q_N(_3560_),
    .Q(\vgademo.linelfsr[1] ));
 sg13g2_dfrbp_1 _7066_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net159),
    .D(net389),
    .Q_N(_3559_),
    .Q(\vgademo.linelfsr[2] ));
 sg13g2_dfrbp_1 _7067_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net157),
    .D(_0115_),
    .Q_N(_3558_),
    .Q(\vgademo.linelfsr[3] ));
 sg13g2_dfrbp_1 _7068_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net155),
    .D(_0116_),
    .Q_N(_3557_),
    .Q(\vgademo.linelfsr[4] ));
 sg13g2_dfrbp_1 _7069_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net153),
    .D(net393),
    .Q_N(_3556_),
    .Q(\vgademo.linelfsr[5] ));
 sg13g2_dfrbp_1 _7070_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net151),
    .D(_0118_),
    .Q_N(_3555_),
    .Q(\vgademo.linelfsr[6] ));
 sg13g2_dfrbp_1 _7071_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net149),
    .D(net376),
    .Q_N(_3554_),
    .Q(\vgademo.linelfsr[7] ));
 sg13g2_dfrbp_1 _7072_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net147),
    .D(_0120_),
    .Q_N(_3553_),
    .Q(\vgademo.linelfsr[8] ));
 sg13g2_dfrbp_1 _7073_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0121_),
    .Q_N(_3552_),
    .Q(\vgademo.linelfsr[9] ));
 sg13g2_dfrbp_1 _7074_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net143),
    .D(net321),
    .Q_N(_3551_),
    .Q(\vgademo.linelfsr[10] ));
 sg13g2_dfrbp_1 _7075_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net141),
    .D(net332),
    .Q_N(_3550_),
    .Q(\vgademo.linelfsr[11] ));
 sg13g2_dfrbp_1 _7076_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net139),
    .D(_0124_),
    .Q_N(_3549_),
    .Q(\vgademo.linelfsr[12] ));
 sg13g2_dfrbp_1 _7077_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1043),
    .D(net210),
    .Q_N(\vgademo.audio_songpos[0] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _7078_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1044),
    .D(_0126_),
    .Q_N(\vgademo.audio_songpos[1] ),
    .Q(_0087_));
 sg13g2_dfrbp_1 _7079_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1044),
    .D(_0127_),
    .Q_N(\vgademo.audio_songpos[2] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 _7080_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1044),
    .D(_0128_),
    .Q_N(\vgademo.audio_songpos[3] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _7081_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1044),
    .D(_0129_),
    .Q_N(\vgademo.audio_songpos[4] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _7082_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1044),
    .D(_0130_),
    .Q_N(\vgademo.audio_songpos[5] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _7083_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1043),
    .D(_0131_),
    .Q_N(\vgademo.audio_songpos[6] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 _7084_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1043),
    .D(_0132_),
    .Q_N(\vgademo.audio_songpos[7] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 _7085_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net121),
    .D(_0133_),
    .Q_N(_0024_),
    .Q(\vgademo.plane_dx[1] ));
 sg13g2_dfrbp_1 _7086_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net119),
    .D(_0134_),
    .Q_N(_0025_),
    .Q(\vgademo.plane_dx[2] ));
 sg13g2_dfrbp_1 _7087_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net117),
    .D(_0135_),
    .Q_N(_0022_),
    .Q(\vgademo.plane_dx[3] ));
 sg13g2_dfrbp_1 _7088_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net115),
    .D(_0136_),
    .Q_N(_0023_),
    .Q(\vgademo.plane_dx_div.q[3] ));
 sg13g2_dfrbp_1 _7089_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net113),
    .D(_0137_),
    .Q_N(_3548_),
    .Q(\vgademo.plane_dx_div.q[4] ));
 sg13g2_dfrbp_1 _7090_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net111),
    .D(_0138_),
    .Q_N(_3547_),
    .Q(\vgademo.plane_dx_div.q[5] ));
 sg13g2_dfrbp_1 _7091_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net109),
    .D(_0139_),
    .Q_N(_3546_),
    .Q(\vgademo.plane_dx_div.q[6] ));
 sg13g2_dfrbp_1 _7092_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net107),
    .D(_0140_),
    .Q_N(_0026_),
    .Q(\vgademo.plane_dx_div.q[7] ));
 sg13g2_dfrbp_1 _7093_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net105),
    .D(_0141_),
    .Q_N(_3545_),
    .Q(\vgademo.plane_dx_div.q[8] ));
 sg13g2_dfrbp_1 _7094_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net103),
    .D(_0142_),
    .Q_N(_3544_),
    .Q(\vgademo.plane_dx_div.q[9] ));
 sg13g2_dfrbp_1 _7095_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net101),
    .D(net169),
    .Q_N(_0085_),
    .Q(\vgademo.plane_dx_div.i[0] ));
 sg13g2_dfrbp_1 _7096_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net99),
    .D(_0144_),
    .Q_N(_3543_),
    .Q(\vgademo.plane_dx_div.i[1] ));
 sg13g2_dfrbp_1 _7097_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net97),
    .D(net540),
    .Q_N(_3542_),
    .Q(\vgademo.plane_dx_div.i[2] ));
 sg13g2_dfrbp_1 _7098_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net26),
    .D(_0146_),
    .Q_N(_3562_),
    .Q(\vgademo.plane_dx_div.i[3] ));
 sg13g2_dfrbp_1 _7099_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1048),
    .D(\vgademo.soundtrack.sigma_delta_accum_[0] ),
    .Q_N(_3563_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[0] ));
 sg13g2_dfrbp_1 _7100_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1045),
    .D(\vgademo.soundtrack.sigma_delta_accum_[1] ),
    .Q_N(_3564_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[1] ));
 sg13g2_dfrbp_1 _7101_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1045),
    .D(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .Q_N(_3565_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[2] ));
 sg13g2_dfrbp_1 _7102_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1056),
    .D(net533),
    .Q_N(_3566_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[3] ));
 sg13g2_dfrbp_1 _7103_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1056),
    .D(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .Q_N(_3567_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[4] ));
 sg13g2_dfrbp_1 _7104_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1056),
    .D(net520),
    .Q_N(_3568_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[5] ));
 sg13g2_dfrbp_1 _7105_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1056),
    .D(\vgademo.soundtrack.sigma_delta_accum_[6] ),
    .Q_N(_3569_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[6] ));
 sg13g2_dfrbp_1 _7106_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1056),
    .D(net517),
    .Q_N(_3570_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[7] ));
 sg13g2_dfrbp_1 _7107_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1056),
    .D(net512),
    .Q_N(_3571_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[8] ));
 sg13g2_dfrbp_1 _7108_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1057),
    .D(net502),
    .Q_N(_3572_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[9] ));
 sg13g2_dfrbp_1 _7109_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1057),
    .D(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .Q_N(_3573_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[10] ));
 sg13g2_dfrbp_1 _7110_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1057),
    .D(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .Q_N(_3574_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[11] ));
 sg13g2_dfrbp_1 _7111_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1047),
    .D(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .Q_N(_3575_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[12] ));
 sg13g2_dfrbp_1 _7112_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1047),
    .D(net514),
    .Q_N(_3576_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[13] ));
 sg13g2_dfrbp_1 _7113_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1047),
    .D(\vgademo.soundtrack.sigma_delta_accum_[14] ),
    .Q_N(_3577_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[14] ));
 sg13g2_dfrbp_1 _7114_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1048),
    .D(\vgademo.soundtrack.sigma_delta_accum_[15] ),
    .Q_N(_3541_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[15] ));
 sg13g2_dfrbp_1 _7115_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1047),
    .D(_0147_),
    .Q_N(_0058_),
    .Q(\vgademo.audio_beat_out[0] ));
 sg13g2_dfrbp_1 _7116_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1047),
    .D(net576),
    .Q_N(_0059_),
    .Q(\vgademo.audio_beat_out[1] ));
 sg13g2_dfrbp_1 _7117_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1046),
    .D(net510),
    .Q_N(_0062_),
    .Q(\vgademo.audio_beat_out[2] ));
 sg13g2_dfrbp_1 _7118_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1046),
    .D(net452),
    .Q_N(_0057_),
    .Q(\vgademo.audio_beat_out[3] ));
 sg13g2_dfrbp_1 _7119_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1046),
    .D(net493),
    .Q_N(_0055_),
    .Q(\vgademo.audio_beat_out[4] ));
 sg13g2_dfrbp_1 _7120_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1043),
    .D(_0152_),
    .Q_N(_3540_),
    .Q(\vgademo.soundtrack.tri_osc_i[0] ));
 sg13g2_dfrbp_1 _7121_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1043),
    .D(_0153_),
    .Q_N(_3539_),
    .Q(\vgademo.soundtrack.tri_osc_i[1] ));
 sg13g2_dfrbp_1 _7122_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1043),
    .D(_0154_),
    .Q_N(_3538_),
    .Q(\vgademo.soundtrack.tri_osc_i[2] ));
 sg13g2_dfrbp_1 _7123_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1043),
    .D(_0155_),
    .Q_N(_3537_),
    .Q(\vgademo.soundtrack.tri_osc_i[3] ));
 sg13g2_dfrbp_1 _7124_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1043),
    .D(_0156_),
    .Q_N(_3536_),
    .Q(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_dfrbp_1 _7125_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1045),
    .D(_0157_),
    .Q_N(_3535_),
    .Q(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_dfrbp_1 _7126_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1045),
    .D(_0158_),
    .Q_N(_3534_),
    .Q(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_dfrbp_1 _7127_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net1045),
    .D(_0159_),
    .Q_N(_3533_),
    .Q(\vgademo.soundtrack.tri_osc_i[7] ));
 sg13g2_dfrbp_1 _7128_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1045),
    .D(net522),
    .Q_N(_3532_),
    .Q(\vgademo.soundtrack.tri_osc_i[8] ));
 sg13g2_dfrbp_1 _7129_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net94),
    .D(net241),
    .Q_N(_3531_),
    .Q(audio));
 sg13g2_dfrbp_1 _7130_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1060),
    .D(net175),
    .Q_N(\vgademo.soundtrack.tick_div_[0] ),
    .Q(\vgademo.soundtrack.tick_div[0] ));
 sg13g2_dfrbp_1 _7131_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1060),
    .D(net498),
    .Q_N(_3530_),
    .Q(\vgademo.soundtrack.tick_div[1] ));
 sg13g2_dfrbp_1 _7132_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1061),
    .D(net243),
    .Q_N(_3529_),
    .Q(\vgademo.soundtrack.tick_div[2] ));
 sg13g2_dfrbp_1 _7133_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1061),
    .D(net251),
    .Q_N(_3528_),
    .Q(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_dfrbp_1 _7134_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1058),
    .D(net214),
    .Q_N(_3527_),
    .Q(\vgademo.soundtrack.tick_div[4] ));
 sg13g2_dfrbp_1 _7135_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1058),
    .D(_0167_),
    .Q_N(_3526_),
    .Q(\vgademo.soundtrack.tick_div[5] ));
 sg13g2_dfrbp_1 _7136_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1058),
    .D(net208),
    .Q_N(_3525_),
    .Q(\vgademo.soundtrack.tick_div[6] ));
 sg13g2_dfrbp_1 _7137_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1046),
    .D(_0169_),
    .Q_N(_3524_),
    .Q(\vgademo.soundtrack.tick_div[7] ));
 sg13g2_dfrbp_1 _7138_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1054),
    .D(net183),
    .Q_N(\vgademo.soundtrack.noise_lfsr[0] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 _7139_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1054),
    .D(net185),
    .Q_N(\vgademo.soundtrack.noise_lfsr[1] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 _7140_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1054),
    .D(net181),
    .Q_N(\vgademo.soundtrack.noise_lfsr[2] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 _7141_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1055),
    .D(net237),
    .Q_N(\vgademo.soundtrack.noise_lfsr[3] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 _7142_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1055),
    .D(net233),
    .Q_N(_0040_),
    .Q(\vgademo.soundtrack.noise_lfsr[4] ));
 sg13g2_dfrbp_1 _7143_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1054),
    .D(net171),
    .Q_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 _7144_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1054),
    .D(net292),
    .Q_N(_0084_),
    .Q(\vgademo.soundtrack.noise_lfsr[6] ));
 sg13g2_dfrbp_1 _7145_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1058),
    .D(net177),
    .Q_N(\vgademo.soundtrack.noise_lfsr[7] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 _7146_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1058),
    .D(net330),
    .Q_N(_0083_),
    .Q(\vgademo.soundtrack.noise_lfsr[8] ));
 sg13g2_dfrbp_1 _7147_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1054),
    .D(net197),
    .Q_N(_3523_),
    .Q(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_dfrbp_1 _7148_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1055),
    .D(net167),
    .Q_N(\vgademo.soundtrack.noise_lfsr[10] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _7149_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1055),
    .D(net195),
    .Q_N(\vgademo.soundtrack.noise_lfsr[11] ),
    .Q(_0101_));
 sg13g2_dfrbp_1 _7150_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1054),
    .D(net173),
    .Q_N(\vgademo.soundtrack.noise_lfsr[12] ),
    .Q(_0102_));
 sg13g2_dfrbp_1 _7151_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1065),
    .D(net226),
    .Q_N(_0082_),
    .Q(\vgademo.soundtrack.noise_lfsr[13] ));
 sg13g2_dfrbp_1 _7152_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1054),
    .D(net308),
    .Q_N(_3522_),
    .Q(\vgademo.soundtrack.noise_lfsr[14] ));
 sg13g2_dfrbp_1 _7153_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1057),
    .D(net262),
    .Q_N(\vgademo.audio_snare_frames[0] ),
    .Q(_0103_));
 sg13g2_dfrbp_1 _7154_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1057),
    .D(_0186_),
    .Q_N(\vgademo.audio_snare_frames[1] ),
    .Q(_0104_));
 sg13g2_dfrbp_1 _7155_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1057),
    .D(_0187_),
    .Q_N(\vgademo.audio_snare_frames[2] ),
    .Q(_0105_));
 sg13g2_dfrbp_1 _7156_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1057),
    .D(net217),
    .Q_N(\vgademo.audio_snare_frames[3] ),
    .Q(_0106_));
 sg13g2_dfrbp_1 _7157_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net64),
    .D(_0189_),
    .Q_N(_3521_),
    .Q(\vgademo.soundtrack.pulse_osc_p[0] ));
 sg13g2_dfrbp_1 _7158_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net63),
    .D(net191),
    .Q_N(_0042_),
    .Q(\vgademo.soundtrack.pulse_osc_p[1] ));
 sg13g2_dfrbp_1 _7159_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net62),
    .D(_0191_),
    .Q_N(_3520_),
    .Q(\vgademo.soundtrack.pulse_osc_p[2] ));
 sg13g2_dfrbp_1 _7160_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net61),
    .D(_0192_),
    .Q_N(_3519_),
    .Q(\vgademo.soundtrack.pulse_osc_p[3] ));
 sg13g2_dfrbp_1 _7161_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net60),
    .D(net343),
    .Q_N(_3518_),
    .Q(\vgademo.soundtrack.pulse_osc_p[4] ));
 sg13g2_dfrbp_1 _7162_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net59),
    .D(_0194_),
    .Q_N(_3517_),
    .Q(\vgademo.soundtrack.pulse_osc_p[5] ));
 sg13g2_dfrbp_1 _7163_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net58),
    .D(net289),
    .Q_N(_3516_),
    .Q(\vgademo.soundtrack.pulse_osc_p[6] ));
 sg13g2_dfrbp_1 _7164_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net57),
    .D(net363),
    .Q_N(_3515_),
    .Q(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_dfrbp_1 _7165_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net56),
    .D(_0197_),
    .Q_N(_3514_),
    .Q(\vgademo.soundtrack.pulse_osc_p[8] ));
 sg13g2_dfrbp_1 _7166_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net55),
    .D(net258),
    .Q_N(_3513_),
    .Q(\vgademo.soundtrack.pulse_osc_p[9] ));
 sg13g2_dfrbp_1 _7167_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net54),
    .D(net223),
    .Q_N(_3512_),
    .Q(\vgademo.soundtrack.pulse_osc_p[10] ));
 sg13g2_dfrbp_1 _7168_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net53),
    .D(_0200_),
    .Q_N(_3511_),
    .Q(\vgademo.soundtrack.pulse_osc_p[11] ));
 sg13g2_dfrbp_1 _7169_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net52),
    .D(_0201_),
    .Q_N(_3510_),
    .Q(\vgademo.soundtrack.pulse_osc_p[12] ));
 sg13g2_dfrbp_1 _7170_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net51),
    .D(net264),
    .Q_N(_3509_),
    .Q(\vgademo.soundtrack.pulse_osc_p[13] ));
 sg13g2_dfrbp_1 _7171_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1046),
    .D(net578),
    .Q_N(_3508_),
    .Q(\vgademo.audio_kick_frames[0] ));
 sg13g2_dfrbp_1 _7172_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1046),
    .D(_0204_),
    .Q_N(_0068_),
    .Q(\vgademo.audio_kick_frames[1] ));
 sg13g2_dfrbp_1 _7173_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1046),
    .D(_0205_),
    .Q_N(_0060_),
    .Q(\vgademo.audio_kick_frames[2] ));
 sg13g2_dfrbp_1 _7174_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1046),
    .D(net179),
    .Q_N(\vgademo.soundtrack.pulse_vol[0] ),
    .Q(_0107_));
 sg13g2_dfrbp_1 _7175_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1048),
    .D(_0207_),
    .Q_N(\vgademo.soundtrack.pulse_vol[1] ),
    .Q(_0108_));
 sg13g2_dfrbp_1 _7176_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1045),
    .D(net193),
    .Q_N(\vgademo.soundtrack.pulse_vol[2] ),
    .Q(_0109_));
 sg13g2_dfrbp_1 _7177_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1047),
    .D(net199),
    .Q_N(\vgademo.soundtrack.pulse_vol[3] ),
    .Q(_0110_));
 sg13g2_dfrbp_1 _7178_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1061),
    .D(net165),
    .Q_N(\vgademo.soundtrack.sample_div_[0] ),
    .Q(\vgademo.soundtrack.sample_div[0] ));
 sg13g2_dfrbp_1 _7179_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1062),
    .D(net255),
    .Q_N(_3578_),
    .Q(\vgademo.soundtrack.sample_div[1] ));
 sg13g2_dfrbp_1 _7180_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1061),
    .D(net455),
    .Q_N(_3579_),
    .Q(\vgademo.soundtrack.sample_div[2] ));
 sg13g2_dfrbp_1 _7181_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1060),
    .D(net245),
    .Q_N(_3580_),
    .Q(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_dfrbp_1 _7182_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1060),
    .D(net229),
    .Q_N(_3581_),
    .Q(\vgademo.soundtrack.sample_div[4] ));
 sg13g2_dfrbp_1 _7183_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1060),
    .D(\vgademo.soundtrack.sample_div_[5] ),
    .Q_N(_3582_),
    .Q(\vgademo.soundtrack.sample_div[5] ));
 sg13g2_dfrbp_1 _7184_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1060),
    .D(\vgademo.soundtrack.sample_div_[6] ),
    .Q_N(_3583_),
    .Q(\vgademo.soundtrack.sample_div[6] ));
 sg13g2_dfrbp_1 _7185_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1065),
    .D(net231),
    .Q_N(_3584_),
    .Q(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_dfrbp_1 _7186_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1060),
    .D(net212),
    .Q_N(_3585_),
    .Q(\vgademo.soundtrack.sample_div[8] ));
 sg13g2_dfrbp_1 _7187_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1060),
    .D(net269),
    .Q_N(_3507_),
    .Q(\vgademo.soundtrack.sample_div[9] ));
 sg13g2_dfrbp_1 _7188_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net42),
    .D(net260),
    .Q_N(_3506_),
    .Q(\vgademo.soundtrack.tri_osc_p[0] ));
 sg13g2_dfrbp_1 _7189_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net41),
    .D(_0211_),
    .Q_N(_3505_),
    .Q(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_dfrbp_1 _7190_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net40),
    .D(_0212_),
    .Q_N(_3504_),
    .Q(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_dfrbp_1 _7191_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net39),
    .D(_0213_),
    .Q_N(_3503_),
    .Q(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_dfrbp_1 _7192_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net38),
    .D(_0214_),
    .Q_N(_3502_),
    .Q(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_dfrbp_1 _7193_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net37),
    .D(_0215_),
    .Q_N(_3501_),
    .Q(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_dfrbp_1 _7194_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net36),
    .D(net471),
    .Q_N(_3500_),
    .Q(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_dfrbp_1 _7195_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net35),
    .D(net429),
    .Q_N(_3499_),
    .Q(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_dfrbp_1 _7196_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net34),
    .D(net421),
    .Q_N(_3498_),
    .Q(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_dfrbp_1 _7197_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net33),
    .D(net387),
    .Q_N(_0041_),
    .Q(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_dfrbp_1 _7198_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net32),
    .D(net282),
    .Q_N(_3497_),
    .Q(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_dfrbp_1 _7199_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net31),
    .D(_0221_),
    .Q_N(_3496_),
    .Q(\vgademo.soundtrack.tri_osc_p[11] ));
 sg13g2_dfrbp_1 _7200_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net30),
    .D(_0222_),
    .Q_N(_3495_),
    .Q(\vgademo.soundtrack.tri_osc_p[12] ));
 sg13g2_dfrbp_1 _7201_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net29),
    .D(net347),
    .Q_N(_3494_),
    .Q(\vgademo.soundtrack.tri_osc_p[13] ));
 sg13g2_dfrbp_1 _7202_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net28),
    .D(net369),
    .Q_N(_3493_),
    .Q(\vgademo.soundtrack.tri_osc_p[14] ));
 sg13g2_dfrbp_1 _7203_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net27),
    .D(_0225_),
    .Q_N(_3492_),
    .Q(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_dfrbp_1 _7204_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net24),
    .D(_0226_),
    .Q_N(_3491_),
    .Q(\vgademo.plane_dx_div.d[16] ));
 sg13g2_dfrbp_1 _7205_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net23),
    .D(_0227_),
    .Q_N(_0070_),
    .Q(\vgademo.plane_dx_div.d[17] ));
 sg13g2_dfrbp_1 _7206_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net22),
    .D(_0228_),
    .Q_N(_0073_),
    .Q(\vgademo.plane_dx_div.d[18] ));
 sg13g2_dfrbp_1 _7207_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net21),
    .D(_0229_),
    .Q_N(_0076_),
    .Q(\vgademo.plane_dx_div.d[19] ));
 sg13g2_dfrbp_1 _7208_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net20),
    .D(_0230_),
    .Q_N(_0079_),
    .Q(\vgademo.plane_dx_div.d[20] ));
 sg13g2_dfrbp_1 _7209_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net19),
    .D(_0231_),
    .Q_N(_0081_),
    .Q(\vgademo.plane_dx_div.d[21] ));
 sg13g2_dfrbp_1 _7210_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net18),
    .D(_0232_),
    .Q_N(_0013_),
    .Q(\vgademo.plane_dx_div.d[22] ));
 sg13g2_dfrbp_1 _7211_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net17),
    .D(_0233_),
    .Q_N(_0017_),
    .Q(\vgademo.plane_dx_div.d[23] ));
 sg13g2_dfrbp_1 _7212_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net90),
    .D(_0234_),
    .Q_N(_0020_),
    .Q(\vgademo.plane_dx_div.d[24] ));
 sg13g2_dfrbp_1 _7213_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net91),
    .D(_0012_),
    .Q_N(_3586_),
    .Q(\vgademo.vsync ));
 sg13g2_dfrbp_1 _7214_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net92),
    .D(_0011_),
    .Q_N(_3587_),
    .Q(hsync));
 sg13g2_dfrbp_1 _7215_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1059),
    .D(net556),
    .Q_N(_3588_),
    .Q(\vgademo.h_count[0] ));
 sg13g2_dfrbp_1 _7216_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1059),
    .D(_0002_),
    .Q_N(_3589_),
    .Q(\vgademo.h_count[1] ));
 sg13g2_dfrbp_1 _7217_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1047),
    .D(_0003_),
    .Q_N(_0033_),
    .Q(\vgademo.h_count[2] ));
 sg13g2_dfrbp_1 _7218_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1051),
    .D(net461),
    .Q_N(_0034_),
    .Q(\vgademo.h_count[3] ));
 sg13g2_dfrbp_1 _7219_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1051),
    .D(_0005_),
    .Q_N(_0044_),
    .Q(\vgademo.h_count[4] ));
 sg13g2_dfrbp_1 _7220_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1051),
    .D(_0006_),
    .Q_N(_0035_),
    .Q(\vgademo.h_count[5] ));
 sg13g2_dfrbp_1 _7221_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1066),
    .D(net553),
    .Q_N(_0036_),
    .Q(\vgademo.h_count[6] ));
 sg13g2_dfrbp_1 _7222_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1066),
    .D(_0008_),
    .Q_N(_0037_),
    .Q(\vgademo.h_count[7] ));
 sg13g2_dfrbp_1 _7223_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1051),
    .D(_0009_),
    .Q_N(_0038_),
    .Q(\vgademo.h_count[8] ));
 sg13g2_dfrbp_1 _7224_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1051),
    .D(net235),
    .Q_N(_0039_),
    .Q(\vgademo.h_count[9] ));
 sg13g2_dfrbp_1 _7225_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1051),
    .D(net274),
    .Q_N(_0061_),
    .Q(\vgademo.h_count[10] ));
 sg13g2_dfrbp_1 _7226_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1049),
    .D(_0235_),
    .Q_N(_0064_),
    .Q(\vgademo.a_scrolly[3] ));
 sg13g2_dfrbp_1 _7227_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1049),
    .D(_0236_),
    .Q_N(_0069_),
    .Q(\vgademo.a_scrolly[4] ));
 sg13g2_dfrbp_1 _7228_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net1049),
    .D(_0237_),
    .Q_N(_0056_),
    .Q(\vgademo.a_scrolly[5] ));
 sg13g2_dfrbp_1 _7229_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1049),
    .D(_0238_),
    .Q_N(_0075_),
    .Q(\vgademo.a_scrolly[6] ));
 sg13g2_dfrbp_1 _7230_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1050),
    .D(_0239_),
    .Q_N(_0078_),
    .Q(\vgademo.a_scrolly[7] ));
 sg13g2_dfrbp_1 _7231_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1049),
    .D(net573),
    .Q_N(_0080_),
    .Q(\vgademo.a_scrolly[8] ));
 sg13g2_dfrbp_1 _7232_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1049),
    .D(net504),
    .Q_N(_0065_),
    .Q(\vgademo.a_scrolly[9] ));
 sg13g2_dfrbp_1 _7233_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1049),
    .D(net424),
    .Q_N(_0015_),
    .Q(\vgademo.a_scrolly[10] ));
 sg13g2_dfrbp_1 _7234_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1050),
    .D(net239),
    .Q_N(_0019_),
    .Q(\vgademo.a_scrolly[11] ));
 sg13g2_dfrbp_1 _7235_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1050),
    .D(net537),
    .Q_N(_0067_),
    .Q(\vgademo.a_scrolly[12] ));
 sg13g2_dfrbp_1 _7236_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1050),
    .D(net404),
    .Q_N(_0066_),
    .Q(\vgademo.a_scrolly[13] ));
 sg13g2_dfrbp_1 _7237_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1066),
    .D(_0246_),
    .Q_N(_3490_),
    .Q(\vgademo.bayer_j[0] ));
 sg13g2_dfrbp_1 _7238_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1066),
    .D(_0247_),
    .Q_N(_0072_),
    .Q(\vgademo.bayer_j[1] ));
 sg13g2_dfrbp_1 _7239_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1066),
    .D(net463),
    .Q_N(_0071_),
    .Q(\vgademo.v_count[2] ));
 sg13g2_dfrbp_1 _7240_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1066),
    .D(net543),
    .Q_N(_0074_),
    .Q(\vgademo.v_count[3] ));
 sg13g2_dfrbp_1 _7241_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1051),
    .D(net266),
    .Q_N(_0077_),
    .Q(\vgademo.v_count[4] ));
 sg13g2_dfrbp_1 _7242_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1066),
    .D(net306),
    .Q_N(_0063_),
    .Q(\vgademo.v_count[5] ));
 sg13g2_dfrbp_1 _7243_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1052),
    .D(net535),
    .Q_N(_0016_),
    .Q(\vgademo.v_count[6] ));
 sg13g2_dfrbp_1 _7244_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1052),
    .D(net478),
    .Q_N(_0014_),
    .Q(\vgademo.v_count[7] ));
 sg13g2_dfrbp_1 _7245_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1052),
    .D(net531),
    .Q_N(_0018_),
    .Q(\vgademo.v_count[8] ));
 sg13g2_dfrbp_1 _7246_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1052),
    .D(_0255_),
    .Q_N(_0021_),
    .Q(\vgademo.v_count[9] ));
 sg13g2_dfrbp_1 _7247_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net16),
    .D(_0256_),
    .Q_N(_3489_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7248_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net15),
    .D(_0257_),
    .Q_N(_3488_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7249_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1061),
    .D(net253),
    .Q_N(_3487_),
    .Q(\vgademo.a_cos[0] ));
 sg13g2_dfrbp_1 _7250_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1063),
    .D(_0259_),
    .Q_N(_3486_),
    .Q(\vgademo.a_cos[1] ));
 sg13g2_dfrbp_1 _7251_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1063),
    .D(_0260_),
    .Q_N(_3485_),
    .Q(\vgademo.a_cos[2] ));
 sg13g2_dfrbp_1 _7252_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1063),
    .D(_0261_),
    .Q_N(_3484_),
    .Q(\vgademo.a_cos[3] ));
 sg13g2_dfrbp_1 _7253_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1067),
    .D(_0262_),
    .Q_N(_3483_),
    .Q(\vgademo.a_cos[4] ));
 sg13g2_dfrbp_1 _7254_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1067),
    .D(_0263_),
    .Q_N(_3482_),
    .Q(\vgademo.a_cos[5] ));
 sg13g2_dfrbp_1 _7255_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1063),
    .D(_0264_),
    .Q_N(_3481_),
    .Q(\vgademo.a_cos[6] ));
 sg13g2_dfrbp_1 _7256_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1062),
    .D(_0265_),
    .Q_N(_3480_),
    .Q(\vgademo.a_cos[7] ));
 sg13g2_dfrbp_1 _7257_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1062),
    .D(_0266_),
    .Q_N(_3479_),
    .Q(\vgademo.a_cos[8] ));
 sg13g2_dfrbp_1 _7258_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1062),
    .D(_0267_),
    .Q_N(_3478_),
    .Q(\vgademo.a_cos[9] ));
 sg13g2_dfrbp_1 _7259_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1059),
    .D(_0268_),
    .Q_N(_3477_),
    .Q(\vgademo.a_cos[10] ));
 sg13g2_dfrbp_1 _7260_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1059),
    .D(_0269_),
    .Q_N(_3476_),
    .Q(\vgademo.a_cos[11] ));
 sg13g2_dfrbp_1 _7261_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1059),
    .D(_0270_),
    .Q_N(_3475_),
    .Q(\vgademo.a_cos[12] ));
 sg13g2_dfrbp_1 _7262_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1059),
    .D(_0271_),
    .Q_N(\vgademo.a_cos[13] ),
    .Q(_0111_));
 sg13g2_dfrbp_1 _7263_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1057),
    .D(_0272_),
    .Q_N(_3474_),
    .Q(\vgademo.a_cos[14] ));
 sg13g2_dfrbp_1 _7264_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1063),
    .D(_0273_),
    .Q_N(_3473_),
    .Q(\vgademo.a_sin[0] ));
 sg13g2_dfrbp_1 _7265_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1061),
    .D(_0274_),
    .Q_N(_3472_),
    .Q(\vgademo.a_sin[1] ));
 sg13g2_dfrbp_1 _7266_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1061),
    .D(net301),
    .Q_N(_3471_),
    .Q(\vgademo.a_sin[2] ));
 sg13g2_dfrbp_1 _7267_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1058),
    .D(_0276_),
    .Q_N(_3470_),
    .Q(\vgademo.a_sin[3] ));
 sg13g2_dfrbp_1 _7268_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1058),
    .D(net367),
    .Q_N(_3469_),
    .Q(\vgademo.a_sin[4] ));
 sg13g2_dfrbp_1 _7269_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1058),
    .D(_0278_),
    .Q_N(_3468_),
    .Q(\vgademo.a_sin[5] ));
 sg13g2_dfrbp_1 _7270_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1061),
    .D(net480),
    .Q_N(_3467_),
    .Q(\vgademo.a_sin[6] ));
 sg13g2_dfrbp_1 _7271_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1062),
    .D(_0280_),
    .Q_N(_3466_),
    .Q(\vgademo.a_sin[7] ));
 sg13g2_dfrbp_1 _7272_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1064),
    .D(_0281_),
    .Q_N(_3465_),
    .Q(\vgademo.a_sin[8] ));
 sg13g2_dfrbp_1 _7273_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1064),
    .D(_0282_),
    .Q_N(_3464_),
    .Q(\vgademo.a_sin[9] ));
 sg13g2_dfrbp_1 _7274_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1063),
    .D(_0283_),
    .Q_N(_3463_),
    .Q(\vgademo.a_sin[10] ));
 sg13g2_dfrbp_1 _7275_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1063),
    .D(_0284_),
    .Q_N(_3462_),
    .Q(\vgademo.a_sin[11] ));
 sg13g2_dfrbp_1 _7276_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1063),
    .D(_0285_),
    .Q_N(_3461_),
    .Q(\vgademo.a_sin[12] ));
 sg13g2_dfrbp_1 _7277_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1062),
    .D(_0286_),
    .Q_N(_3460_),
    .Q(\vgademo.a_sin[13] ));
 sg13g2_dfrbp_1 _7278_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1062),
    .D(_0287_),
    .Q_N(_3459_),
    .Q(\vgademo.a_sin[14] ));
 sg13g2_dfrbp_1 _7279_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net162),
    .D(_0288_),
    .Q_N(_3458_),
    .Q(\vgademo.scanline_audio_sample[0] ));
 sg13g2_dfrbp_1 _7280_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net160),
    .D(_0289_),
    .Q_N(_3457_),
    .Q(\vgademo.scanline_audio_sample[1] ));
 sg13g2_dfrbp_1 _7281_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net158),
    .D(_0290_),
    .Q_N(_3456_),
    .Q(\vgademo.scanline_audio_sample[2] ));
 sg13g2_dfrbp_1 _7282_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net156),
    .D(_0291_),
    .Q_N(_3455_),
    .Q(\vgademo.scanline_audio_sample[3] ));
 sg13g2_dfrbp_1 _7283_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net154),
    .D(_0292_),
    .Q_N(_3454_),
    .Q(\vgademo.scanline_audio_sample[4] ));
 sg13g2_dfrbp_1 _7284_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net152),
    .D(_0293_),
    .Q_N(_0043_),
    .Q(\vgademo.scanline_audio_sample[5] ));
 sg13g2_dfrbp_1 _7285_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net150),
    .D(_0294_),
    .Q_N(_3453_),
    .Q(\vgademo.scanline_audio_sample[6] ));
 sg13g2_dfrbp_1 _7286_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net148),
    .D(net287),
    .Q_N(_3452_),
    .Q(\vgademo.b_cos[0] ));
 sg13g2_dfrbp_1 _7287_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net146),
    .D(net336),
    .Q_N(_3451_),
    .Q(\vgademo.b_cos[1] ));
 sg13g2_dfrbp_1 _7288_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net144),
    .D(_0297_),
    .Q_N(_3450_),
    .Q(\vgademo.b_cos[2] ));
 sg13g2_dfrbp_1 _7289_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net142),
    .D(net345),
    .Q_N(_3449_),
    .Q(\vgademo.b_cos[3] ));
 sg13g2_dfrbp_1 _7290_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net140),
    .D(net444),
    .Q_N(_3448_),
    .Q(\vgademo.b_cos[4] ));
 sg13g2_dfrbp_1 _7291_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net138),
    .D(_0300_),
    .Q_N(_3447_),
    .Q(\vgademo.b_cos[5] ));
 sg13g2_dfrbp_1 _7292_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net137),
    .D(_0301_),
    .Q_N(_3446_),
    .Q(\vgademo.b_cos[6] ));
 sg13g2_dfrbp_1 _7293_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net136),
    .D(net484),
    .Q_N(_3445_),
    .Q(\vgademo.b_cos[7] ));
 sg13g2_dfrbp_1 _7294_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net135),
    .D(net439),
    .Q_N(_3444_),
    .Q(\vgademo.b_cos[8] ));
 sg13g2_dfrbp_1 _7295_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net134),
    .D(_0304_),
    .Q_N(_3443_),
    .Q(\vgademo.b_cos[9] ));
 sg13g2_dfrbp_1 _7296_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net133),
    .D(net411),
    .Q_N(_3442_),
    .Q(\vgademo.b_cos[10] ));
 sg13g2_dfrbp_1 _7297_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net132),
    .D(_0306_),
    .Q_N(_3441_),
    .Q(\vgademo.b_cos[11] ));
 sg13g2_dfrbp_1 _7298_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net131),
    .D(net350),
    .Q_N(_3440_),
    .Q(\vgademo.plane_dx_div.r[16] ));
 sg13g2_dfrbp_1 _7299_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net130),
    .D(_0308_),
    .Q_N(_3439_),
    .Q(\vgademo.plane_dx_div.r[17] ));
 sg13g2_dfrbp_1 _7300_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net129),
    .D(net334),
    .Q_N(_3438_),
    .Q(\vgademo.plane_dx_div.r[18] ));
 sg13g2_dfrbp_1 _7301_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net128),
    .D(net341),
    .Q_N(_3437_),
    .Q(\vgademo.plane_dx_div.r[19] ));
 sg13g2_dfrbp_1 _7302_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net127),
    .D(_0311_),
    .Q_N(_3436_),
    .Q(\vgademo.plane_dx_div.r[20] ));
 sg13g2_dfrbp_1 _7303_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net126),
    .D(_0312_),
    .Q_N(_3435_),
    .Q(\vgademo.plane_dx_div.r[21] ));
 sg13g2_dfrbp_1 _7304_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net125),
    .D(_0313_),
    .Q_N(_3434_),
    .Q(\vgademo.plane_dx_div.r[22] ));
 sg13g2_dfrbp_1 _7305_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net124),
    .D(_0314_),
    .Q_N(_3433_),
    .Q(\vgademo.plane_dx_div.r[23] ));
 sg13g2_dfrbp_1 _7306_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net123),
    .D(_0315_),
    .Q_N(_3432_),
    .Q(\vgademo.plane_dx_div.r[24] ));
 sg13g2_dfrbp_1 _7307_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net122),
    .D(_0316_),
    .Q_N(\vgademo.plane_dx[0] ),
    .Q(\vgademo.plane_dx_div.r[25] ));
 sg13g2_dfrbp_1 _7308_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net120),
    .D(_0317_),
    .Q_N(_3431_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7309_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net118),
    .D(_0318_),
    .Q_N(_3430_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7310_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net116),
    .D(_0319_),
    .Q_N(_3429_),
    .Q(\vgademo.b_sin[0] ));
 sg13g2_dfrbp_1 _7311_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net114),
    .D(net379),
    .Q_N(_3428_),
    .Q(\vgademo.b_sin[1] ));
 sg13g2_dfrbp_1 _7312_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net112),
    .D(_0321_),
    .Q_N(_3427_),
    .Q(\vgademo.b_sin[2] ));
 sg13g2_dfrbp_1 _7313_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net110),
    .D(_0322_),
    .Q_N(_3426_),
    .Q(\vgademo.b_sin[3] ));
 sg13g2_dfrbp_1 _7314_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net108),
    .D(_0323_),
    .Q_N(_3425_),
    .Q(\vgademo.b_sin[4] ));
 sg13g2_dfrbp_1 _7315_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net106),
    .D(net299),
    .Q_N(_3424_),
    .Q(\vgademo.b_sin[5] ));
 sg13g2_dfrbp_1 _7316_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net104),
    .D(_0325_),
    .Q_N(_3423_),
    .Q(\vgademo.b_sin[6] ));
 sg13g2_dfrbp_1 _7317_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net102),
    .D(net359),
    .Q_N(_3422_),
    .Q(\vgademo.b_sin[7] ));
 sg13g2_dfrbp_1 _7318_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net100),
    .D(_0327_),
    .Q_N(_3421_),
    .Q(\vgademo.b_sin[8] ));
 sg13g2_dfrbp_1 _7319_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net98),
    .D(net437),
    .Q_N(_3420_),
    .Q(\vgademo.b_sin[9] ));
 sg13g2_dfrbp_1 _7320_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net96),
    .D(_0329_),
    .Q_N(_3419_),
    .Q(\vgademo.b_sin[10] ));
 sg13g2_dfrbp_1 _7321_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net95),
    .D(net551),
    .Q_N(_3418_),
    .Q(\vgademo.b_sin[11] ));
 sg13g2_dfrbp_1 _7322_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net93),
    .D(net284),
    .Q_N(_3417_),
    .Q(\vgademo.plane_u[1] ));
 sg13g2_dfrbp_1 _7323_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net89),
    .D(_0332_),
    .Q_N(_3416_),
    .Q(\vgademo.plane_u[2] ));
 sg13g2_dfrbp_1 _7324_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net88),
    .D(_0333_),
    .Q_N(_3415_),
    .Q(\vgademo.plane_u[3] ));
 sg13g2_dfrbp_1 _7325_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net87),
    .D(_0334_),
    .Q_N(_3414_),
    .Q(\vgademo.plane_u[4] ));
 sg13g2_dfrbp_1 _7326_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net86),
    .D(_0335_),
    .Q_N(_3413_),
    .Q(\vgademo.plane_u[5] ));
 sg13g2_dfrbp_1 _7327_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net85),
    .D(_0336_),
    .Q_N(_3412_),
    .Q(\vgademo.plane_u[6] ));
 sg13g2_dfrbp_1 _7328_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net84),
    .D(_0337_),
    .Q_N(_3411_),
    .Q(\vgademo.plane_u[7] ));
 sg13g2_dfrbp_1 _7329_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net83),
    .D(_0338_),
    .Q_N(_3410_),
    .Q(\vgademo.plane_u[8] ));
 sg13g2_dfrbp_1 _7330_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net82),
    .D(_0339_),
    .Q_N(_3409_),
    .Q(\vgademo.plane_u[9] ));
 sg13g2_dfrbp_1 _7331_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net81),
    .D(_0340_),
    .Q_N(_3408_),
    .Q(\vgademo.plane_u[10] ));
 sg13g2_dfrbp_1 _7332_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net80),
    .D(net297),
    .Q_N(_0027_),
    .Q(\vgademo.plane_u[11] ));
 sg13g2_dfrbp_1 _7333_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net79),
    .D(net361),
    .Q_N(_0028_),
    .Q(\vgademo.plane_u[12] ));
 sg13g2_dfrbp_1 _7334_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net78),
    .D(net382),
    .Q_N(_0048_),
    .Q(\vgademo.plane_u[13] ));
 sg13g2_dfrbp_1 _7335_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net77),
    .D(_0344_),
    .Q_N(_0029_),
    .Q(\vgademo.plane_u[14] ));
 sg13g2_dfrbp_1 _7336_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net76),
    .D(_0345_),
    .Q_N(_0047_),
    .Q(\vgademo.plane_u[15] ));
 sg13g2_dfrbp_1 _7337_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net75),
    .D(_0346_),
    .Q_N(_0030_),
    .Q(\vgademo.plane_u[16] ));
 sg13g2_dfrbp_1 _7338_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net74),
    .D(_0347_),
    .Q_N(_0046_),
    .Q(\vgademo.plane_u[17] ));
 sg13g2_dfrbp_1 _7339_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net73),
    .D(_0348_),
    .Q_N(_0031_),
    .Q(\vgademo.plane_u[18] ));
 sg13g2_dfrbp_1 _7340_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net72),
    .D(net446),
    .Q_N(_0045_),
    .Q(\vgademo.plane_u[19] ));
 sg13g2_dfrbp_1 _7341_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net71),
    .D(_0350_),
    .Q_N(_0032_),
    .Q(\vgademo.plane_u[20] ));
 sg13g2_dfrbp_1 _7342_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net70),
    .D(net400),
    .Q_N(_3407_),
    .Q(\vgademo.plane_u[21] ));
 sg13g2_dfrbp_1 _7343_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net69),
    .D(_0352_),
    .Q_N(_3406_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7344_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net68),
    .D(_0353_),
    .Q_N(_3405_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7345_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net67),
    .D(net317),
    .Q_N(_3404_),
    .Q(\vgademo.plane_du[0] ));
 sg13g2_dfrbp_1 _7346_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net66),
    .D(net311),
    .Q_N(_3403_),
    .Q(\vgademo.plane_du[1] ));
 sg13g2_dfrbp_1 _7347_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net65),
    .D(net474),
    .Q_N(_3402_),
    .Q(\vgademo.plane_du[2] ));
 sg13g2_dfrbp_1 _7348_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net50),
    .D(_0357_),
    .Q_N(_0050_),
    .Q(\vgademo.plane_du[3] ));
 sg13g2_dfrbp_1 _7349_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net49),
    .D(net500),
    .Q_N(_0049_),
    .Q(\vgademo.plane_du[4] ));
 sg13g2_dfrbp_1 _7350_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net48),
    .D(_0359_),
    .Q_N(_0051_),
    .Q(\vgademo.plane_du[5] ));
 sg13g2_dfrbp_1 _7351_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net47),
    .D(_0360_),
    .Q_N(_0052_),
    .Q(\vgademo.plane_du[6] ));
 sg13g2_dfrbp_1 _7352_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net46),
    .D(_0361_),
    .Q_N(_0053_),
    .Q(\vgademo.plane_du[7] ));
 sg13g2_dfrbp_1 _7353_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net45),
    .D(net568),
    .Q_N(_0054_),
    .Q(\vgademo.plane_du[8] ));
 sg13g2_dfrbp_1 _7354_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net44),
    .D(_0363_),
    .Q_N(_3401_),
    .Q(\vgademo.plane_du[9] ));
 sg13g2_dfrbp_1 _7355_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net43),
    .D(net482),
    .Q_N(_3400_),
    .Q(\vgademo.plane_du[10] ));
 sg13g2_dfrbp_1 _7356_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net163),
    .D(net221),
    .Q_N(_3399_),
    .Q(\vgademo.plane_u[0] ));
 sg13g2_tiehi _7247__16 (.L_HI(net16));
 sg13g2_tiehi _7211__17 (.L_HI(net17));
 sg13g2_tiehi _7210__18 (.L_HI(net18));
 sg13g2_tiehi _7209__19 (.L_HI(net19));
 sg13g2_tiehi _7208__20 (.L_HI(net20));
 sg13g2_tiehi _7207__21 (.L_HI(net21));
 sg13g2_tiehi _7206__22 (.L_HI(net22));
 sg13g2_tiehi _7205__23 (.L_HI(net23));
 sg13g2_tiehi _7204__24 (.L_HI(net24));
 sg13g2_tiehi _7064__25 (.L_HI(net25));
 sg13g2_tiehi _7098__26 (.L_HI(net26));
 sg13g2_tiehi _7203__27 (.L_HI(net27));
 sg13g2_tiehi _7202__28 (.L_HI(net28));
 sg13g2_tiehi _7201__29 (.L_HI(net29));
 sg13g2_tiehi _7200__30 (.L_HI(net30));
 sg13g2_tiehi _7199__31 (.L_HI(net31));
 sg13g2_tiehi _7198__32 (.L_HI(net32));
 sg13g2_tiehi _7197__33 (.L_HI(net33));
 sg13g2_tiehi _7196__34 (.L_HI(net34));
 sg13g2_tiehi _7195__35 (.L_HI(net35));
 sg13g2_tiehi _7194__36 (.L_HI(net36));
 sg13g2_tiehi _7193__37 (.L_HI(net37));
 sg13g2_tiehi _7192__38 (.L_HI(net38));
 sg13g2_tiehi _7191__39 (.L_HI(net39));
 sg13g2_tiehi _7190__40 (.L_HI(net40));
 sg13g2_tiehi _7189__41 (.L_HI(net41));
 sg13g2_tiehi _7188__42 (.L_HI(net42));
 sg13g2_tiehi _7355__43 (.L_HI(net43));
 sg13g2_tiehi _7354__44 (.L_HI(net44));
 sg13g2_tiehi _7353__45 (.L_HI(net45));
 sg13g2_tiehi _7352__46 (.L_HI(net46));
 sg13g2_tiehi _7351__47 (.L_HI(net47));
 sg13g2_tiehi _7350__48 (.L_HI(net48));
 sg13g2_tiehi _7349__49 (.L_HI(net49));
 sg13g2_tiehi _7348__50 (.L_HI(net50));
 sg13g2_tiehi _7170__51 (.L_HI(net51));
 sg13g2_tiehi _7169__52 (.L_HI(net52));
 sg13g2_tiehi _7168__53 (.L_HI(net53));
 sg13g2_tiehi _7167__54 (.L_HI(net54));
 sg13g2_tiehi _7166__55 (.L_HI(net55));
 sg13g2_tiehi _7165__56 (.L_HI(net56));
 sg13g2_tiehi _7164__57 (.L_HI(net57));
 sg13g2_tiehi _7163__58 (.L_HI(net58));
 sg13g2_tiehi _7162__59 (.L_HI(net59));
 sg13g2_tiehi _7161__60 (.L_HI(net60));
 sg13g2_tiehi _7160__61 (.L_HI(net61));
 sg13g2_tiehi _7159__62 (.L_HI(net62));
 sg13g2_tiehi _7158__63 (.L_HI(net63));
 sg13g2_tiehi _7157__64 (.L_HI(net64));
 sg13g2_tiehi _7347__65 (.L_HI(net65));
 sg13g2_tiehi _7346__66 (.L_HI(net66));
 sg13g2_tiehi _7345__67 (.L_HI(net67));
 sg13g2_tiehi _7344__68 (.L_HI(net68));
 sg13g2_tiehi _7343__69 (.L_HI(net69));
 sg13g2_tiehi _7342__70 (.L_HI(net70));
 sg13g2_tiehi _7341__71 (.L_HI(net71));
 sg13g2_tiehi _7340__72 (.L_HI(net72));
 sg13g2_tiehi _7339__73 (.L_HI(net73));
 sg13g2_tiehi _7338__74 (.L_HI(net74));
 sg13g2_tiehi _7337__75 (.L_HI(net75));
 sg13g2_tiehi _7336__76 (.L_HI(net76));
 sg13g2_tiehi _7335__77 (.L_HI(net77));
 sg13g2_tiehi _7334__78 (.L_HI(net78));
 sg13g2_tiehi _7333__79 (.L_HI(net79));
 sg13g2_tiehi _7332__80 (.L_HI(net80));
 sg13g2_tiehi _7331__81 (.L_HI(net81));
 sg13g2_tiehi _7330__82 (.L_HI(net82));
 sg13g2_tiehi _7329__83 (.L_HI(net83));
 sg13g2_tiehi _7328__84 (.L_HI(net84));
 sg13g2_tiehi _7327__85 (.L_HI(net85));
 sg13g2_tiehi _7326__86 (.L_HI(net86));
 sg13g2_tiehi _7325__87 (.L_HI(net87));
 sg13g2_tiehi _7324__88 (.L_HI(net88));
 sg13g2_tiehi _7323__89 (.L_HI(net89));
 sg13g2_tiehi _7212__90 (.L_HI(net90));
 sg13g2_tiehi _7213__91 (.L_HI(net91));
 sg13g2_tiehi _7214__92 (.L_HI(net92));
 sg13g2_tiehi _7322__93 (.L_HI(net93));
 sg13g2_tiehi _7129__94 (.L_HI(net94));
 sg13g2_tiehi _7321__95 (.L_HI(net95));
 sg13g2_tiehi _7320__96 (.L_HI(net96));
 sg13g2_tiehi _7097__97 (.L_HI(net97));
 sg13g2_tiehi _7319__98 (.L_HI(net98));
 sg13g2_tiehi _7096__99 (.L_HI(net99));
 sg13g2_tiehi _7318__100 (.L_HI(net100));
 sg13g2_tiehi _7095__101 (.L_HI(net101));
 sg13g2_tiehi _7317__102 (.L_HI(net102));
 sg13g2_tiehi _7094__103 (.L_HI(net103));
 sg13g2_tiehi _7316__104 (.L_HI(net104));
 sg13g2_tiehi _7093__105 (.L_HI(net105));
 sg13g2_tiehi _7315__106 (.L_HI(net106));
 sg13g2_tiehi _7092__107 (.L_HI(net107));
 sg13g2_tiehi _7314__108 (.L_HI(net108));
 sg13g2_tiehi _7091__109 (.L_HI(net109));
 sg13g2_tiehi _7313__110 (.L_HI(net110));
 sg13g2_tiehi _7090__111 (.L_HI(net111));
 sg13g2_tiehi _7312__112 (.L_HI(net112));
 sg13g2_tiehi _7089__113 (.L_HI(net113));
 sg13g2_tiehi _7311__114 (.L_HI(net114));
 sg13g2_tiehi _7088__115 (.L_HI(net115));
 sg13g2_tiehi _7310__116 (.L_HI(net116));
 sg13g2_tiehi _7087__117 (.L_HI(net117));
 sg13g2_tiehi _7309__118 (.L_HI(net118));
 sg13g2_tiehi _7086__119 (.L_HI(net119));
 sg13g2_tiehi _7308__120 (.L_HI(net120));
 sg13g2_tiehi _7085__121 (.L_HI(net121));
 sg13g2_tiehi _7307__122 (.L_HI(net122));
 sg13g2_tiehi _7306__123 (.L_HI(net123));
 sg13g2_tiehi _7305__124 (.L_HI(net124));
 sg13g2_tiehi _7304__125 (.L_HI(net125));
 sg13g2_tiehi _7303__126 (.L_HI(net126));
 sg13g2_tiehi _7302__127 (.L_HI(net127));
 sg13g2_tiehi _7301__128 (.L_HI(net128));
 sg13g2_tiehi _7300__129 (.L_HI(net129));
 sg13g2_tiehi _7299__130 (.L_HI(net130));
 sg13g2_tiehi _7298__131 (.L_HI(net131));
 sg13g2_tiehi _7297__132 (.L_HI(net132));
 sg13g2_tiehi _7296__133 (.L_HI(net133));
 sg13g2_tiehi _7295__134 (.L_HI(net134));
 sg13g2_tiehi _7294__135 (.L_HI(net135));
 sg13g2_tiehi _7293__136 (.L_HI(net136));
 sg13g2_tiehi _7292__137 (.L_HI(net137));
 sg13g2_tiehi _7291__138 (.L_HI(net138));
 sg13g2_tiehi _7076__139 (.L_HI(net139));
 sg13g2_tiehi _7290__140 (.L_HI(net140));
 sg13g2_tiehi _7075__141 (.L_HI(net141));
 sg13g2_tiehi _7289__142 (.L_HI(net142));
 sg13g2_tiehi _7074__143 (.L_HI(net143));
 sg13g2_tiehi _7288__144 (.L_HI(net144));
 sg13g2_tiehi _7073__145 (.L_HI(net145));
 sg13g2_tiehi _7287__146 (.L_HI(net146));
 sg13g2_tiehi _7072__147 (.L_HI(net147));
 sg13g2_tiehi _7286__148 (.L_HI(net148));
 sg13g2_tiehi _7071__149 (.L_HI(net149));
 sg13g2_tiehi _7285__150 (.L_HI(net150));
 sg13g2_tiehi _7070__151 (.L_HI(net151));
 sg13g2_tiehi _7284__152 (.L_HI(net152));
 sg13g2_tiehi _7069__153 (.L_HI(net153));
 sg13g2_tiehi _7283__154 (.L_HI(net154));
 sg13g2_tiehi _7068__155 (.L_HI(net155));
 sg13g2_tiehi _7282__156 (.L_HI(net156));
 sg13g2_tiehi _7067__157 (.L_HI(net157));
 sg13g2_tiehi _7281__158 (.L_HI(net158));
 sg13g2_tiehi _7066__159 (.L_HI(net159));
 sg13g2_tiehi _7280__160 (.L_HI(net160));
 sg13g2_tiehi _7065__161 (.L_HI(net161));
 sg13g2_tiehi _7279__162 (.L_HI(net162));
 sg13g2_tiehi _7356__163 (.L_HI(net163));
 sg13g2_tiehi tt_um_a1k0n_demo_164 (.L_HI(net164));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_a1k0n_demo_2 (.L_LO(net2));
 sg13g2_tielo tt_um_a1k0n_demo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_a1k0n_demo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_a1k0n_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_a1k0n_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_a1k0n_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_a1k0n_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_a1k0n_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_a1k0n_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_a1k0n_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_a1k0n_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_a1k0n_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_a1k0n_demo_14 (.L_LO(net14));
 sg13g2_tiehi _7248__15 (.L_HI(net15));
 sg13g2_buf_2 _7521_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_1 _7522_ (.A(\vgademo.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7523_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_1786_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_1729_));
 sg13g2_buf_2 fanout814 (.A(net816),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_1660_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_1484_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(net821),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_1488_),
    .X(net821));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(net823));
 sg13g2_buf_2 fanout823 (.A(_2346_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_1487_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_1463_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(net827),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_1380_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_1512_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(net830),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_1461_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_1460_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_1533_),
    .X(net833));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(_1532_));
 sg13g2_buf_2 fanout835 (.A(_1532_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_1453_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_1453_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_0687_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net841),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_2484_),
    .X(net841));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(_1868_));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(_0668_));
 sg13g2_buf_2 fanout844 (.A(net846),
    .X(net844));
 sg13g2_buf_1 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_0626_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_1 fanout848 (.A(_1355_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net851),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_4 fanout851 (.X(net851),
    .A(_1355_));
 sg13g2_buf_2 fanout852 (.A(_1784_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_1353_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(net856),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_1350_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_0869_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_1329_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_0830_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_0829_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(net864),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_0829_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_0592_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_0592_),
    .X(net867));
 sg13g2_buf_1 fanout868 (.A(_0592_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_0575_),
    .X(net869));
 sg13g2_buf_1 fanout870 (.A(_0575_),
    .X(net870));
 sg13g2_buf_4 fanout871 (.X(net871),
    .A(net873));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_0574_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net881),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net881),
    .X(net876));
 sg13g2_buf_1 fanout877 (.A(net881),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(net880),
    .X(net878));
 sg13g2_buf_1 fanout879 (.A(net880),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_2726_),
    .X(net881));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(_2421_));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(_2420_));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(_1227_));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(net886));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(_0583_));
 sg13g2_buf_2 fanout887 (.A(_0583_),
    .X(net887));
 sg13g2_buf_4 fanout888 (.X(net888),
    .A(net889));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(net890));
 sg13g2_buf_2 fanout890 (.A(_2416_),
    .X(net890));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(_2416_));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(_0580_));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net897));
 sg13g2_buf_2 fanout894 (.A(net897),
    .X(net894));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(net897));
 sg13g2_buf_1 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_0580_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_0580_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net900),
    .X(net899));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(net902));
 sg13g2_buf_4 fanout901 (.X(net901),
    .A(net902));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(_0579_));
 sg13g2_buf_2 fanout903 (.A(_1396_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_1079_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_4 fanout906 (.X(net906),
    .A(_0653_));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_0652_),
    .X(net908));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(net915));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_1 fanout911 (.A(net913),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net914),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_0589_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(net919),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net918),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_0588_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(net924),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(net924),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_0582_),
    .X(net924));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(_0581_));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(_0651_));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(net929));
 sg13g2_buf_1 fanout928 (.A(net929),
    .X(net928));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(_0650_));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_4 fanout931 (.X(net931),
    .A(_3216_));
 sg13g2_buf_2 fanout932 (.A(_0701_),
    .X(net932));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(_0632_));
 sg13g2_buf_2 fanout934 (.A(_0624_),
    .X(net934));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(_2236_));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_2177_));
 sg13g2_buf_2 fanout937 (.A(net938),
    .X(net937));
 sg13g2_buf_1 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_3151_),
    .X(net939));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(_3132_));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(_3124_));
 sg13g2_buf_2 fanout942 (.A(_3111_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_3111_),
    .X(net943));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(_3110_));
 sg13g2_buf_4 fanout945 (.X(net945),
    .A(_3109_));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(net550));
 sg13g2_buf_2 fanout947 (.A(\vgademo.b_sin[11] ),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(net949),
    .X(net948));
 sg13g2_buf_1 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_4 fanout950 (.X(net950),
    .A(\vgademo.plane_dx_div.r[25] ));
 sg13g2_buf_2 fanout951 (.A(net952),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(\vgademo.b_cos[10] ),
    .X(net952));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(\vgademo.b_cos[9] ));
 sg13g2_buf_4 fanout954 (.X(net954),
    .A(\vgademo.b_cos[6] ));
 sg13g2_buf_2 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(\vgademo.v_count[9] ),
    .X(net956));
 sg13g2_buf_4 fanout957 (.X(net957),
    .A(\vgademo.v_count[7] ));
 sg13g2_buf_4 fanout958 (.X(net958),
    .A(net534));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(\vgademo.v_count[5] ));
 sg13g2_buf_2 fanout960 (.A(\vgademo.v_count[4] ),
    .X(net960));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(\vgademo.a_scrolly[11] ));
 sg13g2_buf_2 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_4 fanout963 (.X(net963),
    .A(\vgademo.a_scrolly[10] ));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(\vgademo.a_scrolly[9] ));
 sg13g2_buf_2 fanout965 (.A(\vgademo.a_scrolly[9] ),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_4 fanout967 (.X(net967),
    .A(net572));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(net969));
 sg13g2_buf_4 fanout969 (.X(net969),
    .A(net970));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(\vgademo.a_scrolly[7] ));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(net973));
 sg13g2_buf_2 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(\vgademo.a_scrolly[6] ),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net976),
    .X(net974));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(net976));
 sg13g2_buf_2 fanout976 (.A(\vgademo.a_scrolly[5] ),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(net978),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(net979),
    .X(net978));
 sg13g2_buf_1 fanout979 (.A(\vgademo.a_scrolly[4] ),
    .X(net979));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(net981));
 sg13g2_buf_4 fanout981 (.X(net981),
    .A(\vgademo.a_scrolly[3] ));
 sg13g2_buf_2 fanout982 (.A(net272),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(\vgademo.h_count[8] ),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(\vgademo.h_count[6] ),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(\vgademo.h_count[3] ),
    .X(net985));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(\vgademo.h_count[1] ));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(net988));
 sg13g2_buf_4 fanout988 (.X(net988),
    .A(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_buf_2 fanout989 (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(net989));
 sg13g2_buf_1 fanout990 (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(\vgademo.soundtrack.pulse_vol[0] ),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(net994),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(net995),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(\vgademo.audio_snare_frames[3] ),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net998),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_1 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(\vgademo.audio_snare_frames[2] ),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(\vgademo.audio_snare_frames[1] ),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(\vgademo.audio_snare_frames[1] ),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(net1004),
    .X(net1002));
 sg13g2_buf_1 fanout1003 (.A(net1004),
    .X(net1003));
 sg13g2_buf_1 fanout1004 (.A(net1006),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sg13g2_buf_1 fanout1006 (.A(\vgademo.audio_snare_frames[0] ),
    .X(net1006));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(net481));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(net1009));
 sg13g2_buf_4 fanout1009 (.X(net1009),
    .A(net267));
 sg13g2_buf_2 fanout1010 (.A(net567),
    .X(net1010));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(net247));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(net323));
 sg13g2_buf_4 fanout1013 (.X(net1013),
    .A(net1014));
 sg13g2_buf_2 fanout1014 (.A(net246),
    .X(net1014));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(net499));
 sg13g2_buf_2 fanout1016 (.A(net1017),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(\vgademo.audio_songpos[7] ),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(\vgademo.audio_songpos[6] ));
 sg13g2_buf_2 fanout1020 (.A(net1022),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(\vgademo.audio_songpos[5] ),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(net1026),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(net1026),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(\vgademo.audio_songpos[4] ),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(net1029),
    .X(net1027));
 sg13g2_buf_4 fanout1028 (.X(net1028),
    .A(net1029));
 sg13g2_buf_4 fanout1029 (.X(net1029),
    .A(\vgademo.audio_songpos[3] ));
 sg13g2_buf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(net1033),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(\vgademo.audio_songpos[2] ),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net1035),
    .X(net1034));
 sg13g2_buf_4 fanout1035 (.X(net1035),
    .A(\vgademo.audio_songpos[1] ));
 sg13g2_buf_2 fanout1036 (.A(net1037),
    .X(net1036));
 sg13g2_buf_1 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_4 fanout1038 (.X(net1038),
    .A(\vgademo.audio_songpos[0] ));
 sg13g2_buf_4 fanout1039 (.X(net1039),
    .A(\vgademo.linelfsr[1] ));
 sg13g2_buf_1 fanout1040 (.A(\vgademo.linelfsr[1] ),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(net441),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(\vgademo.linelfsr[0] ),
    .X(net1042));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(net1053));
 sg13g2_buf_2 fanout1044 (.A(net1053),
    .X(net1044));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(net1048));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1047));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1048));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(net1053));
 sg13g2_buf_4 fanout1049 (.X(net1049),
    .A(net1053));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(net1053));
 sg13g2_buf_4 fanout1051 (.X(net1051),
    .A(net1052));
 sg13g2_buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(rst_n));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(net1056));
 sg13g2_buf_2 fanout1055 (.A(net1056),
    .X(net1055));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(net1068));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(net1059));
 sg13g2_buf_4 fanout1058 (.X(net1058),
    .A(net1059));
 sg13g2_buf_4 fanout1059 (.X(net1059),
    .A(net1068));
 sg13g2_buf_4 fanout1060 (.X(net1060),
    .A(net1065));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(net1062));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(net1064));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(net1064));
 sg13g2_buf_2 fanout1064 (.A(net1065),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(net1068),
    .X(net1065));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(net1067));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(net1068));
 sg13g2_buf_2 fanout1068 (.A(rst_n),
    .X(net1068));
 sg13g2_tielo tt_um_a1k0n_demo_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_8 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_45_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_48_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_5_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_41_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_43_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_44_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_7_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_11_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_13_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_15_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_39_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_32_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_34_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_16_clk));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload33 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_24_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_30_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vgademo.soundtrack.sample_div_[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold2 (.A(\vgademo.soundtrack.noise_lfsr[11] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0180_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0085_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0143_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0084_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0175_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0082_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0182_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold10 (.A(\vgademo.soundtrack.tick_div_[0] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0162_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0083_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0177_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0107_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0206_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0096_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0172_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0094_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0170_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0095_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0171_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0108_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0089_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0088_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0087_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold26 (.A(\vgademo.soundtrack.pulse_osc_p[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0190_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0109_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0208_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0101_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0181_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold32 (.A(\vgademo.soundtrack.noise_lfsr[10] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0179_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0110_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0209_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0091_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold37 (.A(\vgademo.plane_dx_div.q[7] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0661_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold39 (.A(\vgademo.plane_dx_div.q[3] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0657_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0090_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vgademo.soundtrack.tick_div[6] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0796_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0168_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0086_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0125_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold47 (.A(\vgademo.soundtrack.sample_div[8] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold48 (.A(\vgademo.soundtrack.sample_div_[8] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold49 (.A(\vgademo.soundtrack.tick_div[4] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0166_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0111_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0106_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0188_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vgademo.a_sin[0] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold55 (.A(\vgademo.plane_u[0] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold56 (.A(_3092_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0365_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold58 (.A(\vgademo.soundtrack.pulse_osc_p[10] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0199_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold60 (.A(\vgademo.soundtrack.sigma_delta_accum[0] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold61 (.A(\vgademo.soundtrack.noise_lfsr[13] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0183_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0105_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold64 (.A(\vgademo.soundtrack.sample_div[4] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold65 (.A(\vgademo.soundtrack.sample_div_[4] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold66 (.A(\vgademo.soundtrack.sample_div[7] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold67 (.A(\vgademo.soundtrack.sample_div_[7] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold68 (.A(\vgademo.soundtrack.noise_lfsr[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0174_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0039_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0010_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0097_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0173_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold74 (.A(\vgademo.a_scrolly[11] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0243_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold76 (.A(audio),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0161_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold78 (.A(\vgademo.soundtrack.tick_div[2] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0164_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold80 (.A(\vgademo.soundtrack.sample_div[3] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold81 (.A(\vgademo.soundtrack.sample_div_[3] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold82 (.A(\vgademo.plane_dx_div.q[4] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold83 (.A(\vgademo.plane_dx_div.q[6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0660_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0104_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold86 (.A(\vgademo.soundtrack.tick_div[3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0165_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold88 (.A(\vgademo.a_cos[0] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0258_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold90 (.A(\vgademo.soundtrack.sample_div[0] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold91 (.A(\vgademo.soundtrack.sample_div_[1] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold92 (.A(\vgademo.soundtrack.pulse_osc_p[9] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0953_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0198_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold95 (.A(\vgademo.soundtrack.tri_osc_p[0] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0210_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0103_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0185_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold99 (.A(\vgademo.soundtrack.pulse_osc_p[13] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0202_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold101 (.A(\vgademo.v_count[4] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0250_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vgademo.plane_dx_div.q[8] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold104 (.A(\vgademo.soundtrack.sample_div[9] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold105 (.A(\vgademo.soundtrack.sample_div_[9] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold106 (.A(\vgademo.soundtrack.sample_div[5] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold107 (.A(\vgademo.soundtrack.pulse_osc_p[8] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0061_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold109 (.A(_3237_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0001_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold111 (.A(\vgademo.soundtrack.pulse_osc_p[11] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold112 (.A(\vgademo.soundtrack.tick_div[5] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold113 (.A(\vgademo.plane_dx_div.r[20] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0093_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0092_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold116 (.A(\vgademo.audio_kick_frames[2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold117 (.A(\vgademo.soundtrack.tri_osc_p[10] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0220_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold119 (.A(\vgademo.plane_u[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0331_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold121 (.A(\vgademo.b_cos[0] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold122 (.A(_2422_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0295_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold124 (.A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0195_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold126 (.A(\vgademo.soundtrack.tick_div[7] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold127 (.A(\vgademo.soundtrack.noise_lfsr[7] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0176_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold129 (.A(\vgademo.plane_dx_div.d[23] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold130 (.A(\vgademo.a_sin[1] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold131 (.A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold132 (.A(\vgademo.plane_u[11] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0341_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold134 (.A(\vgademo.b_sin[5] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0324_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold136 (.A(\vgademo.a_sin[2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0275_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold138 (.A(\vgademo.plane_dx_div.d[18] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold139 (.A(\vgademo.plane_dx_div.d[20] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold140 (.A(\vgademo.a_cos[1] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold141 (.A(\vgademo.v_count[5] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0251_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold143 (.A(\vgademo.soundtrack.noise_lfsr[0] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0184_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold145 (.A(\vgademo.soundtrack.pulse_osc_p[2] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold146 (.A(\vgademo.plane_du[1] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0355_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold148 (.A(\vgademo.plane_dx_div.d[22] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold149 (.A(\vgademo.plane_dx_div.r[21] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold150 (.A(\vgademo.plane_dx_div.d[24] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold151 (.A(\vgademo.scanline_audio_sample[0] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold152 (.A(\vgademo.plane_du[0] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0354_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold154 (.A(\vgademo.plane_u[4] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold155 (.A(\vgademo.a_cos[2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold156 (.A(\vgademo.linelfsr[10] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0122_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold158 (.A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold159 (.A(\vgademo.plane_dx_div.q[5] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0659_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold161 (.A(\vgademo.plane_dx_div.r[24] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold162 (.A(\vgademo.audio_beat_out[0] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold163 (.A(\vgademo.plane_u[8] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold164 (.A(\vgademo.plane_u[20] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold165 (.A(\vgademo.soundtrack.noise_lfsr[8] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0178_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold167 (.A(\vgademo.linelfsr[11] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0123_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold169 (.A(\vgademo.plane_dx_div.r[18] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0309_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold171 (.A(\vgademo.b_cos[1] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0296_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold173 (.A(\vgademo.plane_u[5] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold174 (.A(\vgademo.linelfsr[12] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold175 (.A(\vgademo.plane_dx_div.r[23] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold176 (.A(\vgademo.plane_dx_div.r[19] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0310_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold178 (.A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0193_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold180 (.A(\vgademo.b_cos[3] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0298_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold182 (.A(\vgademo.soundtrack.tri_osc_p[13] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0223_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold184 (.A(\vgademo.scanline_audio_sample[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold185 (.A(\vgademo.plane_dx_div.r[16] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0307_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold187 (.A(\vgademo.plane_dx_div.r[22] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold188 (.A(\vgademo.scanline_audio_sample[5] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold189 (.A(\vgademo.plane_u[6] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold190 (.A(\vgademo.scanline_audio_sample[2] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold191 (.A(\vgademo.plane_dx_div.d[21] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold192 (.A(\vgademo.a_cos[12] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold193 (.A(\vgademo.plane_dx_div.d[19] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold194 (.A(\vgademo.b_sin[7] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0326_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold196 (.A(\vgademo.plane_u[12] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0342_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold198 (.A(\vgademo.soundtrack.pulse_osc_p[7] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0196_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold200 (.A(\vgademo.plane_u[7] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold201 (.A(\vgademo.a_sin[5] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold202 (.A(\vgademo.a_sin[4] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0277_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold204 (.A(\vgademo.soundtrack.tri_osc_p[14] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0224_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold206 (.A(\vgademo.linelfsr[9] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold207 (.A(\vgademo.soundtrack.sigma_delta_accum[1] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold208 (.A(\vgademo.a_cos[3] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold209 (.A(\vgademo.plane_u[10] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold210 (.A(\vgademo.soundtrack.tri_osc_p[4] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold211 (.A(\vgademo.linelfsr[7] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0119_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold213 (.A(\vgademo.plane_u[3] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold214 (.A(\vgademo.b_sin[1] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0320_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold216 (.A(\vgademo.b_sin[2] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold217 (.A(\vgademo.plane_u[13] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0343_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold219 (.A(\vgademo.plane_u[2] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold220 (.A(\vgademo.linelfsr[8] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold221 (.A(\vgademo.a_sin[3] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0041_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0219_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold224 (.A(\vgademo.linelfsr[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0114_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold226 (.A(\vgademo.plane_u[14] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold227 (.A(\vgademo.plane_dx_div.d[17] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold228 (.A(\vgademo.linelfsr[5] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0117_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold230 (.A(\vgademo.soundtrack.tri_osc_p[1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold231 (.A(\vgademo.plane_dx_div.r[17] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold232 (.A(\vgademo.plane_dx_div.i[3] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0667_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold234 (.A(\vgademo.linelfsr[4] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold235 (.A(\vgademo.plane_u[21] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0351_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold237 (.A(\vgademo.plane_dx_div.i[0] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0664_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold239 (.A(\vgademo.a_scrolly[13] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0245_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold241 (.A(\vgademo.b_sin[3] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold242 (.A(_2669_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold243 (.A(\vgademo.soundtrack.tri_osc_p[12] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold244 (.A(_1045_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold245 (.A(\vgademo.soundtrack.tri_osc_p[3] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold246 (.A(\vgademo.a_cos[13] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0305_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0021_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold249 (.A(_1283_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold250 (.A(\vgademo.b_sin[0] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold251 (.A(\vgademo.soundtrack.pulse_osc_p[0] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold252 (.A(\vgademo.soundtrack.tri_osc_p[2] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold253 (.A(\vgademo.scanline_audio_sample[6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold254 (.A(\vgademo.b_sin[6] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold255 (.A(_2688_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold256 (.A(\vgademo.soundtrack.tri_osc_p[8] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0218_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0015_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold259 (.A(_1247_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0242_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold261 (.A(\vgademo.plane_u[16] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold262 (.A(_2972_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold263 (.A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold264 (.A(\vgademo.soundtrack.tri_osc_p[7] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0217_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold266 (.A(\vgademo.audio_kick_frames[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold267 (.A(\vgademo.b_cos[2] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold268 (.A(_2432_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0037_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold270 (.A(\vgademo.soundtrack.tri_osc_i[2] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold271 (.A(\vgademo.plane_u[9] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold272 (.A(\vgademo.b_sin[9] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0328_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold274 (.A(\vgademo.a_cos[11] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0303_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold276 (.A(\vgademo.soundtrack.tri_osc_p[11] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold277 (.A(\vgademo.linelfsr[0] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold278 (.A(\vgademo.linelfsr[6] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold279 (.A(\vgademo.b_cos[4] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0299_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold281 (.A(\vgademo.plane_u[19] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0349_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold283 (.A(\vgademo.soundtrack.tri_osc_p[5] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold284 (.A(\vgademo.a_sin[7] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold285 (.A(_2675_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold286 (.A(\vgademo.audio_beat_out[3] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0677_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0150_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold289 (.A(\vgademo.soundtrack.sample_div[2] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0567_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold291 (.A(\vgademo.soundtrack.sample_div_[2] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold292 (.A(\vgademo.soundtrack.sample_div[6] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold293 (.A(\vgademo.plane_du[3] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold294 (.A(\vgademo.plane_dx_div.d[16] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0034_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold296 (.A(_3221_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0004_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold298 (.A(\vgademo.v_count[2] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0248_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold300 (.A(\vgademo.a_cos[14] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold301 (.A(\vgademo.plane_u[17] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold302 (.A(\vgademo.a_sin[9] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold303 (.A(\vgademo.a_sin[13] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold304 (.A(_2719_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0033_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold306 (.A(\vgademo.soundtrack.tri_osc_p[6] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0216_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold308 (.A(\vgademo.b_cos[11] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold309 (.A(\vgademo.plane_du[2] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0356_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0035_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0014_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1277_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0253_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold315 (.A(\vgademo.a_sin[6] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0279_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold317 (.A(\vgademo.plane_dx_div.q[9] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0364_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold319 (.A(\vgademo.a_cos[10] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0302_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold321 (.A(\vgademo.scanline_audio_sample[4] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold322 (.A(\vgademo.a_sin[12] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold323 (.A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold324 (.A(\vgademo.a_sin[11] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold325 (.A(\vgademo.b_sin[8] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold326 (.A(\vgademo.a_sin[12] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold327 (.A(\vgademo.audio_beat_out[4] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0680_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0151_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold330 (.A(\vgademo.a_cos[6] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold331 (.A(\vgademo.soundtrack.pulse_osc_p[12] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold332 (.A(\vgademo.soundtrack.tick_div[1] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0795_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0163_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0023_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0358_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold337 (.A(\vgademo.soundtrack.sigma_delta_accum[9] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold338 (.A(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0065_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0241_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold341 (.A(\vgademo.scanline_audio_sample[3] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold342 (.A(\vgademo.plane_u[18] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold343 (.A(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0062_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0676_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0149_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold347 (.A(\vgademo.soundtrack.sigma_delta_accum[8] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold348 (.A(\vgademo.soundtrack.sigma_delta_accum_[8] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold349 (.A(\vgademo.soundtrack.sigma_delta_accum[13] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold350 (.A(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold351 (.A(\vgademo.a_cos[7] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold352 (.A(\vgademo.soundtrack.sigma_delta_accum[7] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold353 (.A(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold354 (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold355 (.A(\vgademo.soundtrack.sigma_delta_accum[5] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold356 (.A(\vgademo.soundtrack.sigma_delta_accum_[5] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold357 (.A(\vgademo.soundtrack.tri_osc_i[8] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0160_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold359 (.A(\vgademo.a_sin[10] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold360 (.A(\vgademo.soundtrack.sigma_delta_accum[11] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold361 (.A(\vgademo.a_cos[9] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold362 (.A(\vgademo.soundtrack.sigma_delta_accum[12] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold363 (.A(\vgademo.a_cos[5] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold364 (.A(\vgademo.a_cos[4] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold365 (.A(\vgademo.a_sin[8] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold366 (.A(\vgademo.v_count[8] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0254_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold368 (.A(\vgademo.soundtrack.sigma_delta_accum[3] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold369 (.A(\vgademo.soundtrack.sigma_delta_accum_[3] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold370 (.A(\vgademo.v_count[6] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0252_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0067_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0244_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold374 (.A(\vgademo.plane_dx_div.i[2] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0665_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0145_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold377 (.A(\vgademo.h_count[4] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold378 (.A(\vgademo.v_count[3] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0249_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold380 (.A(\vgademo.plane_dx[1] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0655_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold382 (.A(\vgademo.b_cos[5] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold383 (.A(\vgademo.linelfsr[2] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0113_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold385 (.A(\vgademo.soundtrack.sigma_delta_accum[14] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold386 (.A(\vgademo.b_sin[11] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0330_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0036_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0007_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold390 (.A(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold391 (.A(\vgademo.h_count[0] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0000_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold393 (.A(\vgademo.plane_dx[0] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold394 (.A(\vgademo.soundtrack.tri_osc_i[3] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold395 (.A(\vgademo.a_cos[8] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0038_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold397 (.A(_3232_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold398 (.A(\vgademo.plane_du[5] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold399 (.A(\vgademo.soundtrack.sigma_delta_accum[6] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold400 (.A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold401 (.A(\vgademo.soundtrack.sigma_delta_accum[4] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold402 (.A(\vgademo.soundtrack.sigma_delta_accum[2] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0026_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0362_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold405 (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold406 (.A(\vgademo.plane_dx[3] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0656_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold408 (.A(\vgademo.a_scrolly[8] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0240_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold410 (.A(\vgademo.plane_du[6] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold411 (.A(\vgademo.audio_beat_out[1] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0148_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold413 (.A(\vgademo.audio_kick_frames[0] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0203_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold415 (.A(\vgademo.plane_du[7] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold416 (.A(\vgademo.plane_u[15] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0075_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold418 (.A(\vgademo.bayer_j[0] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold419 (.A(_1258_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0078_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold421 (.A(\vgademo.h_count[9] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold422 (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold423 (.A(\vgademo.soundtrack.tri_osc_p[11] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0036_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold425 (.A(\vgademo.a_sin[13] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold426 (.A(\vgademo.audio_beat_out[4] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold427 (.A(\vgademo.plane_dx[3] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold428 (.A(\vgademo.soundtrack.tri_osc_i[2] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold429 (.A(_1003_),
    .X(net593));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_decap_8 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_12_436 ();
 sg13g2_decap_8 FILLER_12_443 ();
 sg13g2_decap_8 FILLER_12_450 ();
 sg13g2_decap_8 FILLER_12_457 ();
 sg13g2_decap_8 FILLER_12_464 ();
 sg13g2_decap_8 FILLER_12_471 ();
 sg13g2_decap_8 FILLER_12_478 ();
 sg13g2_decap_8 FILLER_12_485 ();
 sg13g2_decap_8 FILLER_12_492 ();
 sg13g2_decap_8 FILLER_12_499 ();
 sg13g2_decap_8 FILLER_12_506 ();
 sg13g2_decap_8 FILLER_12_513 ();
 sg13g2_decap_8 FILLER_12_520 ();
 sg13g2_decap_8 FILLER_12_527 ();
 sg13g2_decap_8 FILLER_12_534 ();
 sg13g2_decap_8 FILLER_12_541 ();
 sg13g2_decap_8 FILLER_12_548 ();
 sg13g2_decap_8 FILLER_12_555 ();
 sg13g2_decap_8 FILLER_12_562 ();
 sg13g2_decap_8 FILLER_12_569 ();
 sg13g2_decap_8 FILLER_12_576 ();
 sg13g2_decap_8 FILLER_12_583 ();
 sg13g2_decap_8 FILLER_12_590 ();
 sg13g2_decap_8 FILLER_12_597 ();
 sg13g2_decap_8 FILLER_12_604 ();
 sg13g2_decap_8 FILLER_12_611 ();
 sg13g2_decap_8 FILLER_12_618 ();
 sg13g2_decap_8 FILLER_12_625 ();
 sg13g2_decap_8 FILLER_12_632 ();
 sg13g2_decap_8 FILLER_12_639 ();
 sg13g2_decap_8 FILLER_12_646 ();
 sg13g2_decap_8 FILLER_12_653 ();
 sg13g2_decap_8 FILLER_12_660 ();
 sg13g2_decap_8 FILLER_12_667 ();
 sg13g2_decap_8 FILLER_12_674 ();
 sg13g2_decap_8 FILLER_12_681 ();
 sg13g2_decap_8 FILLER_12_688 ();
 sg13g2_decap_8 FILLER_12_695 ();
 sg13g2_decap_8 FILLER_12_702 ();
 sg13g2_decap_8 FILLER_12_709 ();
 sg13g2_decap_8 FILLER_12_716 ();
 sg13g2_decap_8 FILLER_12_723 ();
 sg13g2_decap_8 FILLER_12_730 ();
 sg13g2_decap_8 FILLER_12_737 ();
 sg13g2_decap_8 FILLER_12_744 ();
 sg13g2_decap_8 FILLER_12_751 ();
 sg13g2_decap_8 FILLER_12_758 ();
 sg13g2_decap_8 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_772 ();
 sg13g2_decap_8 FILLER_12_779 ();
 sg13g2_decap_8 FILLER_12_786 ();
 sg13g2_decap_8 FILLER_12_793 ();
 sg13g2_decap_8 FILLER_12_800 ();
 sg13g2_decap_8 FILLER_12_807 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_8 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_828 ();
 sg13g2_decap_8 FILLER_12_835 ();
 sg13g2_decap_8 FILLER_12_842 ();
 sg13g2_decap_8 FILLER_12_849 ();
 sg13g2_decap_4 FILLER_12_856 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_4 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_298 ();
 sg13g2_decap_4 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_328 ();
 sg13g2_fill_2 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_344 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_decap_8 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_13_415 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_decap_8 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_13_436 ();
 sg13g2_decap_8 FILLER_13_443 ();
 sg13g2_decap_8 FILLER_13_450 ();
 sg13g2_decap_8 FILLER_13_457 ();
 sg13g2_decap_8 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_471 ();
 sg13g2_decap_8 FILLER_13_478 ();
 sg13g2_decap_8 FILLER_13_485 ();
 sg13g2_decap_8 FILLER_13_492 ();
 sg13g2_decap_8 FILLER_13_499 ();
 sg13g2_decap_8 FILLER_13_506 ();
 sg13g2_decap_8 FILLER_13_513 ();
 sg13g2_decap_8 FILLER_13_520 ();
 sg13g2_decap_8 FILLER_13_527 ();
 sg13g2_decap_8 FILLER_13_534 ();
 sg13g2_decap_8 FILLER_13_541 ();
 sg13g2_decap_8 FILLER_13_548 ();
 sg13g2_decap_8 FILLER_13_555 ();
 sg13g2_decap_8 FILLER_13_562 ();
 sg13g2_decap_8 FILLER_13_569 ();
 sg13g2_decap_8 FILLER_13_576 ();
 sg13g2_decap_8 FILLER_13_583 ();
 sg13g2_decap_8 FILLER_13_590 ();
 sg13g2_decap_8 FILLER_13_597 ();
 sg13g2_decap_8 FILLER_13_604 ();
 sg13g2_decap_8 FILLER_13_611 ();
 sg13g2_decap_8 FILLER_13_618 ();
 sg13g2_decap_8 FILLER_13_625 ();
 sg13g2_decap_8 FILLER_13_632 ();
 sg13g2_decap_8 FILLER_13_639 ();
 sg13g2_decap_8 FILLER_13_646 ();
 sg13g2_decap_8 FILLER_13_653 ();
 sg13g2_decap_8 FILLER_13_660 ();
 sg13g2_decap_8 FILLER_13_667 ();
 sg13g2_decap_8 FILLER_13_674 ();
 sg13g2_decap_8 FILLER_13_681 ();
 sg13g2_decap_8 FILLER_13_688 ();
 sg13g2_decap_8 FILLER_13_695 ();
 sg13g2_decap_8 FILLER_13_702 ();
 sg13g2_decap_8 FILLER_13_709 ();
 sg13g2_decap_8 FILLER_13_716 ();
 sg13g2_decap_8 FILLER_13_723 ();
 sg13g2_decap_8 FILLER_13_730 ();
 sg13g2_decap_8 FILLER_13_737 ();
 sg13g2_decap_8 FILLER_13_744 ();
 sg13g2_decap_8 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_772 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_decap_8 FILLER_13_793 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_13_835 ();
 sg13g2_decap_8 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_decap_4 FILLER_13_856 ();
 sg13g2_fill_2 FILLER_13_860 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_41 ();
 sg13g2_decap_8 FILLER_14_48 ();
 sg13g2_fill_1 FILLER_14_55 ();
 sg13g2_decap_8 FILLER_14_61 ();
 sg13g2_decap_8 FILLER_14_68 ();
 sg13g2_decap_8 FILLER_14_75 ();
 sg13g2_fill_1 FILLER_14_82 ();
 sg13g2_fill_2 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_94 ();
 sg13g2_decap_8 FILLER_14_101 ();
 sg13g2_decap_8 FILLER_14_108 ();
 sg13g2_decap_8 FILLER_14_115 ();
 sg13g2_fill_2 FILLER_14_122 ();
 sg13g2_fill_1 FILLER_14_124 ();
 sg13g2_decap_8 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_4 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_fill_2 FILLER_14_378 ();
 sg13g2_fill_1 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_8 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_8 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_14_433 ();
 sg13g2_decap_8 FILLER_14_440 ();
 sg13g2_decap_8 FILLER_14_447 ();
 sg13g2_decap_8 FILLER_14_454 ();
 sg13g2_decap_8 FILLER_14_461 ();
 sg13g2_decap_8 FILLER_14_468 ();
 sg13g2_decap_8 FILLER_14_475 ();
 sg13g2_decap_8 FILLER_14_482 ();
 sg13g2_decap_8 FILLER_14_489 ();
 sg13g2_decap_8 FILLER_14_496 ();
 sg13g2_decap_8 FILLER_14_503 ();
 sg13g2_decap_8 FILLER_14_510 ();
 sg13g2_decap_8 FILLER_14_517 ();
 sg13g2_decap_8 FILLER_14_524 ();
 sg13g2_decap_8 FILLER_14_531 ();
 sg13g2_decap_8 FILLER_14_538 ();
 sg13g2_decap_8 FILLER_14_545 ();
 sg13g2_decap_8 FILLER_14_552 ();
 sg13g2_decap_8 FILLER_14_559 ();
 sg13g2_decap_8 FILLER_14_566 ();
 sg13g2_decap_8 FILLER_14_573 ();
 sg13g2_decap_8 FILLER_14_580 ();
 sg13g2_decap_8 FILLER_14_587 ();
 sg13g2_decap_8 FILLER_14_594 ();
 sg13g2_decap_8 FILLER_14_601 ();
 sg13g2_decap_8 FILLER_14_608 ();
 sg13g2_decap_8 FILLER_14_615 ();
 sg13g2_decap_8 FILLER_14_622 ();
 sg13g2_decap_8 FILLER_14_629 ();
 sg13g2_decap_8 FILLER_14_636 ();
 sg13g2_decap_8 FILLER_14_643 ();
 sg13g2_decap_8 FILLER_14_650 ();
 sg13g2_decap_8 FILLER_14_657 ();
 sg13g2_decap_8 FILLER_14_664 ();
 sg13g2_decap_8 FILLER_14_671 ();
 sg13g2_decap_8 FILLER_14_678 ();
 sg13g2_decap_8 FILLER_14_685 ();
 sg13g2_decap_8 FILLER_14_692 ();
 sg13g2_decap_8 FILLER_14_699 ();
 sg13g2_decap_8 FILLER_14_706 ();
 sg13g2_decap_8 FILLER_14_713 ();
 sg13g2_decap_8 FILLER_14_720 ();
 sg13g2_decap_8 FILLER_14_727 ();
 sg13g2_decap_8 FILLER_14_734 ();
 sg13g2_decap_8 FILLER_14_741 ();
 sg13g2_decap_8 FILLER_14_748 ();
 sg13g2_decap_8 FILLER_14_755 ();
 sg13g2_decap_8 FILLER_14_762 ();
 sg13g2_decap_8 FILLER_14_769 ();
 sg13g2_decap_8 FILLER_14_776 ();
 sg13g2_decap_8 FILLER_14_783 ();
 sg13g2_decap_8 FILLER_14_790 ();
 sg13g2_decap_8 FILLER_14_797 ();
 sg13g2_decap_8 FILLER_14_804 ();
 sg13g2_decap_8 FILLER_14_811 ();
 sg13g2_decap_8 FILLER_14_818 ();
 sg13g2_decap_8 FILLER_14_825 ();
 sg13g2_decap_8 FILLER_14_832 ();
 sg13g2_decap_8 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_8 FILLER_14_853 ();
 sg13g2_fill_2 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_25 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_fill_2 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_fill_1 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_fill_2 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_4 FILLER_15_313 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_decap_4 FILLER_15_344 ();
 sg13g2_fill_2 FILLER_15_395 ();
 sg13g2_fill_1 FILLER_15_397 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_431 ();
 sg13g2_decap_4 FILLER_15_450 ();
 sg13g2_fill_1 FILLER_15_454 ();
 sg13g2_decap_8 FILLER_15_464 ();
 sg13g2_decap_8 FILLER_15_471 ();
 sg13g2_decap_8 FILLER_15_478 ();
 sg13g2_decap_8 FILLER_15_485 ();
 sg13g2_decap_8 FILLER_15_492 ();
 sg13g2_decap_8 FILLER_15_499 ();
 sg13g2_decap_8 FILLER_15_506 ();
 sg13g2_decap_8 FILLER_15_513 ();
 sg13g2_decap_8 FILLER_15_520 ();
 sg13g2_decap_8 FILLER_15_527 ();
 sg13g2_decap_8 FILLER_15_534 ();
 sg13g2_decap_8 FILLER_15_541 ();
 sg13g2_decap_8 FILLER_15_548 ();
 sg13g2_decap_8 FILLER_15_555 ();
 sg13g2_decap_8 FILLER_15_562 ();
 sg13g2_decap_8 FILLER_15_569 ();
 sg13g2_decap_8 FILLER_15_576 ();
 sg13g2_decap_8 FILLER_15_583 ();
 sg13g2_decap_8 FILLER_15_590 ();
 sg13g2_decap_8 FILLER_15_597 ();
 sg13g2_decap_8 FILLER_15_604 ();
 sg13g2_decap_8 FILLER_15_611 ();
 sg13g2_decap_8 FILLER_15_618 ();
 sg13g2_decap_8 FILLER_15_625 ();
 sg13g2_decap_8 FILLER_15_632 ();
 sg13g2_decap_8 FILLER_15_639 ();
 sg13g2_decap_8 FILLER_15_646 ();
 sg13g2_decap_8 FILLER_15_653 ();
 sg13g2_decap_8 FILLER_15_660 ();
 sg13g2_decap_8 FILLER_15_667 ();
 sg13g2_decap_8 FILLER_15_674 ();
 sg13g2_decap_8 FILLER_15_681 ();
 sg13g2_decap_8 FILLER_15_688 ();
 sg13g2_decap_8 FILLER_15_695 ();
 sg13g2_decap_8 FILLER_15_702 ();
 sg13g2_decap_8 FILLER_15_709 ();
 sg13g2_decap_8 FILLER_15_716 ();
 sg13g2_decap_8 FILLER_15_723 ();
 sg13g2_decap_8 FILLER_15_730 ();
 sg13g2_decap_8 FILLER_15_737 ();
 sg13g2_decap_8 FILLER_15_744 ();
 sg13g2_decap_8 FILLER_15_751 ();
 sg13g2_decap_8 FILLER_15_758 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_8 FILLER_15_772 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_8 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_793 ();
 sg13g2_decap_8 FILLER_15_800 ();
 sg13g2_decap_8 FILLER_15_807 ();
 sg13g2_decap_8 FILLER_15_814 ();
 sg13g2_decap_8 FILLER_15_821 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_decap_8 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_849 ();
 sg13g2_decap_4 FILLER_15_856 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_30 ();
 sg13g2_decap_8 FILLER_16_37 ();
 sg13g2_decap_4 FILLER_16_93 ();
 sg13g2_fill_2 FILLER_16_97 ();
 sg13g2_decap_4 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_107 ();
 sg13g2_decap_4 FILLER_16_117 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_decap_4 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_190 ();
 sg13g2_fill_2 FILLER_16_248 ();
 sg13g2_fill_1 FILLER_16_250 ();
 sg13g2_decap_4 FILLER_16_282 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_decap_4 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_356 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_decap_4 FILLER_16_377 ();
 sg13g2_fill_1 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_4 FILLER_16_398 ();
 sg13g2_decap_8 FILLER_16_478 ();
 sg13g2_decap_8 FILLER_16_485 ();
 sg13g2_decap_8 FILLER_16_492 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_506 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_decap_8 FILLER_16_520 ();
 sg13g2_decap_8 FILLER_16_527 ();
 sg13g2_decap_8 FILLER_16_534 ();
 sg13g2_decap_8 FILLER_16_541 ();
 sg13g2_decap_8 FILLER_16_548 ();
 sg13g2_decap_8 FILLER_16_555 ();
 sg13g2_decap_8 FILLER_16_562 ();
 sg13g2_decap_8 FILLER_16_569 ();
 sg13g2_decap_8 FILLER_16_576 ();
 sg13g2_decap_8 FILLER_16_583 ();
 sg13g2_decap_8 FILLER_16_590 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_decap_8 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_611 ();
 sg13g2_decap_8 FILLER_16_618 ();
 sg13g2_decap_8 FILLER_16_625 ();
 sg13g2_decap_8 FILLER_16_632 ();
 sg13g2_decap_8 FILLER_16_639 ();
 sg13g2_decap_8 FILLER_16_646 ();
 sg13g2_decap_8 FILLER_16_653 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_8 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_674 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_decap_8 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_709 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_68 ();
 sg13g2_fill_1 FILLER_17_80 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_208 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_fill_2 FILLER_17_220 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_284 ();
 sg13g2_fill_2 FILLER_17_311 ();
 sg13g2_fill_1 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_4 FILLER_17_341 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_decap_4 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_fill_2 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_405 ();
 sg13g2_decap_4 FILLER_17_415 ();
 sg13g2_fill_2 FILLER_17_424 ();
 sg13g2_decap_4 FILLER_17_435 ();
 sg13g2_fill_1 FILLER_17_439 ();
 sg13g2_decap_8 FILLER_17_445 ();
 sg13g2_decap_8 FILLER_17_452 ();
 sg13g2_fill_1 FILLER_17_477 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_4 FILLER_18_37 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_4 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_decap_8 FILLER_18_139 ();
 sg13g2_decap_4 FILLER_18_146 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_4 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_decap_4 FILLER_18_253 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_1 FILLER_18_294 ();
 sg13g2_fill_2 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_313 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_fill_1 FILLER_18_377 ();
 sg13g2_decap_4 FILLER_18_391 ();
 sg13g2_fill_2 FILLER_18_395 ();
 sg13g2_decap_4 FILLER_18_418 ();
 sg13g2_fill_2 FILLER_18_443 ();
 sg13g2_fill_1 FILLER_18_445 ();
 sg13g2_decap_8 FILLER_18_454 ();
 sg13g2_decap_8 FILLER_18_461 ();
 sg13g2_decap_4 FILLER_18_468 ();
 sg13g2_fill_1 FILLER_18_480 ();
 sg13g2_decap_8 FILLER_18_499 ();
 sg13g2_decap_8 FILLER_18_506 ();
 sg13g2_decap_8 FILLER_18_513 ();
 sg13g2_decap_8 FILLER_18_520 ();
 sg13g2_decap_8 FILLER_18_527 ();
 sg13g2_decap_8 FILLER_18_534 ();
 sg13g2_decap_8 FILLER_18_541 ();
 sg13g2_decap_8 FILLER_18_548 ();
 sg13g2_decap_8 FILLER_18_555 ();
 sg13g2_decap_8 FILLER_18_562 ();
 sg13g2_decap_8 FILLER_18_569 ();
 sg13g2_decap_8 FILLER_18_576 ();
 sg13g2_decap_8 FILLER_18_583 ();
 sg13g2_decap_8 FILLER_18_590 ();
 sg13g2_decap_8 FILLER_18_597 ();
 sg13g2_decap_8 FILLER_18_604 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_decap_8 FILLER_18_632 ();
 sg13g2_decap_8 FILLER_18_639 ();
 sg13g2_decap_8 FILLER_18_646 ();
 sg13g2_decap_8 FILLER_18_653 ();
 sg13g2_decap_8 FILLER_18_660 ();
 sg13g2_decap_8 FILLER_18_667 ();
 sg13g2_decap_8 FILLER_18_674 ();
 sg13g2_decap_8 FILLER_18_681 ();
 sg13g2_decap_8 FILLER_18_688 ();
 sg13g2_decap_8 FILLER_18_695 ();
 sg13g2_decap_8 FILLER_18_702 ();
 sg13g2_decap_8 FILLER_18_709 ();
 sg13g2_decap_8 FILLER_18_716 ();
 sg13g2_decap_8 FILLER_18_723 ();
 sg13g2_decap_8 FILLER_18_730 ();
 sg13g2_decap_8 FILLER_18_737 ();
 sg13g2_decap_8 FILLER_18_744 ();
 sg13g2_decap_8 FILLER_18_751 ();
 sg13g2_decap_8 FILLER_18_758 ();
 sg13g2_decap_8 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_18_849 ();
 sg13g2_decap_4 FILLER_18_856 ();
 sg13g2_fill_2 FILLER_18_860 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_11 ();
 sg13g2_fill_1 FILLER_19_47 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_102 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_fill_1 FILLER_19_157 ();
 sg13g2_decap_8 FILLER_19_173 ();
 sg13g2_decap_4 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_decap_4 FILLER_19_232 ();
 sg13g2_fill_1 FILLER_19_253 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_270 ();
 sg13g2_decap_4 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_316 ();
 sg13g2_decap_4 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_fill_2 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_fill_2 FILLER_19_412 ();
 sg13g2_fill_1 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_428 ();
 sg13g2_fill_1 FILLER_19_435 ();
 sg13g2_decap_8 FILLER_19_454 ();
 sg13g2_fill_2 FILLER_19_461 ();
 sg13g2_fill_1 FILLER_19_463 ();
 sg13g2_fill_1 FILLER_19_481 ();
 sg13g2_decap_8 FILLER_19_508 ();
 sg13g2_decap_8 FILLER_19_515 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_536 ();
 sg13g2_decap_8 FILLER_19_543 ();
 sg13g2_decap_8 FILLER_19_550 ();
 sg13g2_decap_8 FILLER_19_557 ();
 sg13g2_decap_8 FILLER_19_564 ();
 sg13g2_decap_8 FILLER_19_571 ();
 sg13g2_decap_8 FILLER_19_578 ();
 sg13g2_decap_8 FILLER_19_585 ();
 sg13g2_decap_8 FILLER_19_592 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_decap_8 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_620 ();
 sg13g2_decap_8 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_634 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_decap_8 FILLER_19_648 ();
 sg13g2_decap_8 FILLER_19_655 ();
 sg13g2_decap_8 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_676 ();
 sg13g2_decap_8 FILLER_19_683 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_decap_8 FILLER_19_697 ();
 sg13g2_decap_8 FILLER_19_704 ();
 sg13g2_decap_8 FILLER_19_711 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_decap_8 FILLER_19_732 ();
 sg13g2_decap_8 FILLER_19_739 ();
 sg13g2_decap_8 FILLER_19_746 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_767 ();
 sg13g2_decap_8 FILLER_19_774 ();
 sg13g2_decap_8 FILLER_19_781 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_decap_8 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_8 FILLER_19_823 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_decap_8 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_844 ();
 sg13g2_decap_8 FILLER_19_851 ();
 sg13g2_decap_4 FILLER_19_858 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_59 ();
 sg13g2_decap_4 FILLER_20_66 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_83 ();
 sg13g2_decap_8 FILLER_20_90 ();
 sg13g2_decap_4 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_decap_4 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_256 ();
 sg13g2_decap_4 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_decap_4 FILLER_20_379 ();
 sg13g2_fill_1 FILLER_20_383 ();
 sg13g2_decap_4 FILLER_20_389 ();
 sg13g2_fill_1 FILLER_20_393 ();
 sg13g2_fill_1 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_decap_4 FILLER_20_428 ();
 sg13g2_fill_2 FILLER_20_432 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_4 FILLER_20_462 ();
 sg13g2_fill_2 FILLER_20_466 ();
 sg13g2_fill_2 FILLER_20_481 ();
 sg13g2_decap_8 FILLER_20_509 ();
 sg13g2_decap_8 FILLER_20_516 ();
 sg13g2_decap_8 FILLER_20_523 ();
 sg13g2_decap_8 FILLER_20_530 ();
 sg13g2_decap_8 FILLER_20_537 ();
 sg13g2_decap_8 FILLER_20_544 ();
 sg13g2_decap_8 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_558 ();
 sg13g2_decap_8 FILLER_20_565 ();
 sg13g2_decap_8 FILLER_20_572 ();
 sg13g2_decap_8 FILLER_20_579 ();
 sg13g2_decap_8 FILLER_20_586 ();
 sg13g2_decap_8 FILLER_20_593 ();
 sg13g2_decap_8 FILLER_20_600 ();
 sg13g2_decap_8 FILLER_20_607 ();
 sg13g2_decap_8 FILLER_20_614 ();
 sg13g2_decap_8 FILLER_20_621 ();
 sg13g2_decap_8 FILLER_20_628 ();
 sg13g2_decap_8 FILLER_20_635 ();
 sg13g2_decap_8 FILLER_20_642 ();
 sg13g2_decap_8 FILLER_20_649 ();
 sg13g2_decap_8 FILLER_20_656 ();
 sg13g2_decap_8 FILLER_20_663 ();
 sg13g2_decap_8 FILLER_20_670 ();
 sg13g2_decap_8 FILLER_20_677 ();
 sg13g2_decap_8 FILLER_20_684 ();
 sg13g2_decap_8 FILLER_20_691 ();
 sg13g2_decap_8 FILLER_20_698 ();
 sg13g2_decap_8 FILLER_20_705 ();
 sg13g2_decap_8 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_decap_8 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_decap_8 FILLER_20_740 ();
 sg13g2_decap_8 FILLER_20_747 ();
 sg13g2_decap_8 FILLER_20_754 ();
 sg13g2_decap_8 FILLER_20_761 ();
 sg13g2_decap_8 FILLER_20_768 ();
 sg13g2_decap_8 FILLER_20_775 ();
 sg13g2_decap_8 FILLER_20_782 ();
 sg13g2_decap_8 FILLER_20_789 ();
 sg13g2_decap_8 FILLER_20_796 ();
 sg13g2_decap_8 FILLER_20_803 ();
 sg13g2_decap_8 FILLER_20_810 ();
 sg13g2_decap_8 FILLER_20_817 ();
 sg13g2_decap_8 FILLER_20_824 ();
 sg13g2_decap_8 FILLER_20_831 ();
 sg13g2_decap_8 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_845 ();
 sg13g2_decap_8 FILLER_20_852 ();
 sg13g2_fill_2 FILLER_20_859 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_fill_2 FILLER_21_26 ();
 sg13g2_decap_4 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_96 ();
 sg13g2_decap_4 FILLER_21_137 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_160 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_191 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_4 FILLER_21_365 ();
 sg13g2_fill_1 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_373 ();
 sg13g2_decap_4 FILLER_21_395 ();
 sg13g2_fill_1 FILLER_21_411 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_fill_2 FILLER_21_424 ();
 sg13g2_fill_1 FILLER_21_426 ();
 sg13g2_fill_1 FILLER_21_446 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_fill_1 FILLER_21_475 ();
 sg13g2_fill_1 FILLER_21_485 ();
 sg13g2_decap_4 FILLER_21_518 ();
 sg13g2_decap_4 FILLER_21_526 ();
 sg13g2_fill_2 FILLER_21_530 ();
 sg13g2_decap_8 FILLER_21_537 ();
 sg13g2_decap_8 FILLER_21_544 ();
 sg13g2_decap_8 FILLER_21_551 ();
 sg13g2_decap_8 FILLER_21_558 ();
 sg13g2_decap_8 FILLER_21_565 ();
 sg13g2_decap_8 FILLER_21_572 ();
 sg13g2_decap_8 FILLER_21_579 ();
 sg13g2_decap_8 FILLER_21_586 ();
 sg13g2_decap_8 FILLER_21_593 ();
 sg13g2_decap_8 FILLER_21_600 ();
 sg13g2_decap_8 FILLER_21_607 ();
 sg13g2_decap_8 FILLER_21_614 ();
 sg13g2_decap_8 FILLER_21_621 ();
 sg13g2_decap_8 FILLER_21_628 ();
 sg13g2_decap_8 FILLER_21_635 ();
 sg13g2_decap_8 FILLER_21_642 ();
 sg13g2_decap_8 FILLER_21_649 ();
 sg13g2_decap_8 FILLER_21_656 ();
 sg13g2_decap_8 FILLER_21_663 ();
 sg13g2_decap_8 FILLER_21_670 ();
 sg13g2_decap_8 FILLER_21_677 ();
 sg13g2_decap_8 FILLER_21_684 ();
 sg13g2_decap_8 FILLER_21_691 ();
 sg13g2_decap_8 FILLER_21_698 ();
 sg13g2_decap_8 FILLER_21_705 ();
 sg13g2_decap_8 FILLER_21_712 ();
 sg13g2_decap_8 FILLER_21_719 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_decap_8 FILLER_21_740 ();
 sg13g2_decap_8 FILLER_21_747 ();
 sg13g2_decap_8 FILLER_21_754 ();
 sg13g2_decap_8 FILLER_21_761 ();
 sg13g2_decap_8 FILLER_21_768 ();
 sg13g2_decap_8 FILLER_21_775 ();
 sg13g2_decap_8 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_8 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_810 ();
 sg13g2_decap_8 FILLER_21_817 ();
 sg13g2_decap_8 FILLER_21_824 ();
 sg13g2_decap_8 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_838 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_11 ();
 sg13g2_decap_4 FILLER_22_17 ();
 sg13g2_fill_1 FILLER_22_48 ();
 sg13g2_decap_8 FILLER_22_58 ();
 sg13g2_decap_4 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_4 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_fill_1 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_381 ();
 sg13g2_decap_4 FILLER_22_386 ();
 sg13g2_fill_2 FILLER_22_390 ();
 sg13g2_decap_4 FILLER_22_400 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_4 FILLER_22_434 ();
 sg13g2_decap_4 FILLER_22_446 ();
 sg13g2_fill_2 FILLER_22_450 ();
 sg13g2_fill_2 FILLER_22_473 ();
 sg13g2_fill_1 FILLER_22_475 ();
 sg13g2_fill_2 FILLER_22_510 ();
 sg13g2_fill_1 FILLER_22_526 ();
 sg13g2_fill_1 FILLER_22_545 ();
 sg13g2_fill_2 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_571 ();
 sg13g2_decap_8 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_613 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_627 ();
 sg13g2_decap_8 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_decap_8 FILLER_22_648 ();
 sg13g2_decap_8 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_decap_8 FILLER_22_676 ();
 sg13g2_decap_8 FILLER_22_683 ();
 sg13g2_decap_8 FILLER_22_690 ();
 sg13g2_decap_8 FILLER_22_697 ();
 sg13g2_decap_8 FILLER_22_704 ();
 sg13g2_decap_8 FILLER_22_711 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_753 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_decap_8 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_788 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_decap_8 FILLER_22_809 ();
 sg13g2_decap_8 FILLER_22_816 ();
 sg13g2_decap_8 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_4 FILLER_22_858 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_36 ();
 sg13g2_decap_4 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_fill_1 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_decap_4 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_fill_2 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_234 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_fill_2 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_4 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_364 ();
 sg13g2_decap_4 FILLER_23_379 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_1 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_475 ();
 sg13g2_fill_1 FILLER_23_482 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_fill_1 FILLER_23_504 ();
 sg13g2_fill_1 FILLER_23_531 ();
 sg13g2_fill_2 FILLER_23_558 ();
 sg13g2_decap_8 FILLER_23_586 ();
 sg13g2_decap_8 FILLER_23_593 ();
 sg13g2_decap_8 FILLER_23_600 ();
 sg13g2_decap_8 FILLER_23_607 ();
 sg13g2_decap_8 FILLER_23_614 ();
 sg13g2_decap_8 FILLER_23_621 ();
 sg13g2_decap_8 FILLER_23_628 ();
 sg13g2_decap_8 FILLER_23_635 ();
 sg13g2_decap_8 FILLER_23_642 ();
 sg13g2_decap_8 FILLER_23_649 ();
 sg13g2_decap_8 FILLER_23_656 ();
 sg13g2_decap_8 FILLER_23_663 ();
 sg13g2_decap_8 FILLER_23_670 ();
 sg13g2_decap_8 FILLER_23_677 ();
 sg13g2_decap_8 FILLER_23_684 ();
 sg13g2_decap_8 FILLER_23_691 ();
 sg13g2_decap_8 FILLER_23_698 ();
 sg13g2_decap_8 FILLER_23_705 ();
 sg13g2_decap_8 FILLER_23_712 ();
 sg13g2_decap_8 FILLER_23_719 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_decap_8 FILLER_23_733 ();
 sg13g2_decap_8 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_747 ();
 sg13g2_decap_8 FILLER_23_754 ();
 sg13g2_decap_8 FILLER_23_761 ();
 sg13g2_decap_8 FILLER_23_768 ();
 sg13g2_decap_8 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_782 ();
 sg13g2_decap_8 FILLER_23_789 ();
 sg13g2_decap_8 FILLER_23_796 ();
 sg13g2_decap_8 FILLER_23_803 ();
 sg13g2_decap_8 FILLER_23_810 ();
 sg13g2_decap_8 FILLER_23_817 ();
 sg13g2_decap_8 FILLER_23_824 ();
 sg13g2_decap_8 FILLER_23_831 ();
 sg13g2_decap_8 FILLER_23_838 ();
 sg13g2_decap_8 FILLER_23_845 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_fill_2 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_58 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_90 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_110 ();
 sg13g2_decap_8 FILLER_24_117 ();
 sg13g2_decap_8 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_decap_4 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_fill_2 FILLER_24_157 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_206 ();
 sg13g2_decap_4 FILLER_24_213 ();
 sg13g2_decap_4 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_decap_4 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_357 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_4 FILLER_24_399 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_409 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_fill_2 FILLER_24_430 ();
 sg13g2_fill_1 FILLER_24_432 ();
 sg13g2_fill_2 FILLER_24_440 ();
 sg13g2_decap_8 FILLER_24_451 ();
 sg13g2_decap_8 FILLER_24_458 ();
 sg13g2_decap_8 FILLER_24_465 ();
 sg13g2_fill_1 FILLER_24_472 ();
 sg13g2_decap_4 FILLER_24_532 ();
 sg13g2_fill_2 FILLER_24_536 ();
 sg13g2_decap_4 FILLER_24_548 ();
 sg13g2_fill_1 FILLER_24_552 ();
 sg13g2_decap_8 FILLER_24_584 ();
 sg13g2_decap_8 FILLER_24_591 ();
 sg13g2_decap_8 FILLER_24_598 ();
 sg13g2_decap_8 FILLER_24_605 ();
 sg13g2_decap_4 FILLER_24_612 ();
 sg13g2_decap_8 FILLER_24_621 ();
 sg13g2_decap_8 FILLER_24_628 ();
 sg13g2_decap_8 FILLER_24_635 ();
 sg13g2_decap_8 FILLER_24_642 ();
 sg13g2_decap_8 FILLER_24_649 ();
 sg13g2_decap_8 FILLER_24_656 ();
 sg13g2_decap_8 FILLER_24_663 ();
 sg13g2_decap_8 FILLER_24_670 ();
 sg13g2_decap_8 FILLER_24_677 ();
 sg13g2_decap_8 FILLER_24_684 ();
 sg13g2_decap_8 FILLER_24_691 ();
 sg13g2_decap_8 FILLER_24_698 ();
 sg13g2_decap_8 FILLER_24_705 ();
 sg13g2_decap_8 FILLER_24_712 ();
 sg13g2_decap_8 FILLER_24_719 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_747 ();
 sg13g2_decap_8 FILLER_24_754 ();
 sg13g2_decap_8 FILLER_24_761 ();
 sg13g2_decap_8 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_775 ();
 sg13g2_decap_8 FILLER_24_782 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_decap_8 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_8 FILLER_24_831 ();
 sg13g2_decap_8 FILLER_24_838 ();
 sg13g2_decap_8 FILLER_24_845 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_fill_2 FILLER_24_859 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_75 ();
 sg13g2_fill_2 FILLER_25_96 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_fill_1 FILLER_25_127 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_decap_4 FILLER_25_209 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_decap_4 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_fill_1 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_25_418 ();
 sg13g2_decap_8 FILLER_25_443 ();
 sg13g2_fill_2 FILLER_25_450 ();
 sg13g2_fill_1 FILLER_25_452 ();
 sg13g2_decap_8 FILLER_25_457 ();
 sg13g2_fill_2 FILLER_25_464 ();
 sg13g2_fill_1 FILLER_25_466 ();
 sg13g2_decap_8 FILLER_25_491 ();
 sg13g2_decap_4 FILLER_25_498 ();
 sg13g2_fill_1 FILLER_25_502 ();
 sg13g2_fill_1 FILLER_25_521 ();
 sg13g2_fill_2 FILLER_25_548 ();
 sg13g2_fill_1 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_decap_8 FILLER_25_594 ();
 sg13g2_fill_1 FILLER_25_601 ();
 sg13g2_fill_2 FILLER_25_615 ();
 sg13g2_fill_1 FILLER_25_617 ();
 sg13g2_decap_8 FILLER_25_669 ();
 sg13g2_decap_8 FILLER_25_676 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_8 FILLER_25_690 ();
 sg13g2_decap_8 FILLER_25_697 ();
 sg13g2_decap_8 FILLER_25_704 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_8 FILLER_25_718 ();
 sg13g2_decap_8 FILLER_25_725 ();
 sg13g2_decap_8 FILLER_25_732 ();
 sg13g2_decap_8 FILLER_25_739 ();
 sg13g2_decap_8 FILLER_25_746 ();
 sg13g2_decap_8 FILLER_25_753 ();
 sg13g2_decap_8 FILLER_25_760 ();
 sg13g2_decap_8 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_774 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_8 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_8 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_4 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_2 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_fill_2 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_344 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_fill_1 FILLER_26_366 ();
 sg13g2_decap_4 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_fill_1 FILLER_26_417 ();
 sg13g2_fill_1 FILLER_26_437 ();
 sg13g2_decap_4 FILLER_26_443 ();
 sg13g2_fill_1 FILLER_26_447 ();
 sg13g2_decap_8 FILLER_26_468 ();
 sg13g2_fill_2 FILLER_26_475 ();
 sg13g2_decap_8 FILLER_26_486 ();
 sg13g2_fill_2 FILLER_26_493 ();
 sg13g2_fill_1 FILLER_26_495 ();
 sg13g2_fill_2 FILLER_26_542 ();
 sg13g2_fill_1 FILLER_26_544 ();
 sg13g2_fill_2 FILLER_26_559 ();
 sg13g2_fill_1 FILLER_26_570 ();
 sg13g2_fill_2 FILLER_26_618 ();
 sg13g2_fill_1 FILLER_26_620 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_fill_2 FILLER_26_637 ();
 sg13g2_decap_4 FILLER_26_660 ();
 sg13g2_decap_8 FILLER_26_685 ();
 sg13g2_decap_8 FILLER_26_692 ();
 sg13g2_decap_8 FILLER_26_699 ();
 sg13g2_decap_8 FILLER_26_706 ();
 sg13g2_decap_8 FILLER_26_713 ();
 sg13g2_decap_8 FILLER_26_720 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_decap_8 FILLER_26_734 ();
 sg13g2_decap_8 FILLER_26_741 ();
 sg13g2_decap_8 FILLER_26_748 ();
 sg13g2_decap_8 FILLER_26_755 ();
 sg13g2_decap_8 FILLER_26_762 ();
 sg13g2_decap_8 FILLER_26_769 ();
 sg13g2_decap_8 FILLER_26_776 ();
 sg13g2_decap_8 FILLER_26_783 ();
 sg13g2_decap_8 FILLER_26_790 ();
 sg13g2_decap_8 FILLER_26_797 ();
 sg13g2_decap_8 FILLER_26_804 ();
 sg13g2_decap_8 FILLER_26_811 ();
 sg13g2_decap_8 FILLER_26_818 ();
 sg13g2_decap_8 FILLER_26_825 ();
 sg13g2_decap_8 FILLER_26_832 ();
 sg13g2_decap_8 FILLER_26_839 ();
 sg13g2_decap_8 FILLER_26_846 ();
 sg13g2_decap_8 FILLER_26_853 ();
 sg13g2_fill_2 FILLER_26_860 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_16 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_decap_8 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_85 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_decap_4 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_decap_4 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_decap_4 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_230 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_258 ();
 sg13g2_decap_4 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_4 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_4 FILLER_27_386 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_411 ();
 sg13g2_fill_2 FILLER_27_418 ();
 sg13g2_fill_1 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_440 ();
 sg13g2_decap_4 FILLER_27_447 ();
 sg13g2_decap_8 FILLER_27_458 ();
 sg13g2_fill_1 FILLER_27_465 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_4 FILLER_27_497 ();
 sg13g2_fill_1 FILLER_27_501 ();
 sg13g2_fill_2 FILLER_27_554 ();
 sg13g2_decap_8 FILLER_27_705 ();
 sg13g2_decap_8 FILLER_27_712 ();
 sg13g2_decap_8 FILLER_27_719 ();
 sg13g2_decap_8 FILLER_27_726 ();
 sg13g2_decap_8 FILLER_27_733 ();
 sg13g2_decap_8 FILLER_27_740 ();
 sg13g2_decap_8 FILLER_27_747 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_decap_8 FILLER_27_761 ();
 sg13g2_decap_8 FILLER_27_768 ();
 sg13g2_decap_8 FILLER_27_775 ();
 sg13g2_decap_8 FILLER_27_782 ();
 sg13g2_decap_8 FILLER_27_789 ();
 sg13g2_decap_8 FILLER_27_796 ();
 sg13g2_decap_8 FILLER_27_803 ();
 sg13g2_decap_8 FILLER_27_810 ();
 sg13g2_decap_8 FILLER_27_817 ();
 sg13g2_decap_8 FILLER_27_824 ();
 sg13g2_decap_8 FILLER_27_831 ();
 sg13g2_decap_8 FILLER_27_838 ();
 sg13g2_decap_8 FILLER_27_845 ();
 sg13g2_decap_8 FILLER_27_852 ();
 sg13g2_fill_2 FILLER_27_859 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_decap_8 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_66 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_decap_4 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_4 FILLER_28_130 ();
 sg13g2_decap_4 FILLER_28_142 ();
 sg13g2_fill_2 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_4 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_fill_1 FILLER_28_296 ();
 sg13g2_decap_8 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_4 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_decap_4 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_4 FILLER_28_383 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_4 FILLER_28_414 ();
 sg13g2_fill_2 FILLER_28_426 ();
 sg13g2_fill_1 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_4 FILLER_28_441 ();
 sg13g2_fill_2 FILLER_28_445 ();
 sg13g2_decap_4 FILLER_28_466 ();
 sg13g2_fill_2 FILLER_28_470 ();
 sg13g2_fill_2 FILLER_28_486 ();
 sg13g2_fill_1 FILLER_28_514 ();
 sg13g2_fill_1 FILLER_28_565 ();
 sg13g2_fill_2 FILLER_28_576 ();
 sg13g2_fill_2 FILLER_28_613 ();
 sg13g2_fill_1 FILLER_28_615 ();
 sg13g2_fill_1 FILLER_28_630 ();
 sg13g2_decap_4 FILLER_28_640 ();
 sg13g2_fill_2 FILLER_28_644 ();
 sg13g2_fill_2 FILLER_28_660 ();
 sg13g2_fill_1 FILLER_28_662 ();
 sg13g2_decap_4 FILLER_28_666 ();
 sg13g2_fill_2 FILLER_28_670 ();
 sg13g2_decap_8 FILLER_28_698 ();
 sg13g2_decap_8 FILLER_28_705 ();
 sg13g2_decap_8 FILLER_28_712 ();
 sg13g2_decap_8 FILLER_28_719 ();
 sg13g2_decap_8 FILLER_28_726 ();
 sg13g2_decap_8 FILLER_28_733 ();
 sg13g2_decap_8 FILLER_28_740 ();
 sg13g2_decap_8 FILLER_28_747 ();
 sg13g2_decap_8 FILLER_28_754 ();
 sg13g2_decap_8 FILLER_28_761 ();
 sg13g2_decap_8 FILLER_28_768 ();
 sg13g2_decap_8 FILLER_28_775 ();
 sg13g2_decap_8 FILLER_28_782 ();
 sg13g2_decap_8 FILLER_28_789 ();
 sg13g2_decap_8 FILLER_28_796 ();
 sg13g2_decap_8 FILLER_28_803 ();
 sg13g2_decap_8 FILLER_28_810 ();
 sg13g2_decap_8 FILLER_28_817 ();
 sg13g2_decap_8 FILLER_28_824 ();
 sg13g2_decap_8 FILLER_28_831 ();
 sg13g2_decap_8 FILLER_28_838 ();
 sg13g2_decap_8 FILLER_28_845 ();
 sg13g2_decap_8 FILLER_28_852 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_18 ();
 sg13g2_decap_4 FILLER_29_24 ();
 sg13g2_decap_8 FILLER_29_55 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_4 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_decap_4 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_129 ();
 sg13g2_decap_4 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_decap_4 FILLER_29_184 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_decap_4 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_decap_4 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_415 ();
 sg13g2_fill_2 FILLER_29_422 ();
 sg13g2_fill_1 FILLER_29_424 ();
 sg13g2_fill_1 FILLER_29_443 ();
 sg13g2_fill_2 FILLER_29_449 ();
 sg13g2_fill_2 FILLER_29_460 ();
 sg13g2_fill_1 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_482 ();
 sg13g2_decap_4 FILLER_29_489 ();
 sg13g2_fill_1 FILLER_29_493 ();
 sg13g2_fill_2 FILLER_29_548 ();
 sg13g2_fill_2 FILLER_29_569 ();
 sg13g2_fill_2 FILLER_29_580 ();
 sg13g2_fill_1 FILLER_29_582 ();
 sg13g2_decap_4 FILLER_29_620 ();
 sg13g2_fill_1 FILLER_29_624 ();
 sg13g2_decap_4 FILLER_29_633 ();
 sg13g2_fill_2 FILLER_29_671 ();
 sg13g2_decap_8 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_711 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_decap_8 FILLER_29_746 ();
 sg13g2_decap_8 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_decap_8 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_4 FILLER_29_858 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_17 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_30 ();
 sg13g2_fill_2 FILLER_30_41 ();
 sg13g2_fill_1 FILLER_30_43 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_132 ();
 sg13g2_fill_2 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_197 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_4 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_fill_2 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_355 ();
 sg13g2_decap_8 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_4 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_30_409 ();
 sg13g2_decap_4 FILLER_30_416 ();
 sg13g2_fill_2 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_440 ();
 sg13g2_decap_8 FILLER_30_447 ();
 sg13g2_fill_2 FILLER_30_454 ();
 sg13g2_fill_1 FILLER_30_456 ();
 sg13g2_decap_4 FILLER_30_472 ();
 sg13g2_decap_8 FILLER_30_486 ();
 sg13g2_fill_1 FILLER_30_493 ();
 sg13g2_fill_2 FILLER_30_504 ();
 sg13g2_fill_2 FILLER_30_528 ();
 sg13g2_fill_1 FILLER_30_530 ();
 sg13g2_decap_4 FILLER_30_639 ();
 sg13g2_decap_4 FILLER_30_652 ();
 sg13g2_fill_1 FILLER_30_656 ();
 sg13g2_decap_4 FILLER_30_682 ();
 sg13g2_fill_2 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_697 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_725 ();
 sg13g2_decap_8 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_8 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_4 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_39 ();
 sg13g2_decap_4 FILLER_31_44 ();
 sg13g2_decap_8 FILLER_31_52 ();
 sg13g2_decap_8 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_decap_4 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_decap_4 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_120 ();
 sg13g2_decap_4 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_141 ();
 sg13g2_decap_4 FILLER_31_148 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_176 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_223 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_decap_4 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_31_387 ();
 sg13g2_fill_1 FILLER_31_389 ();
 sg13g2_fill_2 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_fill_2 FILLER_31_448 ();
 sg13g2_decap_4 FILLER_31_470 ();
 sg13g2_fill_2 FILLER_31_474 ();
 sg13g2_decap_8 FILLER_31_547 ();
 sg13g2_fill_2 FILLER_31_575 ();
 sg13g2_decap_4 FILLER_31_626 ();
 sg13g2_fill_2 FILLER_31_630 ();
 sg13g2_decap_4 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_685 ();
 sg13g2_decap_8 FILLER_31_692 ();
 sg13g2_decap_8 FILLER_31_699 ();
 sg13g2_decap_8 FILLER_31_706 ();
 sg13g2_decap_8 FILLER_31_713 ();
 sg13g2_decap_8 FILLER_31_720 ();
 sg13g2_decap_8 FILLER_31_727 ();
 sg13g2_decap_8 FILLER_31_734 ();
 sg13g2_decap_8 FILLER_31_741 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_decap_8 FILLER_31_769 ();
 sg13g2_decap_8 FILLER_31_776 ();
 sg13g2_decap_8 FILLER_31_783 ();
 sg13g2_decap_8 FILLER_31_790 ();
 sg13g2_decap_8 FILLER_31_797 ();
 sg13g2_decap_8 FILLER_31_804 ();
 sg13g2_decap_8 FILLER_31_811 ();
 sg13g2_decap_8 FILLER_31_818 ();
 sg13g2_decap_8 FILLER_31_825 ();
 sg13g2_decap_8 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_decap_8 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_853 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_19 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_decap_4 FILLER_32_60 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_fill_2 FILLER_32_75 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_decap_4 FILLER_32_120 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_decap_4 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_182 ();
 sg13g2_decap_4 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_247 ();
 sg13g2_decap_8 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_261 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_2 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_decap_4 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_decap_4 FILLER_32_402 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_decap_4 FILLER_32_418 ();
 sg13g2_decap_8 FILLER_32_444 ();
 sg13g2_decap_8 FILLER_32_451 ();
 sg13g2_fill_1 FILLER_32_458 ();
 sg13g2_fill_2 FILLER_32_468 ();
 sg13g2_decap_4 FILLER_32_486 ();
 sg13g2_fill_1 FILLER_32_490 ();
 sg13g2_decap_4 FILLER_32_514 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_decap_4 FILLER_32_529 ();
 sg13g2_fill_2 FILLER_32_533 ();
 sg13g2_fill_2 FILLER_32_545 ();
 sg13g2_fill_1 FILLER_32_547 ();
 sg13g2_fill_2 FILLER_32_583 ();
 sg13g2_decap_4 FILLER_32_616 ();
 sg13g2_fill_2 FILLER_32_655 ();
 sg13g2_fill_1 FILLER_32_657 ();
 sg13g2_fill_1 FILLER_32_667 ();
 sg13g2_decap_8 FILLER_32_694 ();
 sg13g2_decap_8 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_708 ();
 sg13g2_decap_8 FILLER_32_715 ();
 sg13g2_decap_8 FILLER_32_722 ();
 sg13g2_decap_8 FILLER_32_729 ();
 sg13g2_decap_8 FILLER_32_736 ();
 sg13g2_decap_8 FILLER_32_743 ();
 sg13g2_decap_8 FILLER_32_750 ();
 sg13g2_decap_8 FILLER_32_757 ();
 sg13g2_decap_8 FILLER_32_764 ();
 sg13g2_decap_8 FILLER_32_771 ();
 sg13g2_decap_8 FILLER_32_778 ();
 sg13g2_decap_8 FILLER_32_785 ();
 sg13g2_decap_8 FILLER_32_792 ();
 sg13g2_decap_8 FILLER_32_799 ();
 sg13g2_decap_8 FILLER_32_806 ();
 sg13g2_decap_8 FILLER_32_813 ();
 sg13g2_decap_8 FILLER_32_820 ();
 sg13g2_decap_8 FILLER_32_827 ();
 sg13g2_decap_8 FILLER_32_834 ();
 sg13g2_decap_8 FILLER_32_841 ();
 sg13g2_decap_8 FILLER_32_848 ();
 sg13g2_decap_8 FILLER_32_855 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_25 ();
 sg13g2_decap_4 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_43 ();
 sg13g2_fill_1 FILLER_33_50 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_64 ();
 sg13g2_decap_4 FILLER_33_71 ();
 sg13g2_fill_2 FILLER_33_75 ();
 sg13g2_decap_4 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_2 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_4 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_decap_4 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_decap_8 FILLER_33_325 ();
 sg13g2_decap_4 FILLER_33_339 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_379 ();
 sg13g2_fill_2 FILLER_33_399 ();
 sg13g2_fill_1 FILLER_33_401 ();
 sg13g2_fill_2 FILLER_33_433 ();
 sg13g2_fill_1 FILLER_33_461 ();
 sg13g2_fill_2 FILLER_33_514 ();
 sg13g2_decap_8 FILLER_33_554 ();
 sg13g2_fill_2 FILLER_33_561 ();
 sg13g2_fill_1 FILLER_33_563 ();
 sg13g2_decap_4 FILLER_33_601 ();
 sg13g2_fill_1 FILLER_33_605 ();
 sg13g2_fill_2 FILLER_33_632 ();
 sg13g2_fill_1 FILLER_33_634 ();
 sg13g2_fill_1 FILLER_33_643 ();
 sg13g2_fill_2 FILLER_33_653 ();
 sg13g2_fill_1 FILLER_33_655 ();
 sg13g2_decap_4 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_682 ();
 sg13g2_decap_8 FILLER_33_687 ();
 sg13g2_decap_8 FILLER_33_694 ();
 sg13g2_decap_8 FILLER_33_701 ();
 sg13g2_decap_8 FILLER_33_708 ();
 sg13g2_fill_2 FILLER_33_715 ();
 sg13g2_fill_1 FILLER_33_717 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_38 ();
 sg13g2_decap_8 FILLER_34_55 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_decap_4 FILLER_34_89 ();
 sg13g2_fill_2 FILLER_34_93 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_121 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_fill_1 FILLER_34_130 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_159 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_4 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_decap_4 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_4 FILLER_34_420 ();
 sg13g2_fill_1 FILLER_34_424 ();
 sg13g2_decap_4 FILLER_34_443 ();
 sg13g2_fill_1 FILLER_34_447 ();
 sg13g2_fill_1 FILLER_34_465 ();
 sg13g2_fill_2 FILLER_34_475 ();
 sg13g2_fill_1 FILLER_34_477 ();
 sg13g2_fill_2 FILLER_34_492 ();
 sg13g2_decap_8 FILLER_34_520 ();
 sg13g2_decap_4 FILLER_34_527 ();
 sg13g2_fill_2 FILLER_34_531 ();
 sg13g2_decap_4 FILLER_34_564 ();
 sg13g2_fill_2 FILLER_34_568 ();
 sg13g2_fill_2 FILLER_34_583 ();
 sg13g2_decap_4 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_decap_4 FILLER_34_611 ();
 sg13g2_fill_1 FILLER_34_615 ();
 sg13g2_fill_2 FILLER_34_626 ();
 sg13g2_fill_1 FILLER_34_628 ();
 sg13g2_decap_8 FILLER_34_638 ();
 sg13g2_fill_1 FILLER_34_645 ();
 sg13g2_decap_8 FILLER_34_734 ();
 sg13g2_decap_8 FILLER_34_741 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_decap_8 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_decap_8 FILLER_34_769 ();
 sg13g2_decap_8 FILLER_34_776 ();
 sg13g2_decap_8 FILLER_34_783 ();
 sg13g2_decap_8 FILLER_34_790 ();
 sg13g2_decap_8 FILLER_34_797 ();
 sg13g2_decap_8 FILLER_34_804 ();
 sg13g2_decap_8 FILLER_34_811 ();
 sg13g2_decap_8 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_61 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_117 ();
 sg13g2_decap_4 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_203 ();
 sg13g2_decap_4 FILLER_35_261 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_301 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_fill_2 FILLER_35_409 ();
 sg13g2_fill_2 FILLER_35_460 ();
 sg13g2_fill_1 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_fill_2 FILLER_35_545 ();
 sg13g2_fill_2 FILLER_35_591 ();
 sg13g2_fill_1 FILLER_35_593 ();
 sg13g2_fill_2 FILLER_35_620 ();
 sg13g2_decap_8 FILLER_35_656 ();
 sg13g2_decap_8 FILLER_35_663 ();
 sg13g2_fill_1 FILLER_35_688 ();
 sg13g2_fill_2 FILLER_35_707 ();
 sg13g2_fill_1 FILLER_35_709 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_44 ();
 sg13g2_decap_8 FILLER_36_51 ();
 sg13g2_decap_8 FILLER_36_58 ();
 sg13g2_fill_2 FILLER_36_65 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_4 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_155 ();
 sg13g2_decap_4 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_4 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_362 ();
 sg13g2_decap_4 FILLER_36_369 ();
 sg13g2_fill_2 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_decap_8 FILLER_36_430 ();
 sg13g2_fill_2 FILLER_36_437 ();
 sg13g2_fill_1 FILLER_36_439 ();
 sg13g2_fill_2 FILLER_36_449 ();
 sg13g2_fill_1 FILLER_36_451 ();
 sg13g2_decap_8 FILLER_36_457 ();
 sg13g2_decap_4 FILLER_36_464 ();
 sg13g2_fill_1 FILLER_36_468 ();
 sg13g2_decap_8 FILLER_36_495 ();
 sg13g2_fill_1 FILLER_36_502 ();
 sg13g2_fill_2 FILLER_36_516 ();
 sg13g2_fill_1 FILLER_36_527 ();
 sg13g2_fill_1 FILLER_36_536 ();
 sg13g2_fill_1 FILLER_36_564 ();
 sg13g2_decap_8 FILLER_36_569 ();
 sg13g2_fill_2 FILLER_36_576 ();
 sg13g2_decap_8 FILLER_36_604 ();
 sg13g2_decap_8 FILLER_36_611 ();
 sg13g2_decap_8 FILLER_36_618 ();
 sg13g2_decap_4 FILLER_36_625 ();
 sg13g2_fill_1 FILLER_36_629 ();
 sg13g2_fill_2 FILLER_36_637 ();
 sg13g2_fill_2 FILLER_36_656 ();
 sg13g2_fill_2 FILLER_36_684 ();
 sg13g2_fill_1 FILLER_36_686 ();
 sg13g2_fill_1 FILLER_36_691 ();
 sg13g2_decap_8 FILLER_36_701 ();
 sg13g2_decap_4 FILLER_36_708 ();
 sg13g2_fill_1 FILLER_36_712 ();
 sg13g2_decap_8 FILLER_36_743 ();
 sg13g2_decap_8 FILLER_36_750 ();
 sg13g2_decap_8 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_764 ();
 sg13g2_decap_8 FILLER_36_771 ();
 sg13g2_decap_8 FILLER_36_778 ();
 sg13g2_decap_8 FILLER_36_785 ();
 sg13g2_decap_8 FILLER_36_792 ();
 sg13g2_decap_8 FILLER_36_799 ();
 sg13g2_decap_8 FILLER_36_806 ();
 sg13g2_decap_8 FILLER_36_813 ();
 sg13g2_decap_8 FILLER_36_820 ();
 sg13g2_decap_8 FILLER_36_827 ();
 sg13g2_decap_8 FILLER_36_834 ();
 sg13g2_decap_8 FILLER_36_841 ();
 sg13g2_decap_8 FILLER_36_848 ();
 sg13g2_decap_8 FILLER_36_855 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_18 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_decap_4 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_decap_4 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_322 ();
 sg13g2_decap_4 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_4 FILLER_37_385 ();
 sg13g2_fill_2 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_411 ();
 sg13g2_decap_8 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_425 ();
 sg13g2_fill_2 FILLER_37_455 ();
 sg13g2_fill_1 FILLER_37_457 ();
 sg13g2_decap_4 FILLER_37_463 ();
 sg13g2_fill_2 FILLER_37_467 ();
 sg13g2_decap_4 FILLER_37_474 ();
 sg13g2_decap_4 FILLER_37_486 ();
 sg13g2_decap_8 FILLER_37_519 ();
 sg13g2_fill_2 FILLER_37_531 ();
 sg13g2_fill_1 FILLER_37_533 ();
 sg13g2_fill_2 FILLER_37_558 ();
 sg13g2_fill_1 FILLER_37_560 ();
 sg13g2_decap_4 FILLER_37_575 ();
 sg13g2_fill_2 FILLER_37_584 ();
 sg13g2_fill_1 FILLER_37_586 ();
 sg13g2_decap_8 FILLER_37_596 ();
 sg13g2_decap_4 FILLER_37_603 ();
 sg13g2_decap_8 FILLER_37_610 ();
 sg13g2_decap_4 FILLER_37_622 ();
 sg13g2_decap_8 FILLER_37_671 ();
 sg13g2_fill_2 FILLER_37_678 ();
 sg13g2_fill_2 FILLER_37_720 ();
 sg13g2_fill_1 FILLER_37_722 ();
 sg13g2_decap_8 FILLER_37_741 ();
 sg13g2_decap_8 FILLER_37_748 ();
 sg13g2_decap_8 FILLER_37_755 ();
 sg13g2_decap_8 FILLER_37_762 ();
 sg13g2_decap_8 FILLER_37_769 ();
 sg13g2_decap_8 FILLER_37_776 ();
 sg13g2_decap_8 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_decap_8 FILLER_37_797 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_4 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_39 ();
 sg13g2_decap_8 FILLER_38_54 ();
 sg13g2_fill_1 FILLER_38_61 ();
 sg13g2_decap_8 FILLER_38_89 ();
 sg13g2_fill_1 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_4 FILLER_38_299 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_fill_2 FILLER_38_356 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_decap_4 FILLER_38_442 ();
 sg13g2_fill_1 FILLER_38_446 ();
 sg13g2_decap_4 FILLER_38_456 ();
 sg13g2_fill_2 FILLER_38_486 ();
 sg13g2_decap_4 FILLER_38_496 ();
 sg13g2_fill_1 FILLER_38_515 ();
 sg13g2_decap_4 FILLER_38_526 ();
 sg13g2_fill_1 FILLER_38_538 ();
 sg13g2_decap_4 FILLER_38_547 ();
 sg13g2_fill_1 FILLER_38_551 ();
 sg13g2_decap_4 FILLER_38_570 ();
 sg13g2_fill_2 FILLER_38_589 ();
 sg13g2_fill_1 FILLER_38_617 ();
 sg13g2_fill_2 FILLER_38_644 ();
 sg13g2_fill_1 FILLER_38_646 ();
 sg13g2_decap_8 FILLER_38_671 ();
 sg13g2_decap_4 FILLER_38_694 ();
 sg13g2_fill_1 FILLER_38_698 ();
 sg13g2_fill_2 FILLER_38_703 ();
 sg13g2_fill_1 FILLER_38_705 ();
 sg13g2_fill_2 FILLER_38_710 ();
 sg13g2_decap_8 FILLER_38_738 ();
 sg13g2_decap_8 FILLER_38_745 ();
 sg13g2_decap_8 FILLER_38_752 ();
 sg13g2_decap_8 FILLER_38_759 ();
 sg13g2_decap_8 FILLER_38_766 ();
 sg13g2_decap_8 FILLER_38_773 ();
 sg13g2_decap_8 FILLER_38_780 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_decap_8 FILLER_38_794 ();
 sg13g2_decap_8 FILLER_38_801 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_829 ();
 sg13g2_decap_8 FILLER_38_836 ();
 sg13g2_decap_8 FILLER_38_843 ();
 sg13g2_decap_8 FILLER_38_850 ();
 sg13g2_decap_4 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_fill_2 FILLER_39_49 ();
 sg13g2_decap_4 FILLER_39_99 ();
 sg13g2_fill_2 FILLER_39_103 ();
 sg13g2_decap_8 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_130 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_decap_8 FILLER_39_142 ();
 sg13g2_decap_8 FILLER_39_153 ();
 sg13g2_fill_2 FILLER_39_160 ();
 sg13g2_fill_1 FILLER_39_162 ();
 sg13g2_fill_2 FILLER_39_180 ();
 sg13g2_decap_8 FILLER_39_186 ();
 sg13g2_decap_8 FILLER_39_193 ();
 sg13g2_decap_4 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_204 ();
 sg13g2_fill_2 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_222 ();
 sg13g2_decap_8 FILLER_39_229 ();
 sg13g2_decap_8 FILLER_39_236 ();
 sg13g2_decap_8 FILLER_39_243 ();
 sg13g2_decap_8 FILLER_39_250 ();
 sg13g2_decap_8 FILLER_39_257 ();
 sg13g2_decap_4 FILLER_39_264 ();
 sg13g2_fill_1 FILLER_39_268 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_4 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_fill_2 FILLER_39_338 ();
 sg13g2_decap_8 FILLER_39_354 ();
 sg13g2_decap_8 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_376 ();
 sg13g2_decap_4 FILLER_39_387 ();
 sg13g2_fill_2 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_8 FILLER_39_404 ();
 sg13g2_decap_8 FILLER_39_411 ();
 sg13g2_decap_8 FILLER_39_418 ();
 sg13g2_decap_8 FILLER_39_425 ();
 sg13g2_decap_8 FILLER_39_442 ();
 sg13g2_fill_2 FILLER_39_449 ();
 sg13g2_fill_1 FILLER_39_451 ();
 sg13g2_decap_8 FILLER_39_479 ();
 sg13g2_fill_1 FILLER_39_486 ();
 sg13g2_decap_4 FILLER_39_497 ();
 sg13g2_fill_2 FILLER_39_501 ();
 sg13g2_decap_4 FILLER_39_508 ();
 sg13g2_fill_2 FILLER_39_512 ();
 sg13g2_fill_1 FILLER_39_518 ();
 sg13g2_fill_1 FILLER_39_524 ();
 sg13g2_decap_4 FILLER_39_530 ();
 sg13g2_fill_2 FILLER_39_534 ();
 sg13g2_decap_8 FILLER_39_549 ();
 sg13g2_fill_2 FILLER_39_556 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_fill_1 FILLER_39_574 ();
 sg13g2_fill_1 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_594 ();
 sg13g2_decap_8 FILLER_39_601 ();
 sg13g2_decap_4 FILLER_39_608 ();
 sg13g2_fill_2 FILLER_39_612 ();
 sg13g2_decap_4 FILLER_39_618 ();
 sg13g2_fill_1 FILLER_39_622 ();
 sg13g2_decap_4 FILLER_39_626 ();
 sg13g2_fill_2 FILLER_39_655 ();
 sg13g2_fill_1 FILLER_39_657 ();
 sg13g2_decap_8 FILLER_39_666 ();
 sg13g2_decap_4 FILLER_39_673 ();
 sg13g2_fill_2 FILLER_39_683 ();
 sg13g2_decap_8 FILLER_39_698 ();
 sg13g2_fill_1 FILLER_39_705 ();
 sg13g2_fill_2 FILLER_39_713 ();
 sg13g2_fill_2 FILLER_39_725 ();
 sg13g2_decap_8 FILLER_39_758 ();
 sg13g2_decap_8 FILLER_39_765 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_4 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_39 ();
 sg13g2_fill_2 FILLER_40_45 ();
 sg13g2_fill_1 FILLER_40_47 ();
 sg13g2_decap_8 FILLER_40_57 ();
 sg13g2_decap_8 FILLER_40_64 ();
 sg13g2_decap_8 FILLER_40_71 ();
 sg13g2_fill_2 FILLER_40_78 ();
 sg13g2_fill_1 FILLER_40_80 ();
 sg13g2_fill_1 FILLER_40_112 ();
 sg13g2_fill_2 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_168 ();
 sg13g2_fill_2 FILLER_40_192 ();
 sg13g2_fill_1 FILLER_40_194 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_decap_4 FILLER_40_226 ();
 sg13g2_decap_4 FILLER_40_246 ();
 sg13g2_fill_1 FILLER_40_250 ();
 sg13g2_fill_2 FILLER_40_256 ();
 sg13g2_fill_2 FILLER_40_271 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_292 ();
 sg13g2_fill_2 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_fill_2 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_308 ();
 sg13g2_decap_4 FILLER_40_345 ();
 sg13g2_fill_1 FILLER_40_349 ();
 sg13g2_decap_4 FILLER_40_376 ();
 sg13g2_fill_2 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_4 FILLER_40_434 ();
 sg13g2_fill_2 FILLER_40_459 ();
 sg13g2_fill_1 FILLER_40_461 ();
 sg13g2_decap_4 FILLER_40_470 ();
 sg13g2_fill_1 FILLER_40_474 ();
 sg13g2_fill_1 FILLER_40_483 ();
 sg13g2_fill_1 FILLER_40_492 ();
 sg13g2_decap_8 FILLER_40_506 ();
 sg13g2_fill_1 FILLER_40_513 ();
 sg13g2_fill_2 FILLER_40_519 ();
 sg13g2_fill_1 FILLER_40_529 ();
 sg13g2_fill_1 FILLER_40_587 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_fill_1 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_625 ();
 sg13g2_decap_8 FILLER_40_650 ();
 sg13g2_fill_2 FILLER_40_657 ();
 sg13g2_fill_1 FILLER_40_659 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_fill_2 FILLER_40_679 ();
 sg13g2_fill_1 FILLER_40_681 ();
 sg13g2_fill_1 FILLER_40_697 ();
 sg13g2_fill_2 FILLER_40_711 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_42 ();
 sg13g2_fill_1 FILLER_41_44 ();
 sg13g2_decap_4 FILLER_41_54 ();
 sg13g2_decap_8 FILLER_41_62 ();
 sg13g2_decap_8 FILLER_41_69 ();
 sg13g2_decap_4 FILLER_41_76 ();
 sg13g2_fill_2 FILLER_41_80 ();
 sg13g2_fill_1 FILLER_41_86 ();
 sg13g2_decap_8 FILLER_41_113 ();
 sg13g2_decap_8 FILLER_41_120 ();
 sg13g2_decap_8 FILLER_41_127 ();
 sg13g2_decap_8 FILLER_41_134 ();
 sg13g2_decap_4 FILLER_41_141 ();
 sg13g2_fill_2 FILLER_41_166 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_4 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_205 ();
 sg13g2_decap_8 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_219 ();
 sg13g2_fill_2 FILLER_41_237 ();
 sg13g2_fill_1 FILLER_41_239 ();
 sg13g2_decap_4 FILLER_41_248 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_266 ();
 sg13g2_fill_2 FILLER_41_272 ();
 sg13g2_fill_1 FILLER_41_274 ();
 sg13g2_decap_8 FILLER_41_279 ();
 sg13g2_decap_8 FILLER_41_312 ();
 sg13g2_decap_4 FILLER_41_319 ();
 sg13g2_fill_2 FILLER_41_323 ();
 sg13g2_decap_4 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_349 ();
 sg13g2_decap_4 FILLER_41_359 ();
 sg13g2_fill_2 FILLER_41_363 ();
 sg13g2_decap_4 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_391 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_fill_2 FILLER_41_405 ();
 sg13g2_decap_4 FILLER_41_442 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_fill_2 FILLER_41_478 ();
 sg13g2_fill_1 FILLER_41_480 ();
 sg13g2_decap_8 FILLER_41_500 ();
 sg13g2_decap_8 FILLER_41_507 ();
 sg13g2_fill_2 FILLER_41_514 ();
 sg13g2_fill_2 FILLER_41_529 ();
 sg13g2_fill_1 FILLER_41_540 ();
 sg13g2_decap_8 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_fill_2 FILLER_41_563 ();
 sg13g2_decap_4 FILLER_41_605 ();
 sg13g2_fill_1 FILLER_41_624 ();
 sg13g2_fill_2 FILLER_41_638 ();
 sg13g2_decap_8 FILLER_41_660 ();
 sg13g2_decap_8 FILLER_41_667 ();
 sg13g2_fill_1 FILLER_41_674 ();
 sg13g2_fill_2 FILLER_41_685 ();
 sg13g2_decap_8 FILLER_41_699 ();
 sg13g2_fill_1 FILLER_41_706 ();
 sg13g2_decap_8 FILLER_41_712 ();
 sg13g2_fill_1 FILLER_41_727 ();
 sg13g2_decap_8 FILLER_41_754 ();
 sg13g2_decap_8 FILLER_41_761 ();
 sg13g2_decap_8 FILLER_41_768 ();
 sg13g2_decap_8 FILLER_41_775 ();
 sg13g2_decap_8 FILLER_41_782 ();
 sg13g2_decap_8 FILLER_41_789 ();
 sg13g2_decap_8 FILLER_41_796 ();
 sg13g2_decap_8 FILLER_41_803 ();
 sg13g2_decap_8 FILLER_41_810 ();
 sg13g2_decap_8 FILLER_41_817 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_8 FILLER_41_831 ();
 sg13g2_decap_8 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_fill_2 FILLER_41_859 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_42 ();
 sg13g2_fill_1 FILLER_42_46 ();
 sg13g2_fill_2 FILLER_42_78 ();
 sg13g2_decap_8 FILLER_42_137 ();
 sg13g2_decap_8 FILLER_42_144 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_fill_1 FILLER_42_158 ();
 sg13g2_decap_8 FILLER_42_167 ();
 sg13g2_decap_4 FILLER_42_189 ();
 sg13g2_fill_1 FILLER_42_193 ();
 sg13g2_decap_4 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_decap_8 FILLER_42_215 ();
 sg13g2_fill_2 FILLER_42_222 ();
 sg13g2_fill_2 FILLER_42_231 ();
 sg13g2_fill_1 FILLER_42_233 ();
 sg13g2_decap_8 FILLER_42_239 ();
 sg13g2_decap_4 FILLER_42_246 ();
 sg13g2_decap_8 FILLER_42_255 ();
 sg13g2_decap_4 FILLER_42_267 ();
 sg13g2_fill_2 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_286 ();
 sg13g2_decap_4 FILLER_42_296 ();
 sg13g2_fill_2 FILLER_42_300 ();
 sg13g2_fill_1 FILLER_42_313 ();
 sg13g2_decap_8 FILLER_42_318 ();
 sg13g2_decap_8 FILLER_42_325 ();
 sg13g2_decap_8 FILLER_42_332 ();
 sg13g2_fill_2 FILLER_42_339 ();
 sg13g2_fill_2 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_358 ();
 sg13g2_decap_4 FILLER_42_364 ();
 sg13g2_fill_1 FILLER_42_368 ();
 sg13g2_fill_2 FILLER_42_399 ();
 sg13g2_decap_4 FILLER_42_427 ();
 sg13g2_fill_1 FILLER_42_445 ();
 sg13g2_fill_2 FILLER_42_463 ();
 sg13g2_fill_1 FILLER_42_465 ();
 sg13g2_decap_4 FILLER_42_485 ();
 sg13g2_decap_8 FILLER_42_493 ();
 sg13g2_decap_4 FILLER_42_500 ();
 sg13g2_fill_2 FILLER_42_504 ();
 sg13g2_fill_2 FILLER_42_510 ();
 sg13g2_fill_1 FILLER_42_512 ();
 sg13g2_decap_8 FILLER_42_574 ();
 sg13g2_decap_8 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_588 ();
 sg13g2_fill_2 FILLER_42_595 ();
 sg13g2_fill_2 FILLER_42_614 ();
 sg13g2_fill_1 FILLER_42_616 ();
 sg13g2_decap_8 FILLER_42_626 ();
 sg13g2_fill_1 FILLER_42_633 ();
 sg13g2_fill_2 FILLER_42_649 ();
 sg13g2_fill_2 FILLER_42_677 ();
 sg13g2_fill_1 FILLER_42_692 ();
 sg13g2_decap_8 FILLER_42_698 ();
 sg13g2_fill_1 FILLER_42_705 ();
 sg13g2_decap_8 FILLER_42_710 ();
 sg13g2_decap_8 FILLER_42_717 ();
 sg13g2_decap_8 FILLER_42_724 ();
 sg13g2_decap_4 FILLER_42_731 ();
 sg13g2_fill_1 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_745 ();
 sg13g2_fill_2 FILLER_42_752 ();
 sg13g2_fill_1 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_760 ();
 sg13g2_decap_8 FILLER_42_767 ();
 sg13g2_decap_8 FILLER_42_774 ();
 sg13g2_decap_8 FILLER_42_781 ();
 sg13g2_decap_8 FILLER_42_788 ();
 sg13g2_decap_8 FILLER_42_795 ();
 sg13g2_decap_8 FILLER_42_802 ();
 sg13g2_decap_8 FILLER_42_809 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_42_823 ();
 sg13g2_decap_8 FILLER_42_830 ();
 sg13g2_decap_8 FILLER_42_837 ();
 sg13g2_decap_8 FILLER_42_844 ();
 sg13g2_decap_8 FILLER_42_851 ();
 sg13g2_decap_4 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_4 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_51 ();
 sg13g2_fill_2 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_67 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_fill_2 FILLER_43_94 ();
 sg13g2_fill_2 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_133 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_decap_8 FILLER_43_144 ();
 sg13g2_fill_1 FILLER_43_151 ();
 sg13g2_decap_8 FILLER_43_169 ();
 sg13g2_fill_1 FILLER_43_176 ();
 sg13g2_decap_4 FILLER_43_185 ();
 sg13g2_fill_1 FILLER_43_197 ();
 sg13g2_fill_2 FILLER_43_214 ();
 sg13g2_fill_1 FILLER_43_216 ();
 sg13g2_fill_2 FILLER_43_243 ();
 sg13g2_fill_1 FILLER_43_245 ();
 sg13g2_fill_2 FILLER_43_255 ();
 sg13g2_fill_2 FILLER_43_265 ();
 sg13g2_decap_8 FILLER_43_272 ();
 sg13g2_fill_1 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_317 ();
 sg13g2_fill_2 FILLER_43_338 ();
 sg13g2_fill_1 FILLER_43_340 ();
 sg13g2_fill_2 FILLER_43_349 ();
 sg13g2_decap_4 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_380 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_fill_2 FILLER_43_392 ();
 sg13g2_fill_1 FILLER_43_394 ();
 sg13g2_fill_2 FILLER_43_425 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_4 FILLER_43_448 ();
 sg13g2_fill_1 FILLER_43_452 ();
 sg13g2_decap_8 FILLER_43_457 ();
 sg13g2_fill_2 FILLER_43_464 ();
 sg13g2_fill_1 FILLER_43_466 ();
 sg13g2_fill_2 FILLER_43_493 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_8 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_fill_2 FILLER_43_567 ();
 sg13g2_fill_1 FILLER_43_569 ();
 sg13g2_fill_2 FILLER_43_596 ();
 sg13g2_fill_1 FILLER_43_598 ();
 sg13g2_decap_8 FILLER_43_634 ();
 sg13g2_fill_1 FILLER_43_641 ();
 sg13g2_fill_1 FILLER_43_647 ();
 sg13g2_fill_1 FILLER_43_653 ();
 sg13g2_decap_4 FILLER_43_663 ();
 sg13g2_decap_4 FILLER_43_692 ();
 sg13g2_decap_8 FILLER_43_722 ();
 sg13g2_fill_2 FILLER_43_729 ();
 sg13g2_fill_2 FILLER_43_734 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_decap_8 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_fill_2 FILLER_43_859 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_fill_2 FILLER_44_21 ();
 sg13g2_fill_1 FILLER_44_23 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_fill_1 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_40 ();
 sg13g2_fill_1 FILLER_44_62 ();
 sg13g2_fill_1 FILLER_44_132 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_8 FILLER_44_165 ();
 sg13g2_decap_4 FILLER_44_172 ();
 sg13g2_fill_2 FILLER_44_176 ();
 sg13g2_decap_8 FILLER_44_191 ();
 sg13g2_fill_2 FILLER_44_198 ();
 sg13g2_fill_2 FILLER_44_208 ();
 sg13g2_decap_4 FILLER_44_218 ();
 sg13g2_decap_8 FILLER_44_227 ();
 sg13g2_decap_8 FILLER_44_234 ();
 sg13g2_decap_8 FILLER_44_241 ();
 sg13g2_decap_4 FILLER_44_248 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_4 FILLER_44_277 ();
 sg13g2_fill_2 FILLER_44_290 ();
 sg13g2_decap_4 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_fill_1 FILLER_44_329 ();
 sg13g2_fill_2 FILLER_44_334 ();
 sg13g2_fill_1 FILLER_44_336 ();
 sg13g2_fill_2 FILLER_44_342 ();
 sg13g2_fill_1 FILLER_44_344 ();
 sg13g2_decap_8 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_356 ();
 sg13g2_fill_1 FILLER_44_363 ();
 sg13g2_fill_1 FILLER_44_367 ();
 sg13g2_decap_8 FILLER_44_380 ();
 sg13g2_decap_4 FILLER_44_387 ();
 sg13g2_fill_2 FILLER_44_391 ();
 sg13g2_fill_1 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_432 ();
 sg13g2_decap_8 FILLER_44_488 ();
 sg13g2_decap_4 FILLER_44_495 ();
 sg13g2_fill_1 FILLER_44_499 ();
 sg13g2_fill_2 FILLER_44_539 ();
 sg13g2_decap_8 FILLER_44_545 ();
 sg13g2_decap_8 FILLER_44_552 ();
 sg13g2_decap_8 FILLER_44_559 ();
 sg13g2_fill_2 FILLER_44_566 ();
 sg13g2_fill_1 FILLER_44_568 ();
 sg13g2_decap_8 FILLER_44_597 ();
 sg13g2_fill_2 FILLER_44_604 ();
 sg13g2_fill_1 FILLER_44_606 ();
 sg13g2_fill_1 FILLER_44_672 ();
 sg13g2_fill_2 FILLER_44_713 ();
 sg13g2_fill_1 FILLER_44_715 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_8 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_11 ();
 sg13g2_decap_8 FILLER_45_39 ();
 sg13g2_fill_1 FILLER_45_46 ();
 sg13g2_decap_4 FILLER_45_59 ();
 sg13g2_fill_2 FILLER_45_68 ();
 sg13g2_fill_1 FILLER_45_70 ();
 sg13g2_fill_2 FILLER_45_79 ();
 sg13g2_fill_1 FILLER_45_81 ();
 sg13g2_decap_8 FILLER_45_95 ();
 sg13g2_decap_8 FILLER_45_115 ();
 sg13g2_fill_2 FILLER_45_125 ();
 sg13g2_fill_1 FILLER_45_127 ();
 sg13g2_fill_2 FILLER_45_136 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_decap_4 FILLER_45_143 ();
 sg13g2_fill_2 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_fill_1 FILLER_45_182 ();
 sg13g2_fill_2 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_211 ();
 sg13g2_decap_4 FILLER_45_218 ();
 sg13g2_fill_2 FILLER_45_229 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_fill_2 FILLER_45_250 ();
 sg13g2_decap_4 FILLER_45_268 ();
 sg13g2_fill_1 FILLER_45_272 ();
 sg13g2_fill_2 FILLER_45_325 ();
 sg13g2_fill_1 FILLER_45_327 ();
 sg13g2_fill_2 FILLER_45_344 ();
 sg13g2_decap_4 FILLER_45_357 ();
 sg13g2_fill_1 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_391 ();
 sg13g2_fill_2 FILLER_45_398 ();
 sg13g2_fill_1 FILLER_45_400 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_fill_2 FILLER_45_409 ();
 sg13g2_decap_4 FILLER_45_419 ();
 sg13g2_fill_1 FILLER_45_453 ();
 sg13g2_decap_8 FILLER_45_459 ();
 sg13g2_fill_1 FILLER_45_491 ();
 sg13g2_fill_2 FILLER_45_517 ();
 sg13g2_fill_1 FILLER_45_519 ();
 sg13g2_fill_2 FILLER_45_528 ();
 sg13g2_fill_1 FILLER_45_530 ();
 sg13g2_fill_2 FILLER_45_567 ();
 sg13g2_fill_1 FILLER_45_569 ();
 sg13g2_fill_2 FILLER_45_592 ();
 sg13g2_fill_1 FILLER_45_594 ();
 sg13g2_decap_4 FILLER_45_610 ();
 sg13g2_fill_2 FILLER_45_620 ();
 sg13g2_decap_8 FILLER_45_640 ();
 sg13g2_fill_1 FILLER_45_647 ();
 sg13g2_fill_1 FILLER_45_653 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_fill_2 FILLER_45_672 ();
 sg13g2_fill_2 FILLER_45_693 ();
 sg13g2_fill_1 FILLER_45_695 ();
 sg13g2_fill_2 FILLER_45_701 ();
 sg13g2_fill_1 FILLER_45_703 ();
 sg13g2_decap_8 FILLER_45_775 ();
 sg13g2_decap_8 FILLER_45_782 ();
 sg13g2_decap_8 FILLER_45_789 ();
 sg13g2_decap_8 FILLER_45_796 ();
 sg13g2_decap_8 FILLER_45_803 ();
 sg13g2_decap_8 FILLER_45_810 ();
 sg13g2_decap_8 FILLER_45_817 ();
 sg13g2_decap_8 FILLER_45_824 ();
 sg13g2_decap_8 FILLER_45_831 ();
 sg13g2_decap_8 FILLER_45_838 ();
 sg13g2_decap_8 FILLER_45_845 ();
 sg13g2_decap_8 FILLER_45_852 ();
 sg13g2_fill_2 FILLER_45_859 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_28 ();
 sg13g2_decap_4 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_116 ();
 sg13g2_fill_1 FILLER_46_118 ();
 sg13g2_decap_8 FILLER_46_137 ();
 sg13g2_fill_2 FILLER_46_144 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_168 ();
 sg13g2_decap_4 FILLER_46_175 ();
 sg13g2_fill_1 FILLER_46_192 ();
 sg13g2_decap_8 FILLER_46_213 ();
 sg13g2_fill_1 FILLER_46_225 ();
 sg13g2_decap_4 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_254 ();
 sg13g2_fill_1 FILLER_46_256 ();
 sg13g2_decap_4 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_274 ();
 sg13g2_fill_2 FILLER_46_289 ();
 sg13g2_fill_1 FILLER_46_305 ();
 sg13g2_decap_4 FILLER_46_315 ();
 sg13g2_decap_4 FILLER_46_328 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_fill_1 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_decap_4 FILLER_46_382 ();
 sg13g2_fill_1 FILLER_46_386 ();
 sg13g2_fill_2 FILLER_46_391 ();
 sg13g2_fill_2 FILLER_46_419 ();
 sg13g2_decap_8 FILLER_46_442 ();
 sg13g2_decap_4 FILLER_46_449 ();
 sg13g2_fill_2 FILLER_46_453 ();
 sg13g2_decap_8 FILLER_46_459 ();
 sg13g2_decap_4 FILLER_46_466 ();
 sg13g2_decap_8 FILLER_46_480 ();
 sg13g2_fill_2 FILLER_46_487 ();
 sg13g2_fill_1 FILLER_46_500 ();
 sg13g2_fill_2 FILLER_46_504 ();
 sg13g2_fill_2 FILLER_46_519 ();
 sg13g2_fill_1 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_531 ();
 sg13g2_decap_4 FILLER_46_538 ();
 sg13g2_decap_4 FILLER_46_553 ();
 sg13g2_fill_2 FILLER_46_557 ();
 sg13g2_fill_2 FILLER_46_563 ();
 sg13g2_fill_1 FILLER_46_575 ();
 sg13g2_fill_1 FILLER_46_580 ();
 sg13g2_decap_4 FILLER_46_585 ();
 sg13g2_fill_1 FILLER_46_589 ();
 sg13g2_fill_1 FILLER_46_594 ();
 sg13g2_decap_4 FILLER_46_604 ();
 sg13g2_fill_2 FILLER_46_608 ();
 sg13g2_fill_2 FILLER_46_637 ();
 sg13g2_fill_1 FILLER_46_639 ();
 sg13g2_decap_8 FILLER_46_690 ();
 sg13g2_fill_2 FILLER_46_697 ();
 sg13g2_fill_2 FILLER_46_716 ();
 sg13g2_fill_2 FILLER_46_726 ();
 sg13g2_fill_2 FILLER_46_753 ();
 sg13g2_fill_1 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_773 ();
 sg13g2_decap_8 FILLER_46_780 ();
 sg13g2_decap_8 FILLER_46_787 ();
 sg13g2_decap_8 FILLER_46_794 ();
 sg13g2_decap_8 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_4 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_27 ();
 sg13g2_fill_2 FILLER_47_42 ();
 sg13g2_fill_1 FILLER_47_52 ();
 sg13g2_fill_1 FILLER_47_57 ();
 sg13g2_fill_2 FILLER_47_83 ();
 sg13g2_fill_1 FILLER_47_85 ();
 sg13g2_decap_4 FILLER_47_95 ();
 sg13g2_fill_2 FILLER_47_99 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_fill_2 FILLER_47_131 ();
 sg13g2_fill_1 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_138 ();
 sg13g2_fill_2 FILLER_47_169 ();
 sg13g2_fill_1 FILLER_47_171 ();
 sg13g2_decap_8 FILLER_47_180 ();
 sg13g2_fill_2 FILLER_47_187 ();
 sg13g2_decap_8 FILLER_47_199 ();
 sg13g2_decap_8 FILLER_47_206 ();
 sg13g2_decap_8 FILLER_47_213 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_4 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_decap_4 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_fill_1 FILLER_47_314 ();
 sg13g2_fill_2 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_4 FILLER_47_371 ();
 sg13g2_fill_2 FILLER_47_375 ();
 sg13g2_decap_8 FILLER_47_421 ();
 sg13g2_decap_4 FILLER_47_536 ();
 sg13g2_decap_8 FILLER_47_596 ();
 sg13g2_decap_8 FILLER_47_603 ();
 sg13g2_fill_1 FILLER_47_610 ();
 sg13g2_decap_8 FILLER_47_629 ();
 sg13g2_decap_4 FILLER_47_636 ();
 sg13g2_fill_2 FILLER_47_640 ();
 sg13g2_decap_8 FILLER_47_685 ();
 sg13g2_fill_2 FILLER_47_692 ();
 sg13g2_fill_1 FILLER_47_694 ();
 sg13g2_fill_1 FILLER_47_712 ();
 sg13g2_fill_1 FILLER_47_718 ();
 sg13g2_decap_8 FILLER_47_724 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_15 ();
 sg13g2_fill_2 FILLER_48_22 ();
 sg13g2_fill_1 FILLER_48_24 ();
 sg13g2_fill_2 FILLER_48_39 ();
 sg13g2_fill_1 FILLER_48_41 ();
 sg13g2_decap_8 FILLER_48_47 ();
 sg13g2_decap_4 FILLER_48_54 ();
 sg13g2_fill_2 FILLER_48_58 ();
 sg13g2_decap_4 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_67 ();
 sg13g2_decap_8 FILLER_48_102 ();
 sg13g2_fill_2 FILLER_48_109 ();
 sg13g2_fill_1 FILLER_48_111 ();
 sg13g2_decap_8 FILLER_48_137 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_fill_2 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_166 ();
 sg13g2_decap_4 FILLER_48_173 ();
 sg13g2_fill_1 FILLER_48_177 ();
 sg13g2_decap_4 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_192 ();
 sg13g2_fill_2 FILLER_48_205 ();
 sg13g2_decap_8 FILLER_48_236 ();
 sg13g2_fill_1 FILLER_48_243 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_2 FILLER_48_296 ();
 sg13g2_decap_8 FILLER_48_331 ();
 sg13g2_decap_8 FILLER_48_338 ();
 sg13g2_decap_4 FILLER_48_345 ();
 sg13g2_decap_4 FILLER_48_361 ();
 sg13g2_fill_1 FILLER_48_365 ();
 sg13g2_decap_4 FILLER_48_382 ();
 sg13g2_decap_4 FILLER_48_421 ();
 sg13g2_decap_4 FILLER_48_441 ();
 sg13g2_fill_1 FILLER_48_445 ();
 sg13g2_decap_8 FILLER_48_450 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_fill_2 FILLER_48_483 ();
 sg13g2_fill_1 FILLER_48_485 ();
 sg13g2_decap_8 FILLER_48_502 ();
 sg13g2_decap_4 FILLER_48_513 ();
 sg13g2_fill_2 FILLER_48_517 ();
 sg13g2_decap_8 FILLER_48_533 ();
 sg13g2_fill_2 FILLER_48_540 ();
 sg13g2_decap_8 FILLER_48_550 ();
 sg13g2_fill_2 FILLER_48_562 ();
 sg13g2_fill_1 FILLER_48_582 ();
 sg13g2_decap_4 FILLER_48_635 ();
 sg13g2_decap_4 FILLER_48_653 ();
 sg13g2_fill_2 FILLER_48_657 ();
 sg13g2_decap_4 FILLER_48_674 ();
 sg13g2_fill_2 FILLER_48_678 ();
 sg13g2_fill_1 FILLER_48_683 ();
 sg13g2_fill_1 FILLER_48_696 ();
 sg13g2_fill_1 FILLER_48_710 ();
 sg13g2_decap_8 FILLER_48_752 ();
 sg13g2_fill_2 FILLER_48_759 ();
 sg13g2_fill_1 FILLER_48_761 ();
 sg13g2_decap_8 FILLER_48_788 ();
 sg13g2_decap_8 FILLER_48_795 ();
 sg13g2_decap_8 FILLER_48_802 ();
 sg13g2_decap_8 FILLER_48_809 ();
 sg13g2_decap_8 FILLER_48_816 ();
 sg13g2_decap_8 FILLER_48_823 ();
 sg13g2_decap_8 FILLER_48_830 ();
 sg13g2_decap_8 FILLER_48_837 ();
 sg13g2_decap_8 FILLER_48_844 ();
 sg13g2_decap_8 FILLER_48_851 ();
 sg13g2_decap_4 FILLER_48_858 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_2 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_decap_4 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_fill_2 FILLER_49_116 ();
 sg13g2_fill_2 FILLER_49_122 ();
 sg13g2_fill_1 FILLER_49_124 ();
 sg13g2_decap_4 FILLER_49_138 ();
 sg13g2_fill_2 FILLER_49_152 ();
 sg13g2_decap_4 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_163 ();
 sg13g2_decap_4 FILLER_49_176 ();
 sg13g2_decap_8 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_fill_2 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_226 ();
 sg13g2_decap_4 FILLER_49_233 ();
 sg13g2_fill_2 FILLER_49_237 ();
 sg13g2_decap_8 FILLER_49_261 ();
 sg13g2_decap_8 FILLER_49_268 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_289 ();
 sg13g2_fill_1 FILLER_49_296 ();
 sg13g2_fill_1 FILLER_49_311 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_decap_8 FILLER_49_328 ();
 sg13g2_fill_2 FILLER_49_335 ();
 sg13g2_decap_4 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_fill_1 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_380 ();
 sg13g2_fill_2 FILLER_49_387 ();
 sg13g2_fill_1 FILLER_49_389 ();
 sg13g2_fill_1 FILLER_49_409 ();
 sg13g2_decap_8 FILLER_49_418 ();
 sg13g2_fill_1 FILLER_49_425 ();
 sg13g2_fill_2 FILLER_49_431 ();
 sg13g2_fill_1 FILLER_49_433 ();
 sg13g2_fill_2 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_461 ();
 sg13g2_fill_2 FILLER_49_483 ();
 sg13g2_fill_1 FILLER_49_485 ();
 sg13g2_fill_2 FILLER_49_496 ();
 sg13g2_fill_1 FILLER_49_498 ();
 sg13g2_fill_2 FILLER_49_512 ();
 sg13g2_fill_1 FILLER_49_514 ();
 sg13g2_decap_8 FILLER_49_541 ();
 sg13g2_fill_2 FILLER_49_548 ();
 sg13g2_fill_1 FILLER_49_550 ();
 sg13g2_fill_1 FILLER_49_559 ();
 sg13g2_fill_2 FILLER_49_574 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_fill_2 FILLER_49_593 ();
 sg13g2_decap_4 FILLER_49_605 ();
 sg13g2_fill_2 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_615 ();
 sg13g2_fill_1 FILLER_49_622 ();
 sg13g2_decap_4 FILLER_49_627 ();
 sg13g2_fill_2 FILLER_49_631 ();
 sg13g2_fill_1 FILLER_49_657 ();
 sg13g2_fill_2 FILLER_49_721 ();
 sg13g2_fill_2 FILLER_49_746 ();
 sg13g2_decap_8 FILLER_49_757 ();
 sg13g2_fill_1 FILLER_49_764 ();
 sg13g2_decap_8 FILLER_49_778 ();
 sg13g2_fill_2 FILLER_49_785 ();
 sg13g2_decap_8 FILLER_49_813 ();
 sg13g2_decap_8 FILLER_49_820 ();
 sg13g2_decap_8 FILLER_49_827 ();
 sg13g2_decap_8 FILLER_49_834 ();
 sg13g2_decap_8 FILLER_49_841 ();
 sg13g2_decap_8 FILLER_49_848 ();
 sg13g2_decap_8 FILLER_49_855 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_1 FILLER_50_41 ();
 sg13g2_decap_8 FILLER_50_47 ();
 sg13g2_decap_8 FILLER_50_58 ();
 sg13g2_decap_4 FILLER_50_65 ();
 sg13g2_fill_2 FILLER_50_69 ();
 sg13g2_decap_8 FILLER_50_79 ();
 sg13g2_fill_2 FILLER_50_86 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_117 ();
 sg13g2_decap_8 FILLER_50_124 ();
 sg13g2_decap_4 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_decap_4 FILLER_50_161 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_fill_1 FILLER_50_190 ();
 sg13g2_decap_4 FILLER_50_205 ();
 sg13g2_fill_1 FILLER_50_232 ();
 sg13g2_fill_1 FILLER_50_247 ();
 sg13g2_decap_8 FILLER_50_262 ();
 sg13g2_fill_2 FILLER_50_280 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_decap_4 FILLER_50_366 ();
 sg13g2_fill_1 FILLER_50_430 ();
 sg13g2_decap_4 FILLER_50_454 ();
 sg13g2_decap_4 FILLER_50_463 ();
 sg13g2_fill_1 FILLER_50_467 ();
 sg13g2_decap_8 FILLER_50_473 ();
 sg13g2_fill_2 FILLER_50_480 ();
 sg13g2_decap_8 FILLER_50_503 ();
 sg13g2_fill_1 FILLER_50_510 ();
 sg13g2_decap_8 FILLER_50_515 ();
 sg13g2_fill_2 FILLER_50_522 ();
 sg13g2_fill_1 FILLER_50_524 ();
 sg13g2_decap_4 FILLER_50_540 ();
 sg13g2_fill_1 FILLER_50_544 ();
 sg13g2_decap_4 FILLER_50_561 ();
 sg13g2_fill_1 FILLER_50_565 ();
 sg13g2_fill_2 FILLER_50_577 ();
 sg13g2_fill_2 FILLER_50_588 ();
 sg13g2_fill_1 FILLER_50_590 ();
 sg13g2_fill_2 FILLER_50_611 ();
 sg13g2_fill_2 FILLER_50_623 ();
 sg13g2_fill_1 FILLER_50_625 ();
 sg13g2_decap_8 FILLER_50_634 ();
 sg13g2_fill_1 FILLER_50_641 ();
 sg13g2_decap_8 FILLER_50_655 ();
 sg13g2_fill_2 FILLER_50_662 ();
 sg13g2_fill_1 FILLER_50_664 ();
 sg13g2_fill_1 FILLER_50_684 ();
 sg13g2_decap_8 FILLER_50_711 ();
 sg13g2_fill_1 FILLER_50_718 ();
 sg13g2_fill_1 FILLER_50_729 ();
 sg13g2_decap_4 FILLER_50_771 ();
 sg13g2_fill_2 FILLER_50_775 ();
 sg13g2_fill_2 FILLER_50_796 ();
 sg13g2_fill_1 FILLER_50_798 ();
 sg13g2_decap_8 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_833 ();
 sg13g2_decap_8 FILLER_50_840 ();
 sg13g2_decap_8 FILLER_50_847 ();
 sg13g2_decap_8 FILLER_50_854 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_51_40 ();
 sg13g2_fill_1 FILLER_51_47 ();
 sg13g2_fill_1 FILLER_51_60 ();
 sg13g2_decap_4 FILLER_51_86 ();
 sg13g2_fill_1 FILLER_51_90 ();
 sg13g2_fill_2 FILLER_51_95 ();
 sg13g2_fill_1 FILLER_51_97 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_decap_4 FILLER_51_120 ();
 sg13g2_decap_8 FILLER_51_153 ();
 sg13g2_fill_2 FILLER_51_165 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_decap_8 FILLER_51_173 ();
 sg13g2_decap_4 FILLER_51_180 ();
 sg13g2_fill_1 FILLER_51_192 ();
 sg13g2_decap_8 FILLER_51_207 ();
 sg13g2_decap_4 FILLER_51_214 ();
 sg13g2_fill_2 FILLER_51_218 ();
 sg13g2_fill_2 FILLER_51_225 ();
 sg13g2_fill_1 FILLER_51_227 ();
 sg13g2_decap_8 FILLER_51_231 ();
 sg13g2_decap_8 FILLER_51_238 ();
 sg13g2_decap_4 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_263 ();
 sg13g2_decap_8 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_307 ();
 sg13g2_decap_8 FILLER_51_328 ();
 sg13g2_fill_1 FILLER_51_335 ();
 sg13g2_decap_8 FILLER_51_340 ();
 sg13g2_decap_4 FILLER_51_347 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_fill_2 FILLER_51_377 ();
 sg13g2_fill_1 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_401 ();
 sg13g2_decap_8 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_51_419 ();
 sg13g2_decap_8 FILLER_51_438 ();
 sg13g2_fill_1 FILLER_51_445 ();
 sg13g2_decap_8 FILLER_51_469 ();
 sg13g2_decap_4 FILLER_51_476 ();
 sg13g2_fill_2 FILLER_51_480 ();
 sg13g2_fill_2 FILLER_51_508 ();
 sg13g2_fill_1 FILLER_51_510 ();
 sg13g2_decap_8 FILLER_51_521 ();
 sg13g2_fill_1 FILLER_51_533 ();
 sg13g2_decap_8 FILLER_51_538 ();
 sg13g2_decap_4 FILLER_51_545 ();
 sg13g2_fill_1 FILLER_51_575 ();
 sg13g2_decap_8 FILLER_51_602 ();
 sg13g2_decap_4 FILLER_51_609 ();
 sg13g2_fill_1 FILLER_51_656 ();
 sg13g2_decap_8 FILLER_51_688 ();
 sg13g2_fill_2 FILLER_51_695 ();
 sg13g2_decap_8 FILLER_51_706 ();
 sg13g2_decap_4 FILLER_51_713 ();
 sg13g2_fill_2 FILLER_51_717 ();
 sg13g2_fill_2 FILLER_51_757 ();
 sg13g2_decap_4 FILLER_51_781 ();
 sg13g2_fill_1 FILLER_51_789 ();
 sg13g2_fill_2 FILLER_51_795 ();
 sg13g2_fill_1 FILLER_51_800 ();
 sg13g2_decap_8 FILLER_51_827 ();
 sg13g2_decap_8 FILLER_51_834 ();
 sg13g2_decap_8 FILLER_51_841 ();
 sg13g2_decap_8 FILLER_51_848 ();
 sg13g2_decap_8 FILLER_51_855 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_22 ();
 sg13g2_fill_2 FILLER_52_36 ();
 sg13g2_fill_1 FILLER_52_38 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_decap_4 FILLER_52_70 ();
 sg13g2_fill_2 FILLER_52_74 ();
 sg13g2_fill_1 FILLER_52_89 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_fill_1 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_129 ();
 sg13g2_decap_8 FILLER_52_136 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_fill_2 FILLER_52_158 ();
 sg13g2_decap_4 FILLER_52_172 ();
 sg13g2_fill_2 FILLER_52_176 ();
 sg13g2_decap_4 FILLER_52_199 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_decap_4 FILLER_52_210 ();
 sg13g2_fill_1 FILLER_52_214 ();
 sg13g2_decap_8 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_253 ();
 sg13g2_fill_2 FILLER_52_280 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_1 FILLER_52_319 ();
 sg13g2_decap_8 FILLER_52_334 ();
 sg13g2_decap_4 FILLER_52_341 ();
 sg13g2_fill_2 FILLER_52_350 ();
 sg13g2_fill_1 FILLER_52_352 ();
 sg13g2_decap_4 FILLER_52_359 ();
 sg13g2_decap_8 FILLER_52_372 ();
 sg13g2_decap_8 FILLER_52_379 ();
 sg13g2_fill_1 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_52_409 ();
 sg13g2_decap_8 FILLER_52_416 ();
 sg13g2_decap_8 FILLER_52_423 ();
 sg13g2_decap_4 FILLER_52_430 ();
 sg13g2_decap_4 FILLER_52_438 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_decap_8 FILLER_52_448 ();
 sg13g2_decap_4 FILLER_52_455 ();
 sg13g2_fill_2 FILLER_52_459 ();
 sg13g2_decap_4 FILLER_52_508 ();
 sg13g2_fill_2 FILLER_52_520 ();
 sg13g2_fill_1 FILLER_52_522 ();
 sg13g2_decap_4 FILLER_52_554 ();
 sg13g2_fill_2 FILLER_52_558 ();
 sg13g2_decap_8 FILLER_52_564 ();
 sg13g2_decap_8 FILLER_52_571 ();
 sg13g2_fill_1 FILLER_52_583 ();
 sg13g2_decap_8 FILLER_52_605 ();
 sg13g2_fill_1 FILLER_52_620 ();
 sg13g2_decap_4 FILLER_52_629 ();
 sg13g2_fill_1 FILLER_52_633 ();
 sg13g2_decap_4 FILLER_52_637 ();
 sg13g2_fill_2 FILLER_52_641 ();
 sg13g2_decap_8 FILLER_52_653 ();
 sg13g2_decap_8 FILLER_52_660 ();
 sg13g2_fill_1 FILLER_52_667 ();
 sg13g2_decap_8 FILLER_52_672 ();
 sg13g2_decap_8 FILLER_52_679 ();
 sg13g2_fill_1 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_691 ();
 sg13g2_fill_2 FILLER_52_698 ();
 sg13g2_decap_8 FILLER_52_726 ();
 sg13g2_fill_1 FILLER_52_733 ();
 sg13g2_decap_8 FILLER_52_757 ();
 sg13g2_fill_1 FILLER_52_764 ();
 sg13g2_decap_4 FILLER_52_770 ();
 sg13g2_fill_1 FILLER_52_774 ();
 sg13g2_decap_4 FILLER_52_805 ();
 sg13g2_fill_2 FILLER_52_809 ();
 sg13g2_decap_8 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_822 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_decap_8 FILLER_52_836 ();
 sg13g2_decap_8 FILLER_52_843 ();
 sg13g2_decap_8 FILLER_52_850 ();
 sg13g2_decap_4 FILLER_52_857 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_15 ();
 sg13g2_decap_4 FILLER_53_21 ();
 sg13g2_fill_2 FILLER_53_25 ();
 sg13g2_fill_2 FILLER_53_67 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_86 ();
 sg13g2_fill_2 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_120 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_166 ();
 sg13g2_decap_8 FILLER_53_173 ();
 sg13g2_decap_4 FILLER_53_180 ();
 sg13g2_fill_1 FILLER_53_184 ();
 sg13g2_fill_1 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_229 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_decap_8 FILLER_53_253 ();
 sg13g2_decap_8 FILLER_53_271 ();
 sg13g2_decap_8 FILLER_53_278 ();
 sg13g2_fill_2 FILLER_53_285 ();
 sg13g2_fill_1 FILLER_53_287 ();
 sg13g2_decap_4 FILLER_53_292 ();
 sg13g2_decap_4 FILLER_53_301 ();
 sg13g2_fill_1 FILLER_53_305 ();
 sg13g2_fill_2 FILLER_53_337 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_356 ();
 sg13g2_fill_1 FILLER_53_358 ();
 sg13g2_decap_4 FILLER_53_384 ();
 sg13g2_decap_8 FILLER_53_455 ();
 sg13g2_fill_2 FILLER_53_462 ();
 sg13g2_fill_2 FILLER_53_472 ();
 sg13g2_fill_2 FILLER_53_477 ();
 sg13g2_fill_1 FILLER_53_479 ();
 sg13g2_fill_2 FILLER_53_487 ();
 sg13g2_fill_1 FILLER_53_489 ();
 sg13g2_fill_2 FILLER_53_510 ();
 sg13g2_fill_1 FILLER_53_512 ();
 sg13g2_fill_2 FILLER_53_518 ();
 sg13g2_decap_8 FILLER_53_524 ();
 sg13g2_decap_8 FILLER_53_531 ();
 sg13g2_fill_2 FILLER_53_538 ();
 sg13g2_decap_4 FILLER_53_557 ();
 sg13g2_fill_1 FILLER_53_561 ();
 sg13g2_decap_4 FILLER_53_566 ();
 sg13g2_decap_4 FILLER_53_575 ();
 sg13g2_decap_8 FILLER_53_622 ();
 sg13g2_decap_4 FILLER_53_633 ();
 sg13g2_decap_4 FILLER_53_643 ();
 sg13g2_decap_4 FILLER_53_658 ();
 sg13g2_decap_8 FILLER_53_672 ();
 sg13g2_fill_2 FILLER_53_679 ();
 sg13g2_fill_1 FILLER_53_681 ();
 sg13g2_fill_1 FILLER_53_705 ();
 sg13g2_decap_8 FILLER_53_728 ();
 sg13g2_decap_8 FILLER_53_735 ();
 sg13g2_fill_2 FILLER_53_742 ();
 sg13g2_decap_8 FILLER_53_758 ();
 sg13g2_decap_8 FILLER_53_765 ();
 sg13g2_decap_4 FILLER_53_772 ();
 sg13g2_fill_1 FILLER_53_776 ();
 sg13g2_decap_8 FILLER_53_789 ();
 sg13g2_decap_4 FILLER_53_796 ();
 sg13g2_decap_8 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_833 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_53_847 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_fill_1 FILLER_54_26 ();
 sg13g2_decap_8 FILLER_54_51 ();
 sg13g2_decap_8 FILLER_54_58 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_4 FILLER_54_84 ();
 sg13g2_fill_2 FILLER_54_88 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_4 FILLER_54_105 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_fill_2 FILLER_54_114 ();
 sg13g2_decap_8 FILLER_54_124 ();
 sg13g2_fill_2 FILLER_54_131 ();
 sg13g2_decap_4 FILLER_54_141 ();
 sg13g2_fill_2 FILLER_54_145 ();
 sg13g2_decap_4 FILLER_54_156 ();
 sg13g2_decap_4 FILLER_54_186 ();
 sg13g2_decap_8 FILLER_54_193 ();
 sg13g2_fill_2 FILLER_54_200 ();
 sg13g2_decap_8 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_249 ();
 sg13g2_decap_8 FILLER_54_256 ();
 sg13g2_fill_1 FILLER_54_263 ();
 sg13g2_decap_4 FILLER_54_272 ();
 sg13g2_fill_1 FILLER_54_276 ();
 sg13g2_fill_1 FILLER_54_289 ();
 sg13g2_decap_8 FILLER_54_298 ();
 sg13g2_decap_4 FILLER_54_324 ();
 sg13g2_fill_2 FILLER_54_337 ();
 sg13g2_fill_1 FILLER_54_339 ();
 sg13g2_fill_2 FILLER_54_345 ();
 sg13g2_decap_8 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_fill_2 FILLER_54_377 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_54_422 ();
 sg13g2_decap_4 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_54_433 ();
 sg13g2_fill_1 FILLER_54_470 ();
 sg13g2_fill_2 FILLER_54_499 ();
 sg13g2_fill_2 FILLER_54_557 ();
 sg13g2_decap_8 FILLER_54_580 ();
 sg13g2_decap_8 FILLER_54_587 ();
 sg13g2_decap_8 FILLER_54_594 ();
 sg13g2_decap_4 FILLER_54_601 ();
 sg13g2_fill_2 FILLER_54_605 ();
 sg13g2_decap_8 FILLER_54_611 ();
 sg13g2_fill_2 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_656 ();
 sg13g2_decap_4 FILLER_54_697 ();
 sg13g2_fill_2 FILLER_54_736 ();
 sg13g2_fill_1 FILLER_54_738 ();
 sg13g2_decap_8 FILLER_54_754 ();
 sg13g2_decap_4 FILLER_54_761 ();
 sg13g2_fill_2 FILLER_54_765 ();
 sg13g2_fill_2 FILLER_54_788 ();
 sg13g2_fill_2 FILLER_54_803 ();
 sg13g2_decap_8 FILLER_54_831 ();
 sg13g2_decap_8 FILLER_54_838 ();
 sg13g2_decap_8 FILLER_54_845 ();
 sg13g2_decap_8 FILLER_54_852 ();
 sg13g2_fill_2 FILLER_54_859 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_fill_1 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_43 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_decap_8 FILLER_55_59 ();
 sg13g2_decap_8 FILLER_55_66 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_fill_2 FILLER_55_98 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_decap_8 FILLER_55_171 ();
 sg13g2_decap_4 FILLER_55_178 ();
 sg13g2_fill_1 FILLER_55_182 ();
 sg13g2_fill_1 FILLER_55_187 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_fill_2 FILLER_55_232 ();
 sg13g2_fill_1 FILLER_55_234 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_fill_2 FILLER_55_252 ();
 sg13g2_fill_2 FILLER_55_272 ();
 sg13g2_fill_2 FILLER_55_282 ();
 sg13g2_fill_1 FILLER_55_284 ();
 sg13g2_decap_8 FILLER_55_298 ();
 sg13g2_fill_2 FILLER_55_305 ();
 sg13g2_fill_2 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_355 ();
 sg13g2_decap_8 FILLER_55_372 ();
 sg13g2_fill_2 FILLER_55_379 ();
 sg13g2_decap_8 FILLER_55_434 ();
 sg13g2_decap_4 FILLER_55_441 ();
 sg13g2_fill_1 FILLER_55_445 ();
 sg13g2_decap_8 FILLER_55_450 ();
 sg13g2_fill_1 FILLER_55_482 ();
 sg13g2_decap_8 FILLER_55_486 ();
 sg13g2_fill_2 FILLER_55_493 ();
 sg13g2_fill_1 FILLER_55_495 ();
 sg13g2_decap_8 FILLER_55_501 ();
 sg13g2_decap_4 FILLER_55_508 ();
 sg13g2_fill_2 FILLER_55_512 ();
 sg13g2_decap_8 FILLER_55_517 ();
 sg13g2_decap_8 FILLER_55_524 ();
 sg13g2_decap_8 FILLER_55_531 ();
 sg13g2_decap_4 FILLER_55_538 ();
 sg13g2_fill_2 FILLER_55_542 ();
 sg13g2_decap_8 FILLER_55_552 ();
 sg13g2_decap_8 FILLER_55_559 ();
 sg13g2_decap_8 FILLER_55_579 ();
 sg13g2_decap_4 FILLER_55_586 ();
 sg13g2_decap_8 FILLER_55_613 ();
 sg13g2_fill_1 FILLER_55_620 ();
 sg13g2_fill_2 FILLER_55_626 ();
 sg13g2_fill_2 FILLER_55_647 ();
 sg13g2_fill_1 FILLER_55_649 ();
 sg13g2_fill_2 FILLER_55_667 ();
 sg13g2_fill_2 FILLER_55_673 ();
 sg13g2_decap_4 FILLER_55_684 ();
 sg13g2_fill_2 FILLER_55_688 ();
 sg13g2_decap_8 FILLER_55_695 ();
 sg13g2_decap_8 FILLER_55_702 ();
 sg13g2_decap_4 FILLER_55_709 ();
 sg13g2_fill_2 FILLER_55_713 ();
 sg13g2_decap_8 FILLER_55_732 ();
 sg13g2_fill_2 FILLER_55_739 ();
 sg13g2_decap_4 FILLER_55_754 ();
 sg13g2_fill_1 FILLER_55_787 ();
 sg13g2_fill_2 FILLER_55_796 ();
 sg13g2_fill_1 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_825 ();
 sg13g2_decap_8 FILLER_55_832 ();
 sg13g2_decap_8 FILLER_55_839 ();
 sg13g2_decap_8 FILLER_55_846 ();
 sg13g2_decap_8 FILLER_55_853 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_47 ();
 sg13g2_fill_2 FILLER_56_62 ();
 sg13g2_fill_1 FILLER_56_64 ();
 sg13g2_decap_8 FILLER_56_86 ();
 sg13g2_fill_2 FILLER_56_93 ();
 sg13g2_fill_1 FILLER_56_110 ();
 sg13g2_decap_8 FILLER_56_117 ();
 sg13g2_fill_2 FILLER_56_124 ();
 sg13g2_fill_1 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_144 ();
 sg13g2_decap_4 FILLER_56_173 ();
 sg13g2_fill_1 FILLER_56_177 ();
 sg13g2_decap_4 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_190 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_fill_1 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_213 ();
 sg13g2_decap_8 FILLER_56_220 ();
 sg13g2_decap_8 FILLER_56_227 ();
 sg13g2_fill_1 FILLER_56_234 ();
 sg13g2_fill_1 FILLER_56_243 ();
 sg13g2_decap_8 FILLER_56_253 ();
 sg13g2_decap_8 FILLER_56_260 ();
 sg13g2_decap_4 FILLER_56_270 ();
 sg13g2_decap_8 FILLER_56_283 ();
 sg13g2_decap_8 FILLER_56_290 ();
 sg13g2_fill_1 FILLER_56_297 ();
 sg13g2_decap_8 FILLER_56_319 ();
 sg13g2_decap_4 FILLER_56_326 ();
 sg13g2_fill_1 FILLER_56_330 ();
 sg13g2_decap_8 FILLER_56_348 ();
 sg13g2_fill_2 FILLER_56_355 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_fill_2 FILLER_56_371 ();
 sg13g2_fill_1 FILLER_56_373 ();
 sg13g2_decap_4 FILLER_56_379 ();
 sg13g2_fill_2 FILLER_56_383 ();
 sg13g2_decap_4 FILLER_56_402 ();
 sg13g2_fill_1 FILLER_56_406 ();
 sg13g2_fill_2 FILLER_56_421 ();
 sg13g2_fill_1 FILLER_56_449 ();
 sg13g2_fill_2 FILLER_56_476 ();
 sg13g2_fill_1 FILLER_56_478 ();
 sg13g2_fill_1 FILLER_56_507 ();
 sg13g2_fill_2 FILLER_56_511 ();
 sg13g2_fill_1 FILLER_56_517 ();
 sg13g2_decap_4 FILLER_56_533 ();
 sg13g2_fill_2 FILLER_56_537 ();
 sg13g2_fill_2 FILLER_56_583 ();
 sg13g2_fill_2 FILLER_56_655 ();
 sg13g2_decap_8 FILLER_56_669 ();
 sg13g2_decap_4 FILLER_56_676 ();
 sg13g2_fill_2 FILLER_56_680 ();
 sg13g2_fill_2 FILLER_56_704 ();
 sg13g2_decap_8 FILLER_56_732 ();
 sg13g2_decap_4 FILLER_56_739 ();
 sg13g2_fill_1 FILLER_56_743 ();
 sg13g2_fill_2 FILLER_56_754 ();
 sg13g2_decap_8 FILLER_56_760 ();
 sg13g2_decap_8 FILLER_56_767 ();
 sg13g2_fill_2 FILLER_56_791 ();
 sg13g2_decap_8 FILLER_56_828 ();
 sg13g2_decap_8 FILLER_56_835 ();
 sg13g2_decap_8 FILLER_56_842 ();
 sg13g2_decap_8 FILLER_56_849 ();
 sg13g2_decap_4 FILLER_56_856 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_decap_4 FILLER_57_43 ();
 sg13g2_fill_1 FILLER_57_66 ();
 sg13g2_decap_8 FILLER_57_75 ();
 sg13g2_decap_4 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_1 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_127 ();
 sg13g2_fill_1 FILLER_57_134 ();
 sg13g2_fill_2 FILLER_57_147 ();
 sg13g2_fill_1 FILLER_57_149 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_204 ();
 sg13g2_fill_2 FILLER_57_211 ();
 sg13g2_fill_1 FILLER_57_213 ();
 sg13g2_decap_4 FILLER_57_233 ();
 sg13g2_fill_1 FILLER_57_251 ();
 sg13g2_decap_4 FILLER_57_264 ();
 sg13g2_fill_1 FILLER_57_268 ();
 sg13g2_fill_1 FILLER_57_284 ();
 sg13g2_decap_8 FILLER_57_305 ();
 sg13g2_decap_8 FILLER_57_312 ();
 sg13g2_fill_1 FILLER_57_319 ();
 sg13g2_decap_4 FILLER_57_333 ();
 sg13g2_fill_2 FILLER_57_355 ();
 sg13g2_fill_1 FILLER_57_357 ();
 sg13g2_fill_2 FILLER_57_376 ();
 sg13g2_decap_4 FILLER_57_418 ();
 sg13g2_decap_8 FILLER_57_440 ();
 sg13g2_decap_8 FILLER_57_447 ();
 sg13g2_decap_4 FILLER_57_454 ();
 sg13g2_fill_2 FILLER_57_471 ();
 sg13g2_fill_1 FILLER_57_473 ();
 sg13g2_decap_4 FILLER_57_493 ();
 sg13g2_decap_8 FILLER_57_549 ();
 sg13g2_decap_4 FILLER_57_556 ();
 sg13g2_fill_2 FILLER_57_560 ();
 sg13g2_fill_2 FILLER_57_566 ();
 sg13g2_decap_4 FILLER_57_580 ();
 sg13g2_fill_1 FILLER_57_584 ();
 sg13g2_decap_4 FILLER_57_590 ();
 sg13g2_fill_2 FILLER_57_594 ();
 sg13g2_decap_8 FILLER_57_605 ();
 sg13g2_fill_1 FILLER_57_612 ();
 sg13g2_fill_1 FILLER_57_625 ();
 sg13g2_decap_4 FILLER_57_629 ();
 sg13g2_fill_2 FILLER_57_633 ();
 sg13g2_decap_4 FILLER_57_639 ();
 sg13g2_fill_2 FILLER_57_662 ();
 sg13g2_decap_4 FILLER_57_690 ();
 sg13g2_fill_1 FILLER_57_694 ();
 sg13g2_decap_8 FILLER_57_703 ();
 sg13g2_decap_8 FILLER_57_710 ();
 sg13g2_fill_1 FILLER_57_717 ();
 sg13g2_decap_4 FILLER_57_744 ();
 sg13g2_fill_1 FILLER_57_799 ();
 sg13g2_decap_8 FILLER_57_822 ();
 sg13g2_decap_8 FILLER_57_829 ();
 sg13g2_decap_8 FILLER_57_836 ();
 sg13g2_decap_8 FILLER_57_843 ();
 sg13g2_decap_8 FILLER_57_850 ();
 sg13g2_decap_4 FILLER_57_857 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_19 ();
 sg13g2_fill_2 FILLER_58_26 ();
 sg13g2_fill_1 FILLER_58_41 ();
 sg13g2_decap_8 FILLER_58_50 ();
 sg13g2_decap_8 FILLER_58_57 ();
 sg13g2_fill_2 FILLER_58_64 ();
 sg13g2_decap_4 FILLER_58_78 ();
 sg13g2_fill_1 FILLER_58_82 ();
 sg13g2_fill_2 FILLER_58_87 ();
 sg13g2_decap_8 FILLER_58_97 ();
 sg13g2_decap_4 FILLER_58_104 ();
 sg13g2_decap_8 FILLER_58_113 ();
 sg13g2_fill_2 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_141 ();
 sg13g2_fill_1 FILLER_58_143 ();
 sg13g2_decap_8 FILLER_58_174 ();
 sg13g2_decap_8 FILLER_58_181 ();
 sg13g2_fill_2 FILLER_58_188 ();
 sg13g2_fill_1 FILLER_58_190 ();
 sg13g2_decap_8 FILLER_58_194 ();
 sg13g2_fill_1 FILLER_58_201 ();
 sg13g2_fill_1 FILLER_58_210 ();
 sg13g2_decap_4 FILLER_58_231 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_decap_4 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_276 ();
 sg13g2_decap_8 FILLER_58_282 ();
 sg13g2_decap_4 FILLER_58_289 ();
 sg13g2_fill_1 FILLER_58_293 ();
 sg13g2_decap_4 FILLER_58_298 ();
 sg13g2_fill_2 FILLER_58_302 ();
 sg13g2_fill_2 FILLER_58_317 ();
 sg13g2_decap_8 FILLER_58_335 ();
 sg13g2_decap_8 FILLER_58_342 ();
 sg13g2_fill_2 FILLER_58_349 ();
 sg13g2_fill_1 FILLER_58_351 ();
 sg13g2_decap_4 FILLER_58_368 ();
 sg13g2_fill_2 FILLER_58_372 ();
 sg13g2_fill_2 FILLER_58_391 ();
 sg13g2_fill_1 FILLER_58_397 ();
 sg13g2_decap_8 FILLER_58_403 ();
 sg13g2_fill_1 FILLER_58_422 ();
 sg13g2_decap_4 FILLER_58_475 ();
 sg13g2_fill_2 FILLER_58_500 ();
 sg13g2_decap_8 FILLER_58_507 ();
 sg13g2_decap_4 FILLER_58_514 ();
 sg13g2_fill_1 FILLER_58_531 ();
 sg13g2_fill_1 FILLER_58_545 ();
 sg13g2_fill_2 FILLER_58_600 ();
 sg13g2_decap_8 FILLER_58_628 ();
 sg13g2_fill_1 FILLER_58_655 ();
 sg13g2_fill_2 FILLER_58_668 ();
 sg13g2_fill_2 FILLER_58_683 ();
 sg13g2_decap_4 FILLER_58_711 ();
 sg13g2_fill_2 FILLER_58_715 ();
 sg13g2_fill_2 FILLER_58_726 ();
 sg13g2_fill_2 FILLER_58_732 ();
 sg13g2_decap_8 FILLER_58_763 ();
 sg13g2_decap_4 FILLER_58_770 ();
 sg13g2_fill_2 FILLER_58_774 ();
 sg13g2_decap_8 FILLER_58_824 ();
 sg13g2_decap_8 FILLER_58_831 ();
 sg13g2_decap_8 FILLER_58_838 ();
 sg13g2_decap_8 FILLER_58_845 ();
 sg13g2_decap_8 FILLER_58_852 ();
 sg13g2_fill_2 FILLER_58_859 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_25 ();
 sg13g2_fill_2 FILLER_59_37 ();
 sg13g2_fill_1 FILLER_59_49 ();
 sg13g2_fill_2 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_106 ();
 sg13g2_fill_2 FILLER_59_112 ();
 sg13g2_fill_1 FILLER_59_114 ();
 sg13g2_decap_8 FILLER_59_139 ();
 sg13g2_fill_2 FILLER_59_146 ();
 sg13g2_fill_2 FILLER_59_153 ();
 sg13g2_decap_8 FILLER_59_159 ();
 sg13g2_decap_8 FILLER_59_205 ();
 sg13g2_decap_8 FILLER_59_212 ();
 sg13g2_decap_4 FILLER_59_219 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_decap_8 FILLER_59_234 ();
 sg13g2_decap_4 FILLER_59_241 ();
 sg13g2_fill_1 FILLER_59_245 ();
 sg13g2_fill_2 FILLER_59_250 ();
 sg13g2_decap_8 FILLER_59_265 ();
 sg13g2_decap_4 FILLER_59_272 ();
 sg13g2_fill_1 FILLER_59_276 ();
 sg13g2_fill_1 FILLER_59_282 ();
 sg13g2_fill_2 FILLER_59_295 ();
 sg13g2_decap_8 FILLER_59_305 ();
 sg13g2_decap_8 FILLER_59_312 ();
 sg13g2_decap_8 FILLER_59_345 ();
 sg13g2_fill_2 FILLER_59_352 ();
 sg13g2_fill_1 FILLER_59_354 ();
 sg13g2_fill_2 FILLER_59_359 ();
 sg13g2_fill_1 FILLER_59_361 ();
 sg13g2_decap_4 FILLER_59_368 ();
 sg13g2_fill_2 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_410 ();
 sg13g2_fill_2 FILLER_59_421 ();
 sg13g2_fill_2 FILLER_59_432 ();
 sg13g2_fill_2 FILLER_59_448 ();
 sg13g2_fill_1 FILLER_59_450 ();
 sg13g2_fill_1 FILLER_59_499 ();
 sg13g2_decap_8 FILLER_59_508 ();
 sg13g2_fill_2 FILLER_59_515 ();
 sg13g2_fill_1 FILLER_59_517 ();
 sg13g2_fill_2 FILLER_59_529 ();
 sg13g2_decap_8 FILLER_59_544 ();
 sg13g2_decap_8 FILLER_59_551 ();
 sg13g2_decap_8 FILLER_59_558 ();
 sg13g2_decap_8 FILLER_59_569 ();
 sg13g2_decap_8 FILLER_59_576 ();
 sg13g2_fill_2 FILLER_59_602 ();
 sg13g2_decap_8 FILLER_59_608 ();
 sg13g2_decap_4 FILLER_59_615 ();
 sg13g2_fill_1 FILLER_59_619 ();
 sg13g2_decap_4 FILLER_59_632 ();
 sg13g2_decap_8 FILLER_59_645 ();
 sg13g2_decap_8 FILLER_59_673 ();
 sg13g2_decap_8 FILLER_59_680 ();
 sg13g2_fill_1 FILLER_59_687 ();
 sg13g2_decap_4 FILLER_59_701 ();
 sg13g2_fill_1 FILLER_59_705 ();
 sg13g2_decap_8 FILLER_59_723 ();
 sg13g2_fill_2 FILLER_59_730 ();
 sg13g2_decap_4 FILLER_59_741 ();
 sg13g2_fill_1 FILLER_59_745 ();
 sg13g2_decap_8 FILLER_59_755 ();
 sg13g2_decap_8 FILLER_59_762 ();
 sg13g2_decap_8 FILLER_59_799 ();
 sg13g2_fill_2 FILLER_59_806 ();
 sg13g2_fill_1 FILLER_59_808 ();
 sg13g2_decap_8 FILLER_59_813 ();
 sg13g2_decap_8 FILLER_59_820 ();
 sg13g2_decap_8 FILLER_59_827 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_decap_8 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_fill_1 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_50 ();
 sg13g2_decap_4 FILLER_60_57 ();
 sg13g2_fill_2 FILLER_60_61 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_109 ();
 sg13g2_decap_8 FILLER_60_116 ();
 sg13g2_decap_8 FILLER_60_123 ();
 sg13g2_decap_8 FILLER_60_130 ();
 sg13g2_decap_8 FILLER_60_137 ();
 sg13g2_decap_4 FILLER_60_144 ();
 sg13g2_decap_4 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_165 ();
 sg13g2_decap_8 FILLER_60_176 ();
 sg13g2_decap_8 FILLER_60_183 ();
 sg13g2_decap_8 FILLER_60_190 ();
 sg13g2_decap_8 FILLER_60_197 ();
 sg13g2_fill_1 FILLER_60_204 ();
 sg13g2_fill_1 FILLER_60_217 ();
 sg13g2_decap_4 FILLER_60_245 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_259 ();
 sg13g2_fill_1 FILLER_60_261 ();
 sg13g2_fill_1 FILLER_60_265 ();
 sg13g2_fill_2 FILLER_60_286 ();
 sg13g2_fill_2 FILLER_60_301 ();
 sg13g2_fill_1 FILLER_60_303 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_2 FILLER_60_352 ();
 sg13g2_decap_8 FILLER_60_374 ();
 sg13g2_fill_1 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_407 ();
 sg13g2_decap_4 FILLER_60_414 ();
 sg13g2_decap_4 FILLER_60_422 ();
 sg13g2_decap_8 FILLER_60_452 ();
 sg13g2_decap_8 FILLER_60_459 ();
 sg13g2_fill_1 FILLER_60_466 ();
 sg13g2_fill_2 FILLER_60_481 ();
 sg13g2_fill_1 FILLER_60_483 ();
 sg13g2_decap_8 FILLER_60_506 ();
 sg13g2_fill_2 FILLER_60_513 ();
 sg13g2_fill_1 FILLER_60_515 ();
 sg13g2_decap_4 FILLER_60_537 ();
 sg13g2_fill_1 FILLER_60_541 ();
 sg13g2_fill_2 FILLER_60_554 ();
 sg13g2_fill_1 FILLER_60_556 ();
 sg13g2_fill_2 FILLER_60_562 ();
 sg13g2_fill_1 FILLER_60_564 ();
 sg13g2_fill_2 FILLER_60_578 ();
 sg13g2_decap_8 FILLER_60_588 ();
 sg13g2_decap_4 FILLER_60_595 ();
 sg13g2_fill_1 FILLER_60_599 ();
 sg13g2_decap_8 FILLER_60_610 ();
 sg13g2_decap_4 FILLER_60_617 ();
 sg13g2_fill_2 FILLER_60_621 ();
 sg13g2_decap_4 FILLER_60_633 ();
 sg13g2_fill_2 FILLER_60_637 ();
 sg13g2_decap_8 FILLER_60_651 ();
 sg13g2_decap_4 FILLER_60_676 ();
 sg13g2_fill_2 FILLER_60_688 ();
 sg13g2_decap_8 FILLER_60_703 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_decap_8 FILLER_60_758 ();
 sg13g2_fill_2 FILLER_60_765 ();
 sg13g2_decap_8 FILLER_60_821 ();
 sg13g2_decap_8 FILLER_60_828 ();
 sg13g2_decap_8 FILLER_60_835 ();
 sg13g2_decap_8 FILLER_60_842 ();
 sg13g2_decap_8 FILLER_60_849 ();
 sg13g2_decap_4 FILLER_60_856 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_fill_1 FILLER_61_20 ();
 sg13g2_fill_2 FILLER_61_29 ();
 sg13g2_fill_1 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_38 ();
 sg13g2_decap_8 FILLER_61_44 ();
 sg13g2_decap_8 FILLER_61_51 ();
 sg13g2_fill_1 FILLER_61_58 ();
 sg13g2_decap_4 FILLER_61_70 ();
 sg13g2_fill_2 FILLER_61_74 ();
 sg13g2_fill_1 FILLER_61_84 ();
 sg13g2_fill_1 FILLER_61_95 ();
 sg13g2_fill_1 FILLER_61_115 ();
 sg13g2_fill_2 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_fill_2 FILLER_61_133 ();
 sg13g2_fill_2 FILLER_61_157 ();
 sg13g2_fill_2 FILLER_61_172 ();
 sg13g2_decap_8 FILLER_61_179 ();
 sg13g2_decap_4 FILLER_61_186 ();
 sg13g2_decap_4 FILLER_61_195 ();
 sg13g2_fill_1 FILLER_61_199 ();
 sg13g2_fill_2 FILLER_61_208 ();
 sg13g2_decap_8 FILLER_61_242 ();
 sg13g2_decap_8 FILLER_61_249 ();
 sg13g2_decap_8 FILLER_61_270 ();
 sg13g2_fill_2 FILLER_61_277 ();
 sg13g2_decap_4 FILLER_61_295 ();
 sg13g2_fill_2 FILLER_61_299 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_331 ();
 sg13g2_fill_1 FILLER_61_338 ();
 sg13g2_decap_8 FILLER_61_345 ();
 sg13g2_decap_4 FILLER_61_352 ();
 sg13g2_decap_8 FILLER_61_376 ();
 sg13g2_decap_4 FILLER_61_383 ();
 sg13g2_fill_2 FILLER_61_387 ();
 sg13g2_decap_8 FILLER_61_397 ();
 sg13g2_decap_8 FILLER_61_404 ();
 sg13g2_fill_2 FILLER_61_411 ();
 sg13g2_fill_1 FILLER_61_413 ();
 sg13g2_decap_8 FILLER_61_427 ();
 sg13g2_fill_1 FILLER_61_434 ();
 sg13g2_decap_4 FILLER_61_440 ();
 sg13g2_decap_8 FILLER_61_450 ();
 sg13g2_fill_1 FILLER_61_457 ();
 sg13g2_decap_4 FILLER_61_471 ();
 sg13g2_fill_2 FILLER_61_475 ();
 sg13g2_decap_8 FILLER_61_481 ();
 sg13g2_decap_4 FILLER_61_506 ();
 sg13g2_decap_8 FILLER_61_518 ();
 sg13g2_decap_4 FILLER_61_525 ();
 sg13g2_fill_1 FILLER_61_529 ();
 sg13g2_decap_8 FILLER_61_542 ();
 sg13g2_fill_2 FILLER_61_574 ();
 sg13g2_fill_1 FILLER_61_576 ();
 sg13g2_decap_4 FILLER_61_590 ();
 sg13g2_decap_8 FILLER_61_610 ();
 sg13g2_fill_2 FILLER_61_617 ();
 sg13g2_fill_1 FILLER_61_619 ();
 sg13g2_decap_4 FILLER_61_633 ();
 sg13g2_fill_2 FILLER_61_650 ();
 sg13g2_fill_1 FILLER_61_652 ();
 sg13g2_decap_8 FILLER_61_682 ();
 sg13g2_decap_8 FILLER_61_689 ();
 sg13g2_decap_8 FILLER_61_696 ();
 sg13g2_fill_2 FILLER_61_703 ();
 sg13g2_fill_1 FILLER_61_719 ();
 sg13g2_decap_8 FILLER_61_740 ();
 sg13g2_decap_8 FILLER_61_752 ();
 sg13g2_decap_4 FILLER_61_759 ();
 sg13g2_fill_1 FILLER_61_767 ();
 sg13g2_fill_2 FILLER_61_787 ();
 sg13g2_decap_4 FILLER_61_802 ();
 sg13g2_decap_8 FILLER_61_810 ();
 sg13g2_decap_8 FILLER_61_817 ();
 sg13g2_decap_8 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_decap_8 FILLER_61_838 ();
 sg13g2_decap_8 FILLER_61_845 ();
 sg13g2_decap_8 FILLER_61_852 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_17 ();
 sg13g2_fill_1 FILLER_62_32 ();
 sg13g2_fill_2 FILLER_62_47 ();
 sg13g2_decap_4 FILLER_62_71 ();
 sg13g2_fill_2 FILLER_62_75 ();
 sg13g2_decap_8 FILLER_62_83 ();
 sg13g2_decap_4 FILLER_62_90 ();
 sg13g2_decap_8 FILLER_62_109 ();
 sg13g2_decap_4 FILLER_62_116 ();
 sg13g2_fill_2 FILLER_62_120 ();
 sg13g2_fill_1 FILLER_62_142 ();
 sg13g2_decap_4 FILLER_62_147 ();
 sg13g2_decap_4 FILLER_62_165 ();
 sg13g2_decap_4 FILLER_62_195 ();
 sg13g2_decap_8 FILLER_62_221 ();
 sg13g2_decap_8 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_decap_8 FILLER_62_240 ();
 sg13g2_decap_4 FILLER_62_247 ();
 sg13g2_fill_2 FILLER_62_251 ();
 sg13g2_fill_1 FILLER_62_275 ();
 sg13g2_fill_1 FILLER_62_284 ();
 sg13g2_decap_8 FILLER_62_293 ();
 sg13g2_decap_4 FILLER_62_300 ();
 sg13g2_fill_2 FILLER_62_304 ();
 sg13g2_fill_2 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_62_379 ();
 sg13g2_fill_1 FILLER_62_381 ();
 sg13g2_decap_4 FILLER_62_433 ();
 sg13g2_fill_1 FILLER_62_437 ();
 sg13g2_decap_4 FILLER_62_450 ();
 sg13g2_fill_2 FILLER_62_454 ();
 sg13g2_decap_8 FILLER_62_469 ();
 sg13g2_decap_8 FILLER_62_476 ();
 sg13g2_fill_1 FILLER_62_483 ();
 sg13g2_decap_8 FILLER_62_493 ();
 sg13g2_decap_8 FILLER_62_500 ();
 sg13g2_decap_8 FILLER_62_507 ();
 sg13g2_fill_2 FILLER_62_514 ();
 sg13g2_decap_8 FILLER_62_553 ();
 sg13g2_decap_8 FILLER_62_560 ();
 sg13g2_fill_1 FILLER_62_567 ();
 sg13g2_fill_2 FILLER_62_584 ();
 sg13g2_decap_4 FILLER_62_598 ();
 sg13g2_fill_1 FILLER_62_602 ();
 sg13g2_fill_2 FILLER_62_608 ();
 sg13g2_decap_4 FILLER_62_622 ();
 sg13g2_fill_1 FILLER_62_626 ();
 sg13g2_fill_2 FILLER_62_639 ();
 sg13g2_decap_8 FILLER_62_654 ();
 sg13g2_fill_2 FILLER_62_661 ();
 sg13g2_fill_1 FILLER_62_676 ();
 sg13g2_fill_1 FILLER_62_703 ();
 sg13g2_fill_2 FILLER_62_725 ();
 sg13g2_decap_8 FILLER_62_751 ();
 sg13g2_fill_2 FILLER_62_758 ();
 sg13g2_fill_1 FILLER_62_760 ();
 sg13g2_decap_4 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_814 ();
 sg13g2_decap_8 FILLER_62_821 ();
 sg13g2_decap_8 FILLER_62_828 ();
 sg13g2_decap_8 FILLER_62_835 ();
 sg13g2_decap_8 FILLER_62_842 ();
 sg13g2_decap_8 FILLER_62_849 ();
 sg13g2_decap_4 FILLER_62_856 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_decap_4 FILLER_63_40 ();
 sg13g2_fill_2 FILLER_63_44 ();
 sg13g2_fill_2 FILLER_63_58 ();
 sg13g2_decap_4 FILLER_63_67 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_decap_8 FILLER_63_76 ();
 sg13g2_fill_1 FILLER_63_83 ();
 sg13g2_decap_4 FILLER_63_107 ();
 sg13g2_fill_2 FILLER_63_111 ();
 sg13g2_decap_8 FILLER_63_118 ();
 sg13g2_fill_2 FILLER_63_125 ();
 sg13g2_decap_4 FILLER_63_132 ();
 sg13g2_decap_4 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_149 ();
 sg13g2_decap_8 FILLER_63_159 ();
 sg13g2_decap_4 FILLER_63_166 ();
 sg13g2_fill_1 FILLER_63_170 ();
 sg13g2_fill_1 FILLER_63_179 ();
 sg13g2_decap_8 FILLER_63_185 ();
 sg13g2_fill_2 FILLER_63_192 ();
 sg13g2_fill_1 FILLER_63_194 ();
 sg13g2_decap_8 FILLER_63_207 ();
 sg13g2_decap_8 FILLER_63_214 ();
 sg13g2_decap_4 FILLER_63_221 ();
 sg13g2_decap_8 FILLER_63_246 ();
 sg13g2_decap_4 FILLER_63_258 ();
 sg13g2_decap_8 FILLER_63_270 ();
 sg13g2_fill_2 FILLER_63_277 ();
 sg13g2_fill_1 FILLER_63_279 ();
 sg13g2_decap_8 FILLER_63_285 ();
 sg13g2_decap_8 FILLER_63_292 ();
 sg13g2_decap_8 FILLER_63_299 ();
 sg13g2_fill_2 FILLER_63_311 ();
 sg13g2_fill_2 FILLER_63_322 ();
 sg13g2_fill_2 FILLER_63_346 ();
 sg13g2_fill_1 FILLER_63_348 ();
 sg13g2_fill_2 FILLER_63_374 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_decap_4 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_386 ();
 sg13g2_decap_8 FILLER_63_401 ();
 sg13g2_decap_8 FILLER_63_408 ();
 sg13g2_fill_2 FILLER_63_415 ();
 sg13g2_decap_4 FILLER_63_426 ();
 sg13g2_fill_1 FILLER_63_430 ();
 sg13g2_decap_8 FILLER_63_447 ();
 sg13g2_fill_1 FILLER_63_478 ();
 sg13g2_fill_2 FILLER_63_525 ();
 sg13g2_fill_1 FILLER_63_527 ();
 sg13g2_decap_8 FILLER_63_544 ();
 sg13g2_fill_2 FILLER_63_551 ();
 sg13g2_fill_1 FILLER_63_553 ();
 sg13g2_fill_2 FILLER_63_559 ();
 sg13g2_decap_8 FILLER_63_582 ();
 sg13g2_decap_4 FILLER_63_589 ();
 sg13g2_fill_1 FILLER_63_593 ();
 sg13g2_decap_4 FILLER_63_615 ();
 sg13g2_decap_8 FILLER_63_637 ();
 sg13g2_decap_8 FILLER_63_644 ();
 sg13g2_decap_8 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_658 ();
 sg13g2_decap_8 FILLER_63_665 ();
 sg13g2_decap_4 FILLER_63_672 ();
 sg13g2_fill_2 FILLER_63_685 ();
 sg13g2_fill_1 FILLER_63_687 ();
 sg13g2_decap_8 FILLER_63_692 ();
 sg13g2_decap_8 FILLER_63_699 ();
 sg13g2_fill_2 FILLER_63_706 ();
 sg13g2_fill_1 FILLER_63_708 ();
 sg13g2_decap_8 FILLER_63_758 ();
 sg13g2_fill_1 FILLER_63_776 ();
 sg13g2_fill_2 FILLER_63_791 ();
 sg13g2_fill_2 FILLER_63_796 ();
 sg13g2_fill_1 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_803 ();
 sg13g2_decap_8 FILLER_63_810 ();
 sg13g2_decap_8 FILLER_63_817 ();
 sg13g2_decap_8 FILLER_63_824 ();
 sg13g2_decap_8 FILLER_63_831 ();
 sg13g2_decap_8 FILLER_63_838 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_16 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_fill_1 FILLER_64_28 ();
 sg13g2_fill_2 FILLER_64_38 ();
 sg13g2_fill_1 FILLER_64_40 ();
 sg13g2_decap_4 FILLER_64_49 ();
 sg13g2_fill_1 FILLER_64_53 ();
 sg13g2_fill_2 FILLER_64_62 ();
 sg13g2_fill_1 FILLER_64_70 ();
 sg13g2_decap_4 FILLER_64_87 ();
 sg13g2_fill_2 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_125 ();
 sg13g2_decap_4 FILLER_64_132 ();
 sg13g2_fill_1 FILLER_64_141 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_4 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_172 ();
 sg13g2_decap_4 FILLER_64_194 ();
 sg13g2_fill_1 FILLER_64_198 ();
 sg13g2_decap_4 FILLER_64_215 ();
 sg13g2_fill_2 FILLER_64_219 ();
 sg13g2_decap_8 FILLER_64_249 ();
 sg13g2_decap_8 FILLER_64_256 ();
 sg13g2_fill_2 FILLER_64_263 ();
 sg13g2_fill_2 FILLER_64_271 ();
 sg13g2_decap_8 FILLER_64_302 ();
 sg13g2_decap_4 FILLER_64_309 ();
 sg13g2_fill_1 FILLER_64_313 ();
 sg13g2_decap_8 FILLER_64_372 ();
 sg13g2_fill_2 FILLER_64_379 ();
 sg13g2_fill_1 FILLER_64_381 ();
 sg13g2_fill_1 FILLER_64_390 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_8 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_410 ();
 sg13g2_fill_1 FILLER_64_412 ();
 sg13g2_fill_1 FILLER_64_421 ();
 sg13g2_decap_8 FILLER_64_438 ();
 sg13g2_decap_8 FILLER_64_445 ();
 sg13g2_decap_8 FILLER_64_452 ();
 sg13g2_fill_1 FILLER_64_459 ();
 sg13g2_decap_8 FILLER_64_468 ();
 sg13g2_decap_8 FILLER_64_475 ();
 sg13g2_decap_8 FILLER_64_482 ();
 sg13g2_fill_2 FILLER_64_493 ();
 sg13g2_fill_1 FILLER_64_495 ();
 sg13g2_decap_8 FILLER_64_501 ();
 sg13g2_fill_2 FILLER_64_508 ();
 sg13g2_decap_4 FILLER_64_518 ();
 sg13g2_fill_1 FILLER_64_522 ();
 sg13g2_fill_2 FILLER_64_528 ();
 sg13g2_decap_8 FILLER_64_535 ();
 sg13g2_decap_8 FILLER_64_542 ();
 sg13g2_fill_2 FILLER_64_549 ();
 sg13g2_decap_4 FILLER_64_569 ();
 sg13g2_fill_2 FILLER_64_573 ();
 sg13g2_decap_8 FILLER_64_584 ();
 sg13g2_decap_4 FILLER_64_591 ();
 sg13g2_decap_8 FILLER_64_608 ();
 sg13g2_decap_8 FILLER_64_615 ();
 sg13g2_fill_2 FILLER_64_622 ();
 sg13g2_decap_8 FILLER_64_640 ();
 sg13g2_fill_1 FILLER_64_647 ();
 sg13g2_decap_4 FILLER_64_673 ();
 sg13g2_fill_2 FILLER_64_677 ();
 sg13g2_decap_4 FILLER_64_684 ();
 sg13g2_fill_1 FILLER_64_691 ();
 sg13g2_fill_2 FILLER_64_716 ();
 sg13g2_decap_8 FILLER_64_727 ();
 sg13g2_decap_4 FILLER_64_734 ();
 sg13g2_fill_1 FILLER_64_738 ();
 sg13g2_decap_8 FILLER_64_746 ();
 sg13g2_decap_4 FILLER_64_753 ();
 sg13g2_decap_4 FILLER_64_768 ();
 sg13g2_fill_1 FILLER_64_772 ();
 sg13g2_decap_8 FILLER_64_814 ();
 sg13g2_decap_8 FILLER_64_821 ();
 sg13g2_decap_8 FILLER_64_828 ();
 sg13g2_decap_8 FILLER_64_835 ();
 sg13g2_decap_8 FILLER_64_842 ();
 sg13g2_decap_8 FILLER_64_849 ();
 sg13g2_decap_4 FILLER_64_856 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_fill_2 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_63 ();
 sg13g2_fill_1 FILLER_65_65 ();
 sg13g2_decap_8 FILLER_65_75 ();
 sg13g2_decap_8 FILLER_65_82 ();
 sg13g2_decap_4 FILLER_65_89 ();
 sg13g2_fill_1 FILLER_65_93 ();
 sg13g2_fill_1 FILLER_65_110 ();
 sg13g2_fill_2 FILLER_65_115 ();
 sg13g2_decap_4 FILLER_65_122 ();
 sg13g2_fill_2 FILLER_65_131 ();
 sg13g2_fill_1 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_142 ();
 sg13g2_fill_2 FILLER_65_149 ();
 sg13g2_fill_2 FILLER_65_159 ();
 sg13g2_decap_8 FILLER_65_169 ();
 sg13g2_fill_1 FILLER_65_176 ();
 sg13g2_decap_4 FILLER_65_190 ();
 sg13g2_decap_8 FILLER_65_211 ();
 sg13g2_decap_8 FILLER_65_218 ();
 sg13g2_decap_4 FILLER_65_225 ();
 sg13g2_fill_2 FILLER_65_239 ();
 sg13g2_fill_1 FILLER_65_241 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_fill_2 FILLER_65_252 ();
 sg13g2_decap_4 FILLER_65_270 ();
 sg13g2_fill_2 FILLER_65_274 ();
 sg13g2_decap_4 FILLER_65_299 ();
 sg13g2_fill_2 FILLER_65_303 ();
 sg13g2_decap_4 FILLER_65_315 ();
 sg13g2_fill_1 FILLER_65_319 ();
 sg13g2_fill_2 FILLER_65_338 ();
 sg13g2_fill_1 FILLER_65_340 ();
 sg13g2_decap_4 FILLER_65_354 ();
 sg13g2_fill_2 FILLER_65_358 ();
 sg13g2_fill_2 FILLER_65_370 ();
 sg13g2_decap_4 FILLER_65_377 ();
 sg13g2_fill_1 FILLER_65_381 ();
 sg13g2_decap_4 FILLER_65_387 ();
 sg13g2_fill_2 FILLER_65_401 ();
 sg13g2_decap_4 FILLER_65_418 ();
 sg13g2_fill_2 FILLER_65_422 ();
 sg13g2_fill_2 FILLER_65_441 ();
 sg13g2_fill_2 FILLER_65_458 ();
 sg13g2_fill_1 FILLER_65_460 ();
 sg13g2_fill_2 FILLER_65_478 ();
 sg13g2_fill_2 FILLER_65_499 ();
 sg13g2_decap_4 FILLER_65_508 ();
 sg13g2_fill_1 FILLER_65_512 ();
 sg13g2_decap_8 FILLER_65_518 ();
 sg13g2_decap_8 FILLER_65_525 ();
 sg13g2_decap_8 FILLER_65_532 ();
 sg13g2_decap_8 FILLER_65_539 ();
 sg13g2_fill_2 FILLER_65_554 ();
 sg13g2_fill_1 FILLER_65_556 ();
 sg13g2_decap_8 FILLER_65_560 ();
 sg13g2_fill_2 FILLER_65_567 ();
 sg13g2_decap_4 FILLER_65_593 ();
 sg13g2_fill_2 FILLER_65_600 ();
 sg13g2_fill_1 FILLER_65_610 ();
 sg13g2_fill_2 FILLER_65_619 ();
 sg13g2_fill_1 FILLER_65_621 ();
 sg13g2_fill_1 FILLER_65_636 ();
 sg13g2_decap_8 FILLER_65_673 ();
 sg13g2_fill_1 FILLER_65_680 ();
 sg13g2_decap_8 FILLER_65_726 ();
 sg13g2_decap_8 FILLER_65_733 ();
 sg13g2_fill_2 FILLER_65_740 ();
 sg13g2_fill_2 FILLER_65_777 ();
 sg13g2_fill_1 FILLER_65_779 ();
 sg13g2_fill_1 FILLER_65_789 ();
 sg13g2_fill_2 FILLER_65_798 ();
 sg13g2_fill_1 FILLER_65_800 ();
 sg13g2_decap_8 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_817 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_831 ();
 sg13g2_decap_8 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_845 ();
 sg13g2_decap_8 FILLER_65_852 ();
 sg13g2_fill_2 FILLER_65_859 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_fill_1 FILLER_66_55 ();
 sg13g2_fill_2 FILLER_66_68 ();
 sg13g2_fill_1 FILLER_66_70 ();
 sg13g2_decap_4 FILLER_66_76 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_fill_1 FILLER_66_113 ();
 sg13g2_fill_2 FILLER_66_122 ();
 sg13g2_fill_1 FILLER_66_132 ();
 sg13g2_decap_8 FILLER_66_150 ();
 sg13g2_fill_2 FILLER_66_157 ();
 sg13g2_fill_1 FILLER_66_159 ();
 sg13g2_decap_4 FILLER_66_172 ();
 sg13g2_decap_8 FILLER_66_180 ();
 sg13g2_decap_8 FILLER_66_187 ();
 sg13g2_decap_8 FILLER_66_194 ();
 sg13g2_decap_4 FILLER_66_201 ();
 sg13g2_fill_1 FILLER_66_205 ();
 sg13g2_decap_4 FILLER_66_220 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_250 ();
 sg13g2_decap_8 FILLER_66_265 ();
 sg13g2_decap_8 FILLER_66_272 ();
 sg13g2_decap_8 FILLER_66_298 ();
 sg13g2_decap_8 FILLER_66_305 ();
 sg13g2_decap_8 FILLER_66_312 ();
 sg13g2_fill_2 FILLER_66_319 ();
 sg13g2_fill_1 FILLER_66_321 ();
 sg13g2_fill_1 FILLER_66_365 ();
 sg13g2_decap_8 FILLER_66_374 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_66_414 ();
 sg13g2_decap_8 FILLER_66_421 ();
 sg13g2_fill_1 FILLER_66_428 ();
 sg13g2_decap_8 FILLER_66_438 ();
 sg13g2_decap_4 FILLER_66_445 ();
 sg13g2_fill_2 FILLER_66_449 ();
 sg13g2_fill_1 FILLER_66_459 ();
 sg13g2_fill_2 FILLER_66_464 ();
 sg13g2_fill_1 FILLER_66_466 ();
 sg13g2_fill_2 FILLER_66_470 ();
 sg13g2_decap_8 FILLER_66_498 ();
 sg13g2_fill_1 FILLER_66_531 ();
 sg13g2_decap_8 FILLER_66_583 ();
 sg13g2_decap_4 FILLER_66_590 ();
 sg13g2_decap_8 FILLER_66_602 ();
 sg13g2_decap_8 FILLER_66_609 ();
 sg13g2_fill_2 FILLER_66_616 ();
 sg13g2_decap_8 FILLER_66_638 ();
 sg13g2_fill_2 FILLER_66_645 ();
 sg13g2_fill_2 FILLER_66_656 ();
 sg13g2_decap_8 FILLER_66_683 ();
 sg13g2_fill_1 FILLER_66_690 ();
 sg13g2_decap_8 FILLER_66_697 ();
 sg13g2_fill_2 FILLER_66_704 ();
 sg13g2_fill_1 FILLER_66_706 ();
 sg13g2_fill_2 FILLER_66_758 ();
 sg13g2_fill_1 FILLER_66_760 ();
 sg13g2_decap_8 FILLER_66_770 ();
 sg13g2_fill_2 FILLER_66_777 ();
 sg13g2_fill_1 FILLER_66_779 ();
 sg13g2_fill_1 FILLER_66_792 ();
 sg13g2_decap_8 FILLER_66_827 ();
 sg13g2_decap_8 FILLER_66_834 ();
 sg13g2_decap_8 FILLER_66_841 ();
 sg13g2_decap_8 FILLER_66_848 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_fill_2 FILLER_67_30 ();
 sg13g2_fill_1 FILLER_67_32 ();
 sg13g2_decap_8 FILLER_67_45 ();
 sg13g2_decap_8 FILLER_67_52 ();
 sg13g2_decap_8 FILLER_67_59 ();
 sg13g2_decap_8 FILLER_67_82 ();
 sg13g2_decap_4 FILLER_67_89 ();
 sg13g2_fill_2 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_108 ();
 sg13g2_decap_8 FILLER_67_115 ();
 sg13g2_decap_8 FILLER_67_122 ();
 sg13g2_fill_1 FILLER_67_129 ();
 sg13g2_fill_2 FILLER_67_139 ();
 sg13g2_fill_1 FILLER_67_141 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_fill_2 FILLER_67_159 ();
 sg13g2_decap_4 FILLER_67_169 ();
 sg13g2_fill_2 FILLER_67_191 ();
 sg13g2_decap_8 FILLER_67_209 ();
 sg13g2_decap_8 FILLER_67_216 ();
 sg13g2_fill_2 FILLER_67_223 ();
 sg13g2_fill_1 FILLER_67_231 ();
 sg13g2_fill_2 FILLER_67_236 ();
 sg13g2_decap_8 FILLER_67_242 ();
 sg13g2_fill_2 FILLER_67_249 ();
 sg13g2_decap_8 FILLER_67_257 ();
 sg13g2_decap_8 FILLER_67_264 ();
 sg13g2_fill_2 FILLER_67_271 ();
 sg13g2_fill_2 FILLER_67_301 ();
 sg13g2_decap_4 FILLER_67_317 ();
 sg13g2_fill_1 FILLER_67_321 ();
 sg13g2_fill_2 FILLER_67_335 ();
 sg13g2_fill_1 FILLER_67_337 ();
 sg13g2_decap_8 FILLER_67_346 ();
 sg13g2_decap_8 FILLER_67_353 ();
 sg13g2_fill_2 FILLER_67_360 ();
 sg13g2_decap_8 FILLER_67_375 ();
 sg13g2_fill_2 FILLER_67_422 ();
 sg13g2_decap_4 FILLER_67_442 ();
 sg13g2_decap_8 FILLER_67_464 ();
 sg13g2_fill_2 FILLER_67_471 ();
 sg13g2_decap_8 FILLER_67_499 ();
 sg13g2_fill_2 FILLER_67_523 ();
 sg13g2_fill_2 FILLER_67_530 ();
 sg13g2_fill_2 FILLER_67_541 ();
 sg13g2_decap_8 FILLER_67_552 ();
 sg13g2_decap_4 FILLER_67_559 ();
 sg13g2_fill_2 FILLER_67_563 ();
 sg13g2_decap_4 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_614 ();
 sg13g2_fill_2 FILLER_67_621 ();
 sg13g2_fill_2 FILLER_67_627 ();
 sg13g2_fill_1 FILLER_67_629 ();
 sg13g2_decap_8 FILLER_67_642 ();
 sg13g2_decap_8 FILLER_67_649 ();
 sg13g2_decap_8 FILLER_67_672 ();
 sg13g2_decap_4 FILLER_67_687 ();
 sg13g2_decap_8 FILLER_67_716 ();
 sg13g2_fill_2 FILLER_67_723 ();
 sg13g2_fill_1 FILLER_67_725 ();
 sg13g2_decap_8 FILLER_67_730 ();
 sg13g2_decap_8 FILLER_67_737 ();
 sg13g2_decap_4 FILLER_67_744 ();
 sg13g2_fill_1 FILLER_67_748 ();
 sg13g2_fill_2 FILLER_67_775 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_fill_2 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_33 ();
 sg13g2_fill_2 FILLER_68_52 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_4 FILLER_68_84 ();
 sg13g2_fill_1 FILLER_68_88 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_fill_2 FILLER_68_119 ();
 sg13g2_fill_1 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_138 ();
 sg13g2_decap_8 FILLER_68_145 ();
 sg13g2_decap_4 FILLER_68_152 ();
 sg13g2_fill_1 FILLER_68_160 ();
 sg13g2_decap_4 FILLER_68_170 ();
 sg13g2_fill_1 FILLER_68_174 ();
 sg13g2_fill_2 FILLER_68_189 ();
 sg13g2_fill_2 FILLER_68_219 ();
 sg13g2_decap_4 FILLER_68_237 ();
 sg13g2_decap_4 FILLER_68_273 ();
 sg13g2_fill_1 FILLER_68_277 ();
 sg13g2_fill_2 FILLER_68_281 ();
 sg13g2_fill_1 FILLER_68_283 ();
 sg13g2_decap_8 FILLER_68_292 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_fill_1 FILLER_68_306 ();
 sg13g2_fill_2 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_335 ();
 sg13g2_decap_8 FILLER_68_345 ();
 sg13g2_decap_4 FILLER_68_352 ();
 sg13g2_fill_1 FILLER_68_356 ();
 sg13g2_decap_8 FILLER_68_366 ();
 sg13g2_decap_8 FILLER_68_373 ();
 sg13g2_fill_1 FILLER_68_380 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_fill_2 FILLER_68_409 ();
 sg13g2_decap_8 FILLER_68_416 ();
 sg13g2_decap_8 FILLER_68_423 ();
 sg13g2_fill_1 FILLER_68_430 ();
 sg13g2_decap_8 FILLER_68_436 ();
 sg13g2_decap_4 FILLER_68_443 ();
 sg13g2_fill_2 FILLER_68_447 ();
 sg13g2_decap_8 FILLER_68_465 ();
 sg13g2_decap_8 FILLER_68_472 ();
 sg13g2_decap_4 FILLER_68_479 ();
 sg13g2_fill_1 FILLER_68_483 ();
 sg13g2_decap_4 FILLER_68_488 ();
 sg13g2_fill_2 FILLER_68_492 ();
 sg13g2_fill_2 FILLER_68_537 ();
 sg13g2_fill_1 FILLER_68_554 ();
 sg13g2_fill_2 FILLER_68_559 ();
 sg13g2_fill_1 FILLER_68_561 ();
 sg13g2_fill_1 FILLER_68_566 ();
 sg13g2_fill_2 FILLER_68_577 ();
 sg13g2_fill_2 FILLER_68_609 ();
 sg13g2_decap_4 FILLER_68_619 ();
 sg13g2_decap_4 FILLER_68_631 ();
 sg13g2_fill_2 FILLER_68_656 ();
 sg13g2_fill_2 FILLER_68_666 ();
 sg13g2_fill_1 FILLER_68_668 ();
 sg13g2_decap_8 FILLER_68_678 ();
 sg13g2_fill_2 FILLER_68_685 ();
 sg13g2_fill_2 FILLER_68_719 ();
 sg13g2_decap_8 FILLER_68_747 ();
 sg13g2_decap_4 FILLER_68_754 ();
 sg13g2_fill_1 FILLER_68_758 ();
 sg13g2_decap_4 FILLER_68_772 ();
 sg13g2_decap_8 FILLER_68_819 ();
 sg13g2_decap_8 FILLER_68_826 ();
 sg13g2_decap_8 FILLER_68_833 ();
 sg13g2_decap_8 FILLER_68_840 ();
 sg13g2_decap_8 FILLER_68_847 ();
 sg13g2_decap_8 FILLER_68_854 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_9 ();
 sg13g2_fill_1 FILLER_69_28 ();
 sg13g2_decap_4 FILLER_69_64 ();
 sg13g2_fill_2 FILLER_69_79 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_fill_1 FILLER_69_99 ();
 sg13g2_fill_1 FILLER_69_113 ();
 sg13g2_fill_2 FILLER_69_118 ();
 sg13g2_fill_2 FILLER_69_125 ();
 sg13g2_fill_2 FILLER_69_131 ();
 sg13g2_fill_1 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_156 ();
 sg13g2_fill_2 FILLER_69_177 ();
 sg13g2_fill_1 FILLER_69_179 ();
 sg13g2_decap_4 FILLER_69_192 ();
 sg13g2_fill_2 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_211 ();
 sg13g2_fill_2 FILLER_69_218 ();
 sg13g2_fill_1 FILLER_69_220 ();
 sg13g2_decap_4 FILLER_69_234 ();
 sg13g2_decap_4 FILLER_69_243 ();
 sg13g2_fill_2 FILLER_69_247 ();
 sg13g2_decap_4 FILLER_69_268 ();
 sg13g2_decap_4 FILLER_69_277 ();
 sg13g2_fill_1 FILLER_69_281 ();
 sg13g2_fill_1 FILLER_69_292 ();
 sg13g2_decap_4 FILLER_69_298 ();
 sg13g2_fill_2 FILLER_69_302 ();
 sg13g2_decap_4 FILLER_69_320 ();
 sg13g2_fill_1 FILLER_69_324 ();
 sg13g2_fill_2 FILLER_69_352 ();
 sg13g2_decap_8 FILLER_69_376 ();
 sg13g2_decap_4 FILLER_69_387 ();
 sg13g2_fill_2 FILLER_69_404 ();
 sg13g2_decap_4 FILLER_69_422 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_4 FILLER_69_438 ();
 sg13g2_fill_1 FILLER_69_442 ();
 sg13g2_fill_2 FILLER_69_466 ();
 sg13g2_decap_4 FILLER_69_494 ();
 sg13g2_decap_8 FILLER_69_512 ();
 sg13g2_fill_2 FILLER_69_519 ();
 sg13g2_fill_1 FILLER_69_521 ();
 sg13g2_decap_4 FILLER_69_538 ();
 sg13g2_fill_2 FILLER_69_542 ();
 sg13g2_decap_4 FILLER_69_549 ();
 sg13g2_fill_2 FILLER_69_553 ();
 sg13g2_fill_2 FILLER_69_560 ();
 sg13g2_fill_1 FILLER_69_562 ();
 sg13g2_decap_8 FILLER_69_568 ();
 sg13g2_fill_2 FILLER_69_575 ();
 sg13g2_fill_2 FILLER_69_589 ();
 sg13g2_decap_8 FILLER_69_595 ();
 sg13g2_fill_2 FILLER_69_602 ();
 sg13g2_fill_1 FILLER_69_604 ();
 sg13g2_fill_2 FILLER_69_610 ();
 sg13g2_decap_8 FILLER_69_617 ();
 sg13g2_decap_8 FILLER_69_624 ();
 sg13g2_decap_4 FILLER_69_631 ();
 sg13g2_fill_2 FILLER_69_635 ();
 sg13g2_decap_8 FILLER_69_650 ();
 sg13g2_fill_2 FILLER_69_657 ();
 sg13g2_fill_1 FILLER_69_659 ();
 sg13g2_fill_2 FILLER_69_664 ();
 sg13g2_fill_2 FILLER_69_701 ();
 sg13g2_fill_2 FILLER_69_709 ();
 sg13g2_fill_1 FILLER_69_711 ();
 sg13g2_fill_2 FILLER_69_730 ();
 sg13g2_decap_8 FILLER_69_736 ();
 sg13g2_decap_8 FILLER_69_743 ();
 sg13g2_decap_8 FILLER_69_750 ();
 sg13g2_decap_8 FILLER_69_757 ();
 sg13g2_decap_8 FILLER_69_764 ();
 sg13g2_fill_2 FILLER_69_771 ();
 sg13g2_fill_1 FILLER_69_773 ();
 sg13g2_decap_8 FILLER_69_786 ();
 sg13g2_decap_8 FILLER_69_793 ();
 sg13g2_fill_1 FILLER_69_800 ();
 sg13g2_decap_8 FILLER_69_814 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_decap_8 FILLER_69_842 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_4 FILLER_69_856 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_31 ();
 sg13g2_decap_8 FILLER_70_38 ();
 sg13g2_decap_8 FILLER_70_45 ();
 sg13g2_fill_2 FILLER_70_52 ();
 sg13g2_fill_1 FILLER_70_54 ();
 sg13g2_fill_2 FILLER_70_60 ();
 sg13g2_decap_8 FILLER_70_68 ();
 sg13g2_decap_8 FILLER_70_75 ();
 sg13g2_decap_8 FILLER_70_82 ();
 sg13g2_decap_8 FILLER_70_89 ();
 sg13g2_decap_4 FILLER_70_96 ();
 sg13g2_fill_2 FILLER_70_100 ();
 sg13g2_decap_8 FILLER_70_106 ();
 sg13g2_decap_8 FILLER_70_113 ();
 sg13g2_decap_8 FILLER_70_120 ();
 sg13g2_decap_4 FILLER_70_127 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_1 FILLER_70_151 ();
 sg13g2_decap_8 FILLER_70_158 ();
 sg13g2_decap_8 FILLER_70_165 ();
 sg13g2_decap_4 FILLER_70_172 ();
 sg13g2_fill_1 FILLER_70_176 ();
 sg13g2_fill_2 FILLER_70_182 ();
 sg13g2_fill_1 FILLER_70_184 ();
 sg13g2_fill_2 FILLER_70_192 ();
 sg13g2_fill_2 FILLER_70_208 ();
 sg13g2_fill_2 FILLER_70_218 ();
 sg13g2_fill_1 FILLER_70_220 ();
 sg13g2_fill_2 FILLER_70_226 ();
 sg13g2_fill_1 FILLER_70_228 ();
 sg13g2_fill_1 FILLER_70_235 ();
 sg13g2_decap_8 FILLER_70_249 ();
 sg13g2_fill_1 FILLER_70_256 ();
 sg13g2_decap_8 FILLER_70_262 ();
 sg13g2_decap_8 FILLER_70_281 ();
 sg13g2_decap_8 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_295 ();
 sg13g2_decap_8 FILLER_70_321 ();
 sg13g2_fill_2 FILLER_70_328 ();
 sg13g2_fill_1 FILLER_70_330 ();
 sg13g2_fill_2 FILLER_70_341 ();
 sg13g2_decap_4 FILLER_70_350 ();
 sg13g2_fill_2 FILLER_70_354 ();
 sg13g2_fill_1 FILLER_70_361 ();
 sg13g2_fill_2 FILLER_70_365 ();
 sg13g2_fill_1 FILLER_70_367 ();
 sg13g2_decap_4 FILLER_70_393 ();
 sg13g2_decap_4 FILLER_70_402 ();
 sg13g2_fill_2 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_437 ();
 sg13g2_decap_8 FILLER_70_444 ();
 sg13g2_decap_8 FILLER_70_466 ();
 sg13g2_fill_2 FILLER_70_473 ();
 sg13g2_fill_2 FILLER_70_484 ();
 sg13g2_decap_8 FILLER_70_495 ();
 sg13g2_fill_2 FILLER_70_502 ();
 sg13g2_fill_2 FILLER_70_508 ();
 sg13g2_decap_4 FILLER_70_515 ();
 sg13g2_decap_8 FILLER_70_536 ();
 sg13g2_fill_2 FILLER_70_543 ();
 sg13g2_decap_4 FILLER_70_554 ();
 sg13g2_decap_8 FILLER_70_571 ();
 sg13g2_fill_2 FILLER_70_601 ();
 sg13g2_fill_1 FILLER_70_608 ();
 sg13g2_fill_1 FILLER_70_617 ();
 sg13g2_decap_4 FILLER_70_626 ();
 sg13g2_fill_2 FILLER_70_630 ();
 sg13g2_fill_2 FILLER_70_660 ();
 sg13g2_decap_4 FILLER_70_683 ();
 sg13g2_fill_1 FILLER_70_691 ();
 sg13g2_decap_8 FILLER_70_701 ();
 sg13g2_fill_1 FILLER_70_708 ();
 sg13g2_fill_2 FILLER_70_722 ();
 sg13g2_decap_8 FILLER_70_758 ();
 sg13g2_decap_8 FILLER_70_765 ();
 sg13g2_decap_8 FILLER_70_772 ();
 sg13g2_decap_8 FILLER_70_779 ();
 sg13g2_decap_8 FILLER_70_786 ();
 sg13g2_decap_8 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_800 ();
 sg13g2_decap_8 FILLER_70_807 ();
 sg13g2_decap_8 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_821 ();
 sg13g2_decap_8 FILLER_70_828 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_4 FILLER_71_116 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_decap_8 FILLER_71_134 ();
 sg13g2_decap_4 FILLER_71_141 ();
 sg13g2_fill_2 FILLER_71_171 ();
 sg13g2_fill_2 FILLER_71_183 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_decap_8 FILLER_71_201 ();
 sg13g2_fill_2 FILLER_71_208 ();
 sg13g2_decap_8 FILLER_71_233 ();
 sg13g2_decap_4 FILLER_71_240 ();
 sg13g2_fill_1 FILLER_71_244 ();
 sg13g2_decap_4 FILLER_71_255 ();
 sg13g2_fill_2 FILLER_71_267 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_4 FILLER_71_280 ();
 sg13g2_fill_2 FILLER_71_284 ();
 sg13g2_fill_2 FILLER_71_302 ();
 sg13g2_fill_1 FILLER_71_304 ();
 sg13g2_fill_2 FILLER_71_311 ();
 sg13g2_fill_1 FILLER_71_313 ();
 sg13g2_decap_8 FILLER_71_330 ();
 sg13g2_decap_4 FILLER_71_337 ();
 sg13g2_fill_2 FILLER_71_359 ();
 sg13g2_fill_1 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_fill_1 FILLER_71_389 ();
 sg13g2_fill_2 FILLER_71_403 ();
 sg13g2_fill_1 FILLER_71_405 ();
 sg13g2_decap_4 FILLER_71_413 ();
 sg13g2_fill_2 FILLER_71_417 ();
 sg13g2_decap_8 FILLER_71_431 ();
 sg13g2_decap_8 FILLER_71_438 ();
 sg13g2_decap_4 FILLER_71_445 ();
 sg13g2_fill_1 FILLER_71_449 ();
 sg13g2_decap_4 FILLER_71_466 ();
 sg13g2_fill_1 FILLER_71_522 ();
 sg13g2_fill_1 FILLER_71_545 ();
 sg13g2_decap_8 FILLER_71_572 ();
 sg13g2_fill_1 FILLER_71_579 ();
 sg13g2_decap_8 FILLER_71_597 ();
 sg13g2_fill_2 FILLER_71_604 ();
 sg13g2_decap_8 FILLER_71_614 ();
 sg13g2_decap_4 FILLER_71_621 ();
 sg13g2_fill_2 FILLER_71_625 ();
 sg13g2_fill_2 FILLER_71_670 ();
 sg13g2_decap_8 FILLER_71_740 ();
 sg13g2_decap_8 FILLER_71_747 ();
 sg13g2_decap_8 FILLER_71_754 ();
 sg13g2_decap_8 FILLER_71_761 ();
 sg13g2_decap_8 FILLER_71_768 ();
 sg13g2_decap_8 FILLER_71_775 ();
 sg13g2_decap_8 FILLER_71_782 ();
 sg13g2_decap_8 FILLER_71_789 ();
 sg13g2_decap_8 FILLER_71_796 ();
 sg13g2_decap_8 FILLER_71_803 ();
 sg13g2_decap_8 FILLER_71_810 ();
 sg13g2_decap_8 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_824 ();
 sg13g2_decap_8 FILLER_71_831 ();
 sg13g2_decap_8 FILLER_71_838 ();
 sg13g2_decap_8 FILLER_71_845 ();
 sg13g2_decap_8 FILLER_71_852 ();
 sg13g2_fill_2 FILLER_71_859 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_91 ();
 sg13g2_fill_1 FILLER_72_93 ();
 sg13g2_fill_2 FILLER_72_100 ();
 sg13g2_decap_8 FILLER_72_114 ();
 sg13g2_fill_2 FILLER_72_121 ();
 sg13g2_fill_1 FILLER_72_123 ();
 sg13g2_fill_2 FILLER_72_129 ();
 sg13g2_fill_1 FILLER_72_131 ();
 sg13g2_decap_8 FILLER_72_142 ();
 sg13g2_decap_8 FILLER_72_153 ();
 sg13g2_fill_2 FILLER_72_160 ();
 sg13g2_decap_8 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_174 ();
 sg13g2_decap_4 FILLER_72_181 ();
 sg13g2_fill_1 FILLER_72_185 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_fill_2 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_4 FILLER_72_224 ();
 sg13g2_fill_1 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_234 ();
 sg13g2_fill_2 FILLER_72_247 ();
 sg13g2_fill_2 FILLER_72_257 ();
 sg13g2_fill_1 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_4 FILLER_72_280 ();
 sg13g2_decap_4 FILLER_72_300 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_decap_8 FILLER_72_323 ();
 sg13g2_decap_8 FILLER_72_335 ();
 sg13g2_decap_8 FILLER_72_342 ();
 sg13g2_decap_4 FILLER_72_349 ();
 sg13g2_fill_1 FILLER_72_353 ();
 sg13g2_decap_4 FILLER_72_359 ();
 sg13g2_fill_1 FILLER_72_363 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_fill_1 FILLER_72_385 ();
 sg13g2_decap_4 FILLER_72_391 ();
 sg13g2_fill_1 FILLER_72_395 ();
 sg13g2_fill_2 FILLER_72_409 ();
 sg13g2_decap_8 FILLER_72_418 ();
 sg13g2_decap_8 FILLER_72_443 ();
 sg13g2_decap_4 FILLER_72_450 ();
 sg13g2_fill_2 FILLER_72_454 ();
 sg13g2_decap_8 FILLER_72_466 ();
 sg13g2_fill_1 FILLER_72_473 ();
 sg13g2_fill_2 FILLER_72_478 ();
 sg13g2_fill_1 FILLER_72_480 ();
 sg13g2_fill_1 FILLER_72_485 ();
 sg13g2_decap_8 FILLER_72_495 ();
 sg13g2_decap_8 FILLER_72_502 ();
 sg13g2_fill_1 FILLER_72_509 ();
 sg13g2_fill_1 FILLER_72_515 ();
 sg13g2_fill_2 FILLER_72_521 ();
 sg13g2_fill_1 FILLER_72_523 ();
 sg13g2_fill_2 FILLER_72_536 ();
 sg13g2_decap_8 FILLER_72_543 ();
 sg13g2_decap_4 FILLER_72_550 ();
 sg13g2_fill_2 FILLER_72_554 ();
 sg13g2_decap_4 FILLER_72_592 ();
 sg13g2_fill_1 FILLER_72_596 ();
 sg13g2_decap_8 FILLER_72_601 ();
 sg13g2_decap_4 FILLER_72_608 ();
 sg13g2_fill_2 FILLER_72_612 ();
 sg13g2_fill_2 FILLER_72_618 ();
 sg13g2_fill_2 FILLER_72_626 ();
 sg13g2_fill_2 FILLER_72_641 ();
 sg13g2_fill_2 FILLER_72_658 ();
 sg13g2_fill_2 FILLER_72_674 ();
 sg13g2_decap_8 FILLER_72_702 ();
 sg13g2_decap_8 FILLER_72_709 ();
 sg13g2_decap_8 FILLER_72_716 ();
 sg13g2_decap_8 FILLER_72_723 ();
 sg13g2_decap_8 FILLER_72_730 ();
 sg13g2_decap_8 FILLER_72_737 ();
 sg13g2_decap_8 FILLER_72_744 ();
 sg13g2_decap_8 FILLER_72_751 ();
 sg13g2_decap_8 FILLER_72_758 ();
 sg13g2_decap_8 FILLER_72_765 ();
 sg13g2_decap_8 FILLER_72_772 ();
 sg13g2_decap_8 FILLER_72_779 ();
 sg13g2_decap_8 FILLER_72_786 ();
 sg13g2_decap_8 FILLER_72_793 ();
 sg13g2_decap_8 FILLER_72_800 ();
 sg13g2_decap_8 FILLER_72_807 ();
 sg13g2_decap_8 FILLER_72_814 ();
 sg13g2_decap_8 FILLER_72_821 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_4 FILLER_72_856 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_4 FILLER_73_70 ();
 sg13g2_fill_2 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_86 ();
 sg13g2_decap_4 FILLER_73_104 ();
 sg13g2_fill_2 FILLER_73_125 ();
 sg13g2_fill_1 FILLER_73_127 ();
 sg13g2_decap_8 FILLER_73_148 ();
 sg13g2_fill_2 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_fill_1 FILLER_73_225 ();
 sg13g2_fill_1 FILLER_73_235 ();
 sg13g2_decap_8 FILLER_73_243 ();
 sg13g2_decap_8 FILLER_73_250 ();
 sg13g2_fill_2 FILLER_73_257 ();
 sg13g2_fill_2 FILLER_73_274 ();
 sg13g2_fill_1 FILLER_73_276 ();
 sg13g2_decap_8 FILLER_73_288 ();
 sg13g2_decap_4 FILLER_73_295 ();
 sg13g2_decap_8 FILLER_73_319 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_decap_8 FILLER_73_345 ();
 sg13g2_decap_8 FILLER_73_352 ();
 sg13g2_fill_1 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_fill_1 FILLER_73_405 ();
 sg13g2_decap_4 FILLER_73_412 ();
 sg13g2_fill_1 FILLER_73_416 ();
 sg13g2_decap_8 FILLER_73_422 ();
 sg13g2_fill_2 FILLER_73_429 ();
 sg13g2_fill_1 FILLER_73_431 ();
 sg13g2_fill_2 FILLER_73_445 ();
 sg13g2_fill_1 FILLER_73_447 ();
 sg13g2_decap_8 FILLER_73_471 ();
 sg13g2_decap_8 FILLER_73_478 ();
 sg13g2_fill_2 FILLER_73_485 ();
 sg13g2_fill_1 FILLER_73_511 ();
 sg13g2_fill_2 FILLER_73_527 ();
 sg13g2_fill_2 FILLER_73_549 ();
 sg13g2_fill_1 FILLER_73_551 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_585 ();
 sg13g2_decap_4 FILLER_73_592 ();
 sg13g2_fill_1 FILLER_73_612 ();
 sg13g2_fill_1 FILLER_73_621 ();
 sg13g2_fill_2 FILLER_73_677 ();
 sg13g2_fill_1 FILLER_73_679 ();
 sg13g2_decap_8 FILLER_73_698 ();
 sg13g2_decap_8 FILLER_73_705 ();
 sg13g2_decap_8 FILLER_73_712 ();
 sg13g2_decap_8 FILLER_73_719 ();
 sg13g2_decap_8 FILLER_73_726 ();
 sg13g2_decap_8 FILLER_73_733 ();
 sg13g2_decap_8 FILLER_73_740 ();
 sg13g2_decap_8 FILLER_73_747 ();
 sg13g2_decap_8 FILLER_73_754 ();
 sg13g2_decap_8 FILLER_73_761 ();
 sg13g2_decap_8 FILLER_73_768 ();
 sg13g2_decap_8 FILLER_73_775 ();
 sg13g2_decap_8 FILLER_73_782 ();
 sg13g2_decap_8 FILLER_73_789 ();
 sg13g2_decap_8 FILLER_73_796 ();
 sg13g2_decap_8 FILLER_73_803 ();
 sg13g2_decap_8 FILLER_73_810 ();
 sg13g2_decap_8 FILLER_73_817 ();
 sg13g2_decap_8 FILLER_73_824 ();
 sg13g2_decap_8 FILLER_73_831 ();
 sg13g2_decap_8 FILLER_73_838 ();
 sg13g2_decap_8 FILLER_73_845 ();
 sg13g2_decap_8 FILLER_73_852 ();
 sg13g2_fill_2 FILLER_73_859 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_4 FILLER_74_63 ();
 sg13g2_fill_2 FILLER_74_67 ();
 sg13g2_fill_1 FILLER_74_92 ();
 sg13g2_fill_1 FILLER_74_97 ();
 sg13g2_decap_8 FILLER_74_108 ();
 sg13g2_decap_8 FILLER_74_115 ();
 sg13g2_decap_8 FILLER_74_122 ();
 sg13g2_decap_4 FILLER_74_129 ();
 sg13g2_fill_1 FILLER_74_133 ();
 sg13g2_decap_4 FILLER_74_142 ();
 sg13g2_fill_1 FILLER_74_146 ();
 sg13g2_decap_8 FILLER_74_155 ();
 sg13g2_decap_8 FILLER_74_167 ();
 sg13g2_decap_4 FILLER_74_174 ();
 sg13g2_fill_2 FILLER_74_178 ();
 sg13g2_fill_2 FILLER_74_186 ();
 sg13g2_fill_1 FILLER_74_188 ();
 sg13g2_decap_8 FILLER_74_193 ();
 sg13g2_fill_2 FILLER_74_200 ();
 sg13g2_decap_8 FILLER_74_211 ();
 sg13g2_decap_8 FILLER_74_218 ();
 sg13g2_decap_8 FILLER_74_225 ();
 sg13g2_decap_4 FILLER_74_249 ();
 sg13g2_decap_8 FILLER_74_260 ();
 sg13g2_decap_4 FILLER_74_267 ();
 sg13g2_fill_1 FILLER_74_271 ();
 sg13g2_decap_8 FILLER_74_293 ();
 sg13g2_fill_2 FILLER_74_300 ();
 sg13g2_decap_8 FILLER_74_314 ();
 sg13g2_decap_4 FILLER_74_321 ();
 sg13g2_fill_1 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_360 ();
 sg13g2_decap_8 FILLER_74_367 ();
 sg13g2_fill_2 FILLER_74_374 ();
 sg13g2_fill_1 FILLER_74_376 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_fill_2 FILLER_74_405 ();
 sg13g2_decap_4 FILLER_74_414 ();
 sg13g2_fill_1 FILLER_74_418 ();
 sg13g2_decap_8 FILLER_74_439 ();
 sg13g2_decap_8 FILLER_74_463 ();
 sg13g2_decap_4 FILLER_74_470 ();
 sg13g2_fill_2 FILLER_74_474 ();
 sg13g2_decap_4 FILLER_74_502 ();
 sg13g2_fill_1 FILLER_74_506 ();
 sg13g2_fill_2 FILLER_74_512 ();
 sg13g2_fill_1 FILLER_74_514 ();
 sg13g2_decap_8 FILLER_74_524 ();
 sg13g2_decap_8 FILLER_74_531 ();
 sg13g2_fill_2 FILLER_74_538 ();
 sg13g2_fill_1 FILLER_74_549 ();
 sg13g2_fill_1 FILLER_74_562 ();
 sg13g2_fill_2 FILLER_74_567 ();
 sg13g2_decap_4 FILLER_74_583 ();
 sg13g2_decap_4 FILLER_74_615 ();
 sg13g2_decap_8 FILLER_74_622 ();
 sg13g2_decap_8 FILLER_74_629 ();
 sg13g2_fill_2 FILLER_74_636 ();
 sg13g2_fill_1 FILLER_74_647 ();
 sg13g2_decap_8 FILLER_74_651 ();
 sg13g2_fill_1 FILLER_74_658 ();
 sg13g2_decap_8 FILLER_74_663 ();
 sg13g2_decap_8 FILLER_74_670 ();
 sg13g2_decap_8 FILLER_74_677 ();
 sg13g2_decap_8 FILLER_74_684 ();
 sg13g2_decap_8 FILLER_74_691 ();
 sg13g2_decap_8 FILLER_74_698 ();
 sg13g2_decap_8 FILLER_74_705 ();
 sg13g2_decap_8 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_719 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_740 ();
 sg13g2_decap_8 FILLER_74_747 ();
 sg13g2_decap_8 FILLER_74_754 ();
 sg13g2_decap_8 FILLER_74_761 ();
 sg13g2_decap_8 FILLER_74_768 ();
 sg13g2_decap_8 FILLER_74_775 ();
 sg13g2_decap_8 FILLER_74_782 ();
 sg13g2_decap_8 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_796 ();
 sg13g2_decap_8 FILLER_74_803 ();
 sg13g2_decap_8 FILLER_74_810 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_8 FILLER_74_824 ();
 sg13g2_decap_8 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_77 ();
 sg13g2_fill_2 FILLER_75_92 ();
 sg13g2_decap_4 FILLER_75_99 ();
 sg13g2_decap_4 FILLER_75_128 ();
 sg13g2_fill_1 FILLER_75_137 ();
 sg13g2_decap_4 FILLER_75_154 ();
 sg13g2_fill_2 FILLER_75_158 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_decap_4 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_186 ();
 sg13g2_decap_4 FILLER_75_195 ();
 sg13g2_fill_2 FILLER_75_202 ();
 sg13g2_fill_1 FILLER_75_204 ();
 sg13g2_decap_8 FILLER_75_209 ();
 sg13g2_decap_4 FILLER_75_216 ();
 sg13g2_fill_1 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_246 ();
 sg13g2_decap_8 FILLER_75_268 ();
 sg13g2_decap_8 FILLER_75_275 ();
 sg13g2_fill_1 FILLER_75_282 ();
 sg13g2_decap_4 FILLER_75_300 ();
 sg13g2_fill_2 FILLER_75_304 ();
 sg13g2_decap_4 FILLER_75_310 ();
 sg13g2_fill_2 FILLER_75_314 ();
 sg13g2_decap_8 FILLER_75_334 ();
 sg13g2_decap_8 FILLER_75_341 ();
 sg13g2_fill_2 FILLER_75_366 ();
 sg13g2_fill_1 FILLER_75_368 ();
 sg13g2_fill_2 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_fill_2 FILLER_75_398 ();
 sg13g2_fill_1 FILLER_75_400 ();
 sg13g2_decap_8 FILLER_75_414 ();
 sg13g2_fill_2 FILLER_75_421 ();
 sg13g2_fill_2 FILLER_75_433 ();
 sg13g2_fill_1 FILLER_75_435 ();
 sg13g2_decap_4 FILLER_75_441 ();
 sg13g2_fill_1 FILLER_75_445 ();
 sg13g2_fill_2 FILLER_75_451 ();
 sg13g2_fill_1 FILLER_75_456 ();
 sg13g2_fill_1 FILLER_75_461 ();
 sg13g2_decap_8 FILLER_75_471 ();
 sg13g2_decap_8 FILLER_75_478 ();
 sg13g2_decap_8 FILLER_75_485 ();
 sg13g2_fill_2 FILLER_75_492 ();
 sg13g2_decap_8 FILLER_75_498 ();
 sg13g2_fill_2 FILLER_75_541 ();
 sg13g2_fill_2 FILLER_75_564 ();
 sg13g2_fill_2 FILLER_75_575 ();
 sg13g2_fill_1 FILLER_75_577 ();
 sg13g2_fill_1 FILLER_75_586 ();
 sg13g2_fill_1 FILLER_75_609 ();
 sg13g2_decap_8 FILLER_75_641 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_8 FILLER_75_655 ();
 sg13g2_decap_8 FILLER_75_662 ();
 sg13g2_decap_8 FILLER_75_669 ();
 sg13g2_decap_8 FILLER_75_676 ();
 sg13g2_decap_8 FILLER_75_683 ();
 sg13g2_decap_8 FILLER_75_690 ();
 sg13g2_decap_8 FILLER_75_697 ();
 sg13g2_decap_8 FILLER_75_704 ();
 sg13g2_decap_8 FILLER_75_711 ();
 sg13g2_decap_8 FILLER_75_718 ();
 sg13g2_decap_8 FILLER_75_725 ();
 sg13g2_decap_8 FILLER_75_732 ();
 sg13g2_decap_8 FILLER_75_739 ();
 sg13g2_decap_8 FILLER_75_746 ();
 sg13g2_decap_8 FILLER_75_753 ();
 sg13g2_decap_8 FILLER_75_760 ();
 sg13g2_decap_8 FILLER_75_767 ();
 sg13g2_decap_8 FILLER_75_774 ();
 sg13g2_decap_8 FILLER_75_781 ();
 sg13g2_decap_8 FILLER_75_788 ();
 sg13g2_decap_8 FILLER_75_795 ();
 sg13g2_decap_8 FILLER_75_802 ();
 sg13g2_decap_8 FILLER_75_809 ();
 sg13g2_decap_8 FILLER_75_816 ();
 sg13g2_decap_8 FILLER_75_823 ();
 sg13g2_decap_8 FILLER_75_830 ();
 sg13g2_decap_8 FILLER_75_837 ();
 sg13g2_decap_8 FILLER_75_844 ();
 sg13g2_decap_8 FILLER_75_851 ();
 sg13g2_decap_4 FILLER_75_858 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_101 ();
 sg13g2_decap_8 FILLER_76_116 ();
 sg13g2_fill_1 FILLER_76_123 ();
 sg13g2_fill_2 FILLER_76_152 ();
 sg13g2_fill_2 FILLER_76_159 ();
 sg13g2_fill_1 FILLER_76_176 ();
 sg13g2_decap_8 FILLER_76_187 ();
 sg13g2_decap_4 FILLER_76_194 ();
 sg13g2_fill_1 FILLER_76_198 ();
 sg13g2_decap_4 FILLER_76_238 ();
 sg13g2_fill_2 FILLER_76_242 ();
 sg13g2_decap_8 FILLER_76_272 ();
 sg13g2_decap_4 FILLER_76_279 ();
 sg13g2_fill_2 FILLER_76_283 ();
 sg13g2_fill_1 FILLER_76_302 ();
 sg13g2_fill_2 FILLER_76_316 ();
 sg13g2_fill_1 FILLER_76_318 ();
 sg13g2_fill_2 FILLER_76_326 ();
 sg13g2_decap_4 FILLER_76_333 ();
 sg13g2_fill_2 FILLER_76_337 ();
 sg13g2_fill_2 FILLER_76_358 ();
 sg13g2_fill_1 FILLER_76_360 ();
 sg13g2_fill_2 FILLER_76_371 ();
 sg13g2_fill_2 FILLER_76_384 ();
 sg13g2_fill_1 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_391 ();
 sg13g2_decap_4 FILLER_76_398 ();
 sg13g2_fill_2 FILLER_76_402 ();
 sg13g2_fill_2 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_426 ();
 sg13g2_decap_4 FILLER_76_433 ();
 sg13g2_fill_2 FILLER_76_437 ();
 sg13g2_fill_1 FILLER_76_449 ();
 sg13g2_decap_8 FILLER_76_476 ();
 sg13g2_fill_1 FILLER_76_544 ();
 sg13g2_fill_1 FILLER_76_553 ();
 sg13g2_fill_2 FILLER_76_559 ();
 sg13g2_fill_2 FILLER_76_589 ();
 sg13g2_fill_1 FILLER_76_626 ();
 sg13g2_decap_8 FILLER_76_636 ();
 sg13g2_decap_8 FILLER_76_643 ();
 sg13g2_decap_8 FILLER_76_650 ();
 sg13g2_decap_8 FILLER_76_657 ();
 sg13g2_decap_8 FILLER_76_664 ();
 sg13g2_decap_8 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_678 ();
 sg13g2_decap_8 FILLER_76_685 ();
 sg13g2_decap_8 FILLER_76_692 ();
 sg13g2_decap_8 FILLER_76_699 ();
 sg13g2_decap_8 FILLER_76_706 ();
 sg13g2_decap_8 FILLER_76_713 ();
 sg13g2_decap_8 FILLER_76_720 ();
 sg13g2_decap_8 FILLER_76_727 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_decap_8 FILLER_76_741 ();
 sg13g2_decap_8 FILLER_76_748 ();
 sg13g2_decap_8 FILLER_76_755 ();
 sg13g2_decap_8 FILLER_76_762 ();
 sg13g2_decap_8 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_776 ();
 sg13g2_decap_8 FILLER_76_783 ();
 sg13g2_decap_8 FILLER_76_790 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_804 ();
 sg13g2_decap_8 FILLER_76_811 ();
 sg13g2_decap_8 FILLER_76_818 ();
 sg13g2_decap_8 FILLER_76_825 ();
 sg13g2_decap_8 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_839 ();
 sg13g2_decap_8 FILLER_76_846 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_86 ();
 sg13g2_decap_8 FILLER_77_108 ();
 sg13g2_decap_8 FILLER_77_115 ();
 sg13g2_decap_8 FILLER_77_122 ();
 sg13g2_decap_8 FILLER_77_129 ();
 sg13g2_decap_4 FILLER_77_136 ();
 sg13g2_fill_1 FILLER_77_140 ();
 sg13g2_fill_2 FILLER_77_146 ();
 sg13g2_decap_8 FILLER_77_166 ();
 sg13g2_fill_1 FILLER_77_173 ();
 sg13g2_decap_8 FILLER_77_195 ();
 sg13g2_decap_4 FILLER_77_202 ();
 sg13g2_decap_8 FILLER_77_218 ();
 sg13g2_fill_1 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_237 ();
 sg13g2_decap_8 FILLER_77_244 ();
 sg13g2_fill_1 FILLER_77_251 ();
 sg13g2_decap_8 FILLER_77_268 ();
 sg13g2_decap_8 FILLER_77_275 ();
 sg13g2_decap_4 FILLER_77_282 ();
 sg13g2_fill_1 FILLER_77_286 ();
 sg13g2_decap_8 FILLER_77_305 ();
 sg13g2_decap_8 FILLER_77_312 ();
 sg13g2_fill_2 FILLER_77_326 ();
 sg13g2_fill_1 FILLER_77_328 ();
 sg13g2_decap_8 FILLER_77_338 ();
 sg13g2_fill_2 FILLER_77_345 ();
 sg13g2_decap_8 FILLER_77_352 ();
 sg13g2_decap_4 FILLER_77_364 ();
 sg13g2_decap_4 FILLER_77_377 ();
 sg13g2_fill_1 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_413 ();
 sg13g2_decap_4 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_443 ();
 sg13g2_decap_4 FILLER_77_450 ();
 sg13g2_fill_2 FILLER_77_454 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_476 ();
 sg13g2_decap_8 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_490 ();
 sg13g2_decap_8 FILLER_77_497 ();
 sg13g2_decap_4 FILLER_77_504 ();
 sg13g2_decap_8 FILLER_77_517 ();
 sg13g2_fill_2 FILLER_77_524 ();
 sg13g2_fill_1 FILLER_77_526 ();
 sg13g2_decap_8 FILLER_77_553 ();
 sg13g2_decap_8 FILLER_77_595 ();
 sg13g2_fill_2 FILLER_77_606 ();
 sg13g2_fill_1 FILLER_77_608 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_fill_1 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_630 ();
 sg13g2_decap_8 FILLER_77_637 ();
 sg13g2_decap_8 FILLER_77_644 ();
 sg13g2_decap_8 FILLER_77_651 ();
 sg13g2_decap_8 FILLER_77_658 ();
 sg13g2_decap_8 FILLER_77_665 ();
 sg13g2_decap_8 FILLER_77_672 ();
 sg13g2_decap_8 FILLER_77_679 ();
 sg13g2_decap_8 FILLER_77_686 ();
 sg13g2_decap_8 FILLER_77_693 ();
 sg13g2_decap_8 FILLER_77_700 ();
 sg13g2_decap_8 FILLER_77_707 ();
 sg13g2_decap_8 FILLER_77_714 ();
 sg13g2_decap_8 FILLER_77_721 ();
 sg13g2_decap_8 FILLER_77_728 ();
 sg13g2_decap_8 FILLER_77_735 ();
 sg13g2_decap_8 FILLER_77_742 ();
 sg13g2_decap_8 FILLER_77_749 ();
 sg13g2_decap_8 FILLER_77_756 ();
 sg13g2_decap_8 FILLER_77_763 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_decap_8 FILLER_77_791 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_4 FILLER_78_84 ();
 sg13g2_fill_2 FILLER_78_88 ();
 sg13g2_fill_2 FILLER_78_95 ();
 sg13g2_decap_8 FILLER_78_101 ();
 sg13g2_fill_1 FILLER_78_108 ();
 sg13g2_decap_8 FILLER_78_135 ();
 sg13g2_decap_8 FILLER_78_142 ();
 sg13g2_decap_4 FILLER_78_158 ();
 sg13g2_fill_1 FILLER_78_162 ();
 sg13g2_decap_4 FILLER_78_168 ();
 sg13g2_fill_1 FILLER_78_172 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_fill_2 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_4 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_fill_2 FILLER_78_287 ();
 sg13g2_fill_1 FILLER_78_289 ();
 sg13g2_decap_8 FILLER_78_295 ();
 sg13g2_decap_4 FILLER_78_302 ();
 sg13g2_fill_2 FILLER_78_324 ();
 sg13g2_fill_2 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_356 ();
 sg13g2_decap_4 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_78_380 ();
 sg13g2_decap_4 FILLER_78_387 ();
 sg13g2_decap_4 FILLER_78_396 ();
 sg13g2_fill_1 FILLER_78_400 ();
 sg13g2_fill_2 FILLER_78_415 ();
 sg13g2_fill_2 FILLER_78_431 ();
 sg13g2_fill_1 FILLER_78_433 ();
 sg13g2_fill_2 FILLER_78_452 ();
 sg13g2_decap_8 FILLER_78_470 ();
 sg13g2_decap_8 FILLER_78_477 ();
 sg13g2_decap_8 FILLER_78_484 ();
 sg13g2_decap_8 FILLER_78_491 ();
 sg13g2_decap_8 FILLER_78_498 ();
 sg13g2_decap_8 FILLER_78_505 ();
 sg13g2_decap_8 FILLER_78_512 ();
 sg13g2_decap_8 FILLER_78_519 ();
 sg13g2_decap_8 FILLER_78_526 ();
 sg13g2_decap_4 FILLER_78_533 ();
 sg13g2_decap_8 FILLER_78_550 ();
 sg13g2_decap_8 FILLER_78_557 ();
 sg13g2_decap_8 FILLER_78_564 ();
 sg13g2_decap_8 FILLER_78_579 ();
 sg13g2_decap_8 FILLER_78_586 ();
 sg13g2_decap_8 FILLER_78_593 ();
 sg13g2_decap_8 FILLER_78_600 ();
 sg13g2_decap_8 FILLER_78_607 ();
 sg13g2_decap_8 FILLER_78_614 ();
 sg13g2_decap_8 FILLER_78_621 ();
 sg13g2_decap_8 FILLER_78_628 ();
 sg13g2_decap_8 FILLER_78_635 ();
 sg13g2_decap_8 FILLER_78_642 ();
 sg13g2_decap_8 FILLER_78_649 ();
 sg13g2_decap_8 FILLER_78_656 ();
 sg13g2_decap_8 FILLER_78_663 ();
 sg13g2_decap_8 FILLER_78_670 ();
 sg13g2_decap_8 FILLER_78_677 ();
 sg13g2_decap_8 FILLER_78_684 ();
 sg13g2_decap_8 FILLER_78_691 ();
 sg13g2_decap_8 FILLER_78_698 ();
 sg13g2_decap_8 FILLER_78_705 ();
 sg13g2_decap_8 FILLER_78_712 ();
 sg13g2_decap_8 FILLER_78_719 ();
 sg13g2_decap_8 FILLER_78_726 ();
 sg13g2_decap_8 FILLER_78_733 ();
 sg13g2_decap_8 FILLER_78_740 ();
 sg13g2_decap_8 FILLER_78_747 ();
 sg13g2_decap_8 FILLER_78_754 ();
 sg13g2_decap_8 FILLER_78_761 ();
 sg13g2_decap_8 FILLER_78_768 ();
 sg13g2_decap_8 FILLER_78_775 ();
 sg13g2_decap_8 FILLER_78_782 ();
 sg13g2_decap_8 FILLER_78_789 ();
 sg13g2_decap_8 FILLER_78_796 ();
 sg13g2_decap_8 FILLER_78_803 ();
 sg13g2_decap_8 FILLER_78_810 ();
 sg13g2_decap_8 FILLER_78_817 ();
 sg13g2_decap_8 FILLER_78_824 ();
 sg13g2_decap_8 FILLER_78_831 ();
 sg13g2_decap_8 FILLER_78_838 ();
 sg13g2_decap_8 FILLER_78_845 ();
 sg13g2_decap_8 FILLER_78_852 ();
 sg13g2_fill_2 FILLER_78_859 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_fill_2 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_86 ();
 sg13g2_decap_8 FILLER_79_113 ();
 sg13g2_decap_8 FILLER_79_124 ();
 sg13g2_decap_8 FILLER_79_131 ();
 sg13g2_decap_8 FILLER_79_138 ();
 sg13g2_decap_8 FILLER_79_145 ();
 sg13g2_decap_4 FILLER_79_152 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_fill_2 FILLER_79_166 ();
 sg13g2_fill_1 FILLER_79_181 ();
 sg13g2_decap_8 FILLER_79_208 ();
 sg13g2_decap_8 FILLER_79_219 ();
 sg13g2_decap_4 FILLER_79_226 ();
 sg13g2_fill_2 FILLER_79_230 ();
 sg13g2_decap_4 FILLER_79_236 ();
 sg13g2_fill_2 FILLER_79_240 ();
 sg13g2_decap_4 FILLER_79_247 ();
 sg13g2_fill_2 FILLER_79_251 ();
 sg13g2_decap_8 FILLER_79_299 ();
 sg13g2_fill_2 FILLER_79_306 ();
 sg13g2_decap_4 FILLER_79_312 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_decap_8 FILLER_79_323 ();
 sg13g2_decap_4 FILLER_79_330 ();
 sg13g2_fill_2 FILLER_79_339 ();
 sg13g2_fill_1 FILLER_79_348 ();
 sg13g2_fill_1 FILLER_79_354 ();
 sg13g2_fill_2 FILLER_79_380 ();
 sg13g2_fill_1 FILLER_79_382 ();
 sg13g2_fill_1 FILLER_79_416 ();
 sg13g2_fill_2 FILLER_79_432 ();
 sg13g2_fill_1 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_445 ();
 sg13g2_fill_1 FILLER_79_452 ();
 sg13g2_decap_8 FILLER_79_458 ();
 sg13g2_decap_8 FILLER_79_465 ();
 sg13g2_decap_8 FILLER_79_472 ();
 sg13g2_decap_8 FILLER_79_479 ();
 sg13g2_decap_8 FILLER_79_486 ();
 sg13g2_decap_8 FILLER_79_493 ();
 sg13g2_decap_8 FILLER_79_500 ();
 sg13g2_decap_8 FILLER_79_507 ();
 sg13g2_decap_8 FILLER_79_514 ();
 sg13g2_decap_8 FILLER_79_521 ();
 sg13g2_decap_8 FILLER_79_528 ();
 sg13g2_decap_8 FILLER_79_535 ();
 sg13g2_decap_8 FILLER_79_542 ();
 sg13g2_decap_8 FILLER_79_549 ();
 sg13g2_decap_8 FILLER_79_556 ();
 sg13g2_decap_8 FILLER_79_563 ();
 sg13g2_decap_8 FILLER_79_570 ();
 sg13g2_decap_8 FILLER_79_577 ();
 sg13g2_decap_8 FILLER_79_584 ();
 sg13g2_decap_8 FILLER_79_591 ();
 sg13g2_decap_8 FILLER_79_598 ();
 sg13g2_decap_8 FILLER_79_605 ();
 sg13g2_decap_8 FILLER_79_612 ();
 sg13g2_decap_8 FILLER_79_619 ();
 sg13g2_decap_8 FILLER_79_626 ();
 sg13g2_decap_8 FILLER_79_633 ();
 sg13g2_decap_8 FILLER_79_640 ();
 sg13g2_decap_8 FILLER_79_647 ();
 sg13g2_decap_8 FILLER_79_654 ();
 sg13g2_decap_8 FILLER_79_661 ();
 sg13g2_decap_8 FILLER_79_668 ();
 sg13g2_decap_8 FILLER_79_675 ();
 sg13g2_decap_8 FILLER_79_682 ();
 sg13g2_decap_8 FILLER_79_689 ();
 sg13g2_decap_8 FILLER_79_696 ();
 sg13g2_decap_8 FILLER_79_703 ();
 sg13g2_decap_8 FILLER_79_710 ();
 sg13g2_decap_8 FILLER_79_717 ();
 sg13g2_decap_8 FILLER_79_724 ();
 sg13g2_decap_8 FILLER_79_731 ();
 sg13g2_decap_8 FILLER_79_738 ();
 sg13g2_decap_8 FILLER_79_745 ();
 sg13g2_decap_8 FILLER_79_752 ();
 sg13g2_decap_8 FILLER_79_759 ();
 sg13g2_decap_8 FILLER_79_766 ();
 sg13g2_decap_8 FILLER_79_773 ();
 sg13g2_decap_8 FILLER_79_780 ();
 sg13g2_decap_8 FILLER_79_787 ();
 sg13g2_decap_8 FILLER_79_794 ();
 sg13g2_decap_8 FILLER_79_801 ();
 sg13g2_decap_8 FILLER_79_808 ();
 sg13g2_decap_8 FILLER_79_815 ();
 sg13g2_decap_8 FILLER_79_822 ();
 sg13g2_decap_8 FILLER_79_829 ();
 sg13g2_decap_8 FILLER_79_836 ();
 sg13g2_decap_8 FILLER_79_843 ();
 sg13g2_decap_8 FILLER_79_850 ();
 sg13g2_decap_4 FILLER_79_857 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_fill_2 FILLER_80_132 ();
 sg13g2_fill_1 FILLER_80_134 ();
 sg13g2_decap_8 FILLER_80_186 ();
 sg13g2_decap_8 FILLER_80_197 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_decap_8 FILLER_80_274 ();
 sg13g2_fill_2 FILLER_80_281 ();
 sg13g2_fill_1 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_fill_2 FILLER_80_341 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_decap_4 FILLER_80_349 ();
 sg13g2_decap_8 FILLER_80_358 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_4 FILLER_80_401 ();
 sg13g2_fill_2 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_417 ();
 sg13g2_decap_8 FILLER_80_424 ();
 sg13g2_decap_4 FILLER_80_431 ();
 sg13g2_decap_8 FILLER_80_440 ();
 sg13g2_decap_8 FILLER_80_447 ();
 sg13g2_fill_2 FILLER_80_454 ();
 sg13g2_decap_8 FILLER_80_461 ();
 sg13g2_decap_8 FILLER_80_468 ();
 sg13g2_decap_8 FILLER_80_475 ();
 sg13g2_decap_8 FILLER_80_482 ();
 sg13g2_decap_8 FILLER_80_489 ();
 sg13g2_decap_8 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_503 ();
 sg13g2_decap_8 FILLER_80_510 ();
 sg13g2_decap_8 FILLER_80_517 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_decap_8 FILLER_80_531 ();
 sg13g2_decap_8 FILLER_80_538 ();
 sg13g2_decap_8 FILLER_80_545 ();
 sg13g2_decap_8 FILLER_80_552 ();
 sg13g2_decap_8 FILLER_80_559 ();
 sg13g2_decap_8 FILLER_80_566 ();
 sg13g2_decap_8 FILLER_80_573 ();
 sg13g2_decap_8 FILLER_80_580 ();
 sg13g2_decap_8 FILLER_80_587 ();
 sg13g2_decap_8 FILLER_80_594 ();
 sg13g2_decap_8 FILLER_80_601 ();
 sg13g2_decap_8 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_615 ();
 sg13g2_decap_8 FILLER_80_622 ();
 sg13g2_decap_8 FILLER_80_629 ();
 sg13g2_decap_8 FILLER_80_636 ();
 sg13g2_decap_8 FILLER_80_643 ();
 sg13g2_decap_8 FILLER_80_650 ();
 sg13g2_decap_8 FILLER_80_657 ();
 sg13g2_decap_8 FILLER_80_664 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_685 ();
 sg13g2_decap_8 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_720 ();
 sg13g2_decap_8 FILLER_80_727 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_8 FILLER_80_741 ();
 sg13g2_decap_8 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_797 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net164;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule
