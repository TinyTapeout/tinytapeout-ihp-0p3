module tt_um_algofoogle_fun_vga_clock (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire \clock_color_offset[0] ;
 wire \clock_color_offset[1] ;
 wire \clock_color_offset[2] ;
 wire \clock_hrs_d[0] ;
 wire \clock_hrs_d[1] ;
 wire \clock_hrs_u[0] ;
 wire \clock_hrs_u[1] ;
 wire \clock_hrs_u[2] ;
 wire \clock_hrs_u[3] ;
 wire \clock_min_d[0] ;
 wire \clock_min_d[1] ;
 wire \clock_min_d[2] ;
 wire \clock_min_u[0] ;
 wire \clock_min_u[1] ;
 wire \clock_min_u[2] ;
 wire \clock_min_u[3] ;
 wire \clock_sec_d[0] ;
 wire \clock_sec_d[1] ;
 wire \clock_sec_d[2] ;
 wire \clock_sec_u[0] ;
 wire \clock_sec_u[1] ;
 wire \clock_sec_u[2] ;
 wire \clock_sec_u[3] ;
 wire dx;
 wire \h[0] ;
 wire \h[1] ;
 wire \h[2] ;
 wire \h[3] ;
 wire \h[4] ;
 wire \h[5] ;
 wire hblank;
 wire hmax;
 wire \matt_venn_clock.pulse_hrs.comp[0] ;
 wire \matt_venn_clock.pulse_hrs.comp[1] ;
 wire \matt_venn_clock.pulse_hrs.comp[2] ;
 wire \matt_venn_clock.pulse_hrs.comp[3] ;
 wire \matt_venn_clock.pulse_hrs.comp[4] ;
 wire \matt_venn_clock.pulse_hrs.count[0] ;
 wire \matt_venn_clock.pulse_hrs.count[1] ;
 wire \matt_venn_clock.pulse_hrs.count[2] ;
 wire \matt_venn_clock.pulse_hrs.count[3] ;
 wire \matt_venn_clock.pulse_hrs.count[4] ;
 wire \matt_venn_clock.pulse_min.comp[0] ;
 wire \matt_venn_clock.pulse_min.comp[1] ;
 wire \matt_venn_clock.pulse_min.comp[2] ;
 wire \matt_venn_clock.pulse_min.comp[3] ;
 wire \matt_venn_clock.pulse_min.comp[4] ;
 wire \matt_venn_clock.pulse_min.count[0] ;
 wire \matt_venn_clock.pulse_min.count[1] ;
 wire \matt_venn_clock.pulse_min.count[2] ;
 wire \matt_venn_clock.pulse_min.count[3] ;
 wire \matt_venn_clock.pulse_min.count[4] ;
 wire \matt_venn_clock.pulse_sec.comp[0] ;
 wire \matt_venn_clock.pulse_sec.comp[1] ;
 wire \matt_venn_clock.pulse_sec.comp[2] ;
 wire \matt_venn_clock.pulse_sec.comp[3] ;
 wire \matt_venn_clock.pulse_sec.comp[4] ;
 wire \matt_venn_clock.pulse_sec.count[0] ;
 wire \matt_venn_clock.pulse_sec.count[1] ;
 wire \matt_venn_clock.pulse_sec.count[2] ;
 wire \matt_venn_clock.pulse_sec.count[3] ;
 wire \matt_venn_clock.pulse_sec.count[4] ;
 wire \matt_venn_clock.sec_counter[0] ;
 wire \matt_venn_clock.sec_counter[10] ;
 wire \matt_venn_clock.sec_counter[11] ;
 wire \matt_venn_clock.sec_counter[12] ;
 wire \matt_venn_clock.sec_counter[13] ;
 wire \matt_venn_clock.sec_counter[14] ;
 wire \matt_venn_clock.sec_counter[15] ;
 wire \matt_venn_clock.sec_counter[16] ;
 wire \matt_venn_clock.sec_counter[17] ;
 wire \matt_venn_clock.sec_counter[18] ;
 wire \matt_venn_clock.sec_counter[19] ;
 wire \matt_venn_clock.sec_counter[1] ;
 wire \matt_venn_clock.sec_counter[20] ;
 wire \matt_venn_clock.sec_counter[21] ;
 wire \matt_venn_clock.sec_counter[22] ;
 wire \matt_venn_clock.sec_counter[23] ;
 wire \matt_venn_clock.sec_counter[24] ;
 wire \matt_venn_clock.sec_counter[2] ;
 wire \matt_venn_clock.sec_counter[3] ;
 wire \matt_venn_clock.sec_counter[4] ;
 wire \matt_venn_clock.sec_counter[5] ;
 wire \matt_venn_clock.sec_counter[6] ;
 wire \matt_venn_clock.sec_counter[7] ;
 wire \matt_venn_clock.sec_counter[8] ;
 wire \matt_venn_clock.sec_counter[9] ;
 wire \matt_venn_vga.activevideo ;
 wire \matt_venn_vga.col_index[0] ;
 wire \matt_venn_vga.col_index[1] ;
 wire \matt_venn_vga.col_index_q[0] ;
 wire \matt_venn_vga.col_index_q[1] ;
 wire \matt_venn_vga.color[0] ;
 wire \matt_venn_vga.color[1] ;
 wire \matt_venn_vga.color[2] ;
 wire \matt_venn_vga.color[3] ;
 wire \matt_venn_vga.color[4] ;
 wire \matt_venn_vga.color[5] ;
 wire \matt_venn_vga.digit_0.char[0] ;
 wire \matt_venn_vga.digit_0.digit_index[0] ;
 wire \matt_venn_vga.digit_0.digit_index[1] ;
 wire \matt_venn_vga.digit_0.digit_index[2] ;
 wire \matt_venn_vga.digit_0.digit_index[3] ;
 wire \matt_venn_vga.digit_0.digit_index[4] ;
 wire \matt_venn_vga.digit_0.digit_index[5] ;
 wire \matt_venn_vga.draw ;
 wire \matt_venn_vga.font_0.dout[1] ;
 wire \matt_venn_vga.font_0.dout[2] ;
 wire \matt_venn_vga.font_0.dout[3] ;
 wire \matt_venn_vga.x_block_q[5] ;
 wire \matt_venn_vga.x_px[6] ;
 wire \matt_venn_vga.x_px[7] ;
 wire \matt_venn_vga.x_px[8] ;
 wire \matt_venn_vga.x_px[9] ;
 wire \matt_venn_vga.y_block_q[0] ;
 wire \matt_venn_vga.y_block_q[1] ;
 wire \matt_venn_vga.y_block_q[2] ;
 wire \matt_venn_vga.y_block_q[3] ;
 wire \matt_venn_vga.y_block_q[4] ;
 wire \matt_venn_vga.y_block_q[5] ;
 wire \matt_venn_vga.y_px[0] ;
 wire \matt_venn_vga.y_px[1] ;
 wire \matt_venn_vga.y_px[2] ;
 wire \matt_venn_vga.y_px[3] ;
 wire \matt_venn_vga.y_px[4] ;
 wire \matt_venn_vga.y_px[5] ;
 wire \matt_venn_vga.y_px[6] ;
 wire \matt_venn_vga.y_px[7] ;
 wire \matt_venn_vga.y_px[8] ;
 wire \matt_venn_vga.y_px[9] ;
 wire \matt_venn_vga_shadow.col_index[0] ;
 wire \matt_venn_vga_shadow.col_index[1] ;
 wire \matt_venn_vga_shadow.col_index_q[0] ;
 wire \matt_venn_vga_shadow.col_index_q[1] ;
 wire \matt_venn_vga_shadow.color[0] ;
 wire \matt_venn_vga_shadow.color[1] ;
 wire \matt_venn_vga_shadow.color[2] ;
 wire \matt_venn_vga_shadow.color[3] ;
 wire \matt_venn_vga_shadow.color[4] ;
 wire \matt_venn_vga_shadow.color[5] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[0] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[1] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[2] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[3] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[4] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[5] ;
 wire \matt_venn_vga_shadow.draw ;
 wire \matt_venn_vga_shadow.font_0.dout[1] ;
 wire \matt_venn_vga_shadow.font_0.dout[2] ;
 wire \matt_venn_vga_shadow.font_0.dout[3] ;
 wire \matt_venn_vga_shadow.x_block_q[5] ;
 wire \matt_venn_vga_shadow.y_block_q[0] ;
 wire \matt_venn_vga_shadow.y_block_q[1] ;
 wire \matt_venn_vga_shadow.y_block_q[2] ;
 wire \matt_venn_vga_shadow.y_block_q[3] ;
 wire \matt_venn_vga_shadow.y_block_q[4] ;
 wire \matt_venn_vga_shadow.y_block_q[5] ;
 wire \product_comp[0] ;
 wire \product_comp[10] ;
 wire \product_comp[1] ;
 wire \product_comp[2] ;
 wire \product_comp[3] ;
 wire \product_comp[4] ;
 wire \product_comp[5] ;
 wire \product_comp[6] ;
 wire \product_comp[7] ;
 wire \product_comp[8] ;
 wire \product_comp[9] ;
 wire \px[0] ;
 wire \px[1] ;
 wire \px[2] ;
 wire \px[3] ;
 wire \px[4] ;
 wire \px[5] ;
 wire \px[6] ;
 wire \px[7] ;
 wire \px[8] ;
 wire \px[9] ;
 wire \pxm[0] ;
 wire \pxm[1] ;
 wire \py[0] ;
 wire \py[1] ;
 wire \py[2] ;
 wire \py[3] ;
 wire \py[4] ;
 wire \py[5] ;
 wire \py[6] ;
 wire \py[7] ;
 wire \py[8] ;
 wire \py[9] ;
 wire \pym[10] ;
 wire \pym[11] ;
 wire \t[0] ;
 wire \t[1] ;
 wire \t[2] ;
 wire \t[3] ;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire clknet_leaf_0_clk;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire vblank;
 wire \vga_sync.hsync ;
 wire \vga_sync.o_vmax ;
 wire \vga_sync.vsync ;
 wire \ydelta[0] ;
 wire \ydelta[1] ;
 wire \ydelta[2] ;
 wire \ydelta[3] ;
 wire \ydelta[4] ;
 wire \ydelta[5] ;
 wire \ydelta[6] ;
 wire \ydelta[7] ;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;

 sg13g2_inv_1 _2195_ (.Y(_1349_),
    .A(net258));
 sg13g2_inv_1 _2196_ (.Y(_1350_),
    .A(\clock_min_d[1] ));
 sg13g2_inv_1 _2197_ (.Y(_1351_),
    .A(net425));
 sg13g2_inv_1 _2198_ (.Y(_1352_),
    .A(net228));
 sg13g2_inv_1 _2199_ (.Y(_1353_),
    .A(\matt_venn_clock.pulse_sec.count[4] ));
 sg13g2_inv_2 _2200_ (.Y(_1354_),
    .A(net248));
 sg13g2_inv_1 _2201_ (.Y(_1355_),
    .A(net427));
 sg13g2_inv_1 _2202_ (.Y(_1356_),
    .A(net373));
 sg13g2_inv_1 _2203_ (.Y(_1357_),
    .A(net443));
 sg13g2_inv_1 _2204_ (.Y(_1358_),
    .A(\matt_venn_clock.pulse_min.count[4] ));
 sg13g2_inv_1 _2205_ (.Y(_1359_),
    .A(net276));
 sg13g2_inv_1 _2206_ (.Y(_1360_),
    .A(\matt_venn_clock.pulse_min.count[1] ));
 sg13g2_inv_1 _2207_ (.Y(_1361_),
    .A(\matt_venn_clock.pulse_min.comp[4] ));
 sg13g2_inv_1 _2208_ (.Y(_1362_),
    .A(\matt_venn_clock.pulse_min.comp[3] ));
 sg13g2_inv_1 _2209_ (.Y(_1363_),
    .A(net418));
 sg13g2_inv_1 _2210_ (.Y(_1364_),
    .A(\matt_venn_clock.pulse_hrs.count[2] ));
 sg13g2_inv_1 _2211_ (.Y(_1365_),
    .A(\matt_venn_clock.pulse_hrs.count[1] ));
 sg13g2_inv_1 _2212_ (.Y(_1366_),
    .A(net450));
 sg13g2_inv_1 _2213_ (.Y(_1367_),
    .A(\matt_venn_clock.pulse_hrs.comp[1] ));
 sg13g2_inv_2 _2214_ (.Y(_1368_),
    .A(net323));
 sg13g2_inv_2 _2215_ (.Y(_1369_),
    .A(net328));
 sg13g2_inv_2 _2216_ (.Y(_1370_),
    .A(\matt_venn_vga.y_px[6] ));
 sg13g2_inv_1 _2217_ (.Y(_1371_),
    .A(net333));
 sg13g2_inv_4 _2218_ (.A(net334),
    .Y(_1372_));
 sg13g2_inv_1 _2219_ (.Y(_1373_),
    .A(net338));
 sg13g2_inv_2 _2220_ (.Y(_1374_),
    .A(net340));
 sg13g2_inv_2 _2221_ (.Y(_1375_),
    .A(dx));
 sg13g2_inv_1 _2222_ (.Y(_1376_),
    .A(\product_comp[10] ));
 sg13g2_inv_1 _2223_ (.Y(_1377_),
    .A(\product_comp[3] ));
 sg13g2_inv_1 _2224_ (.Y(_1378_),
    .A(net278));
 sg13g2_inv_1 _2225_ (.Y(_1379_),
    .A(net456));
 sg13g2_inv_1 _2226_ (.Y(_1380_),
    .A(\pym[10] ));
 sg13g2_inv_1 _2227_ (.Y(_1381_),
    .A(net513));
 sg13g2_inv_1 _2228_ (.Y(_1382_),
    .A(\py[6] ));
 sg13g2_inv_1 _2229_ (.Y(_1383_),
    .A(net548));
 sg13g2_inv_1 _2230_ (.Y(_1384_),
    .A(net350));
 sg13g2_inv_1 _2231_ (.Y(_1385_),
    .A(\px[2] ));
 sg13g2_inv_1 _2232_ (.Y(_1386_),
    .A(net354));
 sg13g2_inv_1 _2233_ (.Y(_1387_),
    .A(net355));
 sg13g2_inv_1 _2234_ (.Y(_1388_),
    .A(net475));
 sg13g2_inv_1 _2235_ (.Y(_1389_),
    .A(net498));
 sg13g2_inv_2 _2236_ (.Y(_1390_),
    .A(net550));
 sg13g2_inv_2 _2237_ (.Y(_1391_),
    .A(net312));
 sg13g2_inv_1 _2238_ (.Y(_1392_),
    .A(net318));
 sg13g2_inv_1 _2239_ (.Y(_1393_),
    .A(net556));
 sg13g2_inv_1 _2240_ (.Y(_1394_),
    .A(\h[1] ));
 sg13g2_inv_2 _2241_ (.Y(_1395_),
    .A(net6));
 sg13g2_inv_1 _2242_ (.Y(_1396_),
    .A(_0063_));
 sg13g2_inv_1 _2243_ (.Y(_1397_),
    .A(_0065_));
 sg13g2_inv_1 _2244_ (.Y(_1398_),
    .A(net370));
 sg13g2_inv_2 _2245_ (.Y(_1399_),
    .A(net3));
 sg13g2_inv_1 _2246_ (.Y(_1400_),
    .A(net2));
 sg13g2_inv_1 _2247_ (.Y(_1401_),
    .A(net1));
 sg13g2_inv_1 _2248_ (.Y(_1402_),
    .A(_0069_));
 sg13g2_inv_1 _2249_ (.Y(_1403_),
    .A(net361));
 sg13g2_inv_1 _2250_ (.Y(_1404_),
    .A(_0044_));
 sg13g2_inv_1 _2251_ (.Y(_1405_),
    .A(_0043_));
 sg13g2_inv_1 _2252_ (.Y(_1406_),
    .A(\matt_venn_vga.font_0.dout[2] ));
 sg13g2_inv_1 _2253_ (.Y(_1407_),
    .A(\matt_venn_vga.col_index_q[1] ));
 sg13g2_inv_1 _2254_ (.Y(_1408_),
    .A(\matt_venn_vga_shadow.font_0.dout[2] ));
 sg13g2_inv_1 _2255_ (.Y(_1409_),
    .A(\matt_venn_vga_shadow.col_index_q[1] ));
 sg13g2_nand2_1 _2256_ (.Y(_1410_),
    .A(net318),
    .B(net536));
 sg13g2_and2_1 _2257_ (.A(\h[0] ),
    .B(net532),
    .X(_1411_));
 sg13g2_nand2_2 _2258_ (.Y(_1412_),
    .A(net545),
    .B(net321));
 sg13g2_nor4_1 _2259_ (.A(net317),
    .B(_0055_),
    .C(_1410_),
    .D(_1412_),
    .Y(_1413_));
 sg13g2_nor2_1 _2260_ (.A(_1391_),
    .B(_1395_),
    .Y(_1414_));
 sg13g2_a21o_1 _2261_ (.A2(net310),
    .A1(\h[2] ),
    .B1(_1414_),
    .X(_1415_));
 sg13g2_nor2_2 _2262_ (.A(net313),
    .B(net558),
    .Y(_1416_));
 sg13g2_nand2_2 _2263_ (.Y(_1417_),
    .A(net313),
    .B(\matt_venn_vga.x_px[7] ));
 sg13g2_nand2b_2 _2264_ (.Y(_1418_),
    .B(_1417_),
    .A_N(_1416_));
 sg13g2_nand2_1 _2265_ (.Y(_1419_),
    .A(_1391_),
    .B(_1395_));
 sg13g2_o21ai_1 _2266_ (.B1(_1419_),
    .Y(_1420_),
    .A1(\h[2] ),
    .A2(net310));
 sg13g2_nand4_1 _2267_ (.B(_1415_),
    .C(_1418_),
    .A(_1413_),
    .Y(_1421_),
    .D(_1420_));
 sg13g2_inv_1 _2268_ (.Y(hmax),
    .A(_1421_));
 sg13g2_and2_1 _2269_ (.A(net335),
    .B(net337),
    .X(_1422_));
 sg13g2_nand2_2 _2270_ (.Y(_1423_),
    .A(net335),
    .B(net336));
 sg13g2_nor4_1 _2271_ (.A(net326),
    .B(\matt_venn_vga.y_px[7] ),
    .C(net331),
    .D(net6),
    .Y(_1424_));
 sg13g2_a21oi_1 _2272_ (.A1(_1422_),
    .A2(_1424_),
    .Y(_1425_),
    .B1(\matt_venn_vga.y_px[1] ));
 sg13g2_nand2_1 _2273_ (.Y(_1426_),
    .A(net339),
    .B(_1374_));
 sg13g2_xor2_1 _2274_ (.B(net340),
    .A(net338),
    .X(_1427_));
 sg13g2_nor4_1 _2275_ (.A(net329),
    .B(net333),
    .C(_0057_),
    .D(_1427_),
    .Y(_1428_));
 sg13g2_and2_2 _2276_ (.A(net325),
    .B(net328),
    .X(_1429_));
 sg13g2_nand2_1 _2277_ (.Y(_1430_),
    .A(net325),
    .B(net328));
 sg13g2_nor2_1 _2278_ (.A(net334),
    .B(net337),
    .Y(_1431_));
 sg13g2_nand4_1 _2279_ (.B(net6),
    .C(_1429_),
    .A(net331),
    .Y(_1432_),
    .D(_1431_));
 sg13g2_a21oi_1 _2280_ (.A1(\matt_venn_vga.y_px[1] ),
    .A2(_1432_),
    .Y(_1433_),
    .B1(_1425_));
 sg13g2_nand2_2 _2281_ (.Y(_1434_),
    .A(_1428_),
    .B(_1433_));
 sg13g2_inv_1 _2282_ (.Y(\vga_sync.o_vmax ),
    .A(_1434_));
 sg13g2_a21oi_1 _2283_ (.A1(net310),
    .A2(_1419_),
    .Y(_1435_),
    .B1(\matt_venn_vga.x_px[8] ));
 sg13g2_or2_1 _2284_ (.X(_1436_),
    .B(net319),
    .A(net318));
 sg13g2_nand4_1 _2285_ (.B(net316),
    .C(net6),
    .A(net314),
    .Y(_1437_),
    .D(_1436_));
 sg13g2_nor2_1 _2286_ (.A(net310),
    .B(_1414_),
    .Y(_1438_));
 sg13g2_a21oi_1 _2287_ (.A1(_1437_),
    .A2(_1438_),
    .Y(hblank),
    .B1(_1435_));
 sg13g2_nor2_2 _2288_ (.A(net330),
    .B(net332),
    .Y(_1439_));
 sg13g2_nor2_1 _2289_ (.A(net333),
    .B(net335),
    .Y(_1440_));
 sg13g2_nor4_2 _2290_ (.A(\matt_venn_vga.y_px[6] ),
    .B(net331),
    .C(net332),
    .Y(_1441_),
    .D(net335));
 sg13g2_nand2b_1 _2291_ (.Y(_1442_),
    .B(_1441_),
    .A_N(net337));
 sg13g2_nor2_2 _2292_ (.A(net338),
    .B(net340),
    .Y(_1443_));
 sg13g2_nor3_2 _2293_ (.A(net336),
    .B(net338),
    .C(net340),
    .Y(_1444_));
 sg13g2_and2_2 _2294_ (.A(_1372_),
    .B(_1444_),
    .X(_1445_));
 sg13g2_nand3_1 _2295_ (.B(_1429_),
    .C(_1442_),
    .A(net324),
    .Y(_1446_));
 sg13g2_and4_1 _2296_ (.A(net328),
    .B(net329),
    .C(net331),
    .D(_1371_),
    .X(_1447_));
 sg13g2_nand3_1 _2297_ (.B(_1445_),
    .C(_1447_),
    .A(net325),
    .Y(_1448_));
 sg13g2_nor2_1 _2298_ (.A(_1370_),
    .B(_0069_),
    .Y(_1449_));
 sg13g2_a21oi_1 _2299_ (.A1(_1429_),
    .A2(_1449_),
    .Y(_1450_),
    .B1(net324));
 sg13g2_a22oi_1 _2300_ (.Y(vblank),
    .B1(_1448_),
    .B2(_1450_),
    .A2(_1446_),
    .A1(net6));
 sg13g2_nor2_2 _2301_ (.A(hblank),
    .B(vblank),
    .Y(\matt_venn_vga.activevideo ));
 sg13g2_nand2_1 _2302_ (.Y(_1451_),
    .A(_0070_),
    .B(net361));
 sg13g2_nand2_2 _2303_ (.Y(_1452_),
    .A(_1403_),
    .B(\matt_venn_vga.activevideo ));
 sg13g2_inv_1 _2304_ (.Y(_1453_),
    .A(_1452_));
 sg13g2_nand3_1 _2305_ (.B(_1370_),
    .C(_1439_),
    .A(net328),
    .Y(_1454_));
 sg13g2_inv_1 _2306_ (.Y(_1455_),
    .A(_1454_));
 sg13g2_nor4_2 _2307_ (.A(_1369_),
    .B(net329),
    .C(net331),
    .Y(_1456_),
    .D(_1371_));
 sg13g2_nand2_1 _2308_ (.Y(_1457_),
    .A(net338),
    .B(net340));
 sg13g2_nand2_1 _2309_ (.Y(_1458_),
    .A(_1368_),
    .B(net325));
 sg13g2_nor2_1 _2310_ (.A(_1426_),
    .B(_1458_),
    .Y(_1459_));
 sg13g2_a21oi_1 _2311_ (.A1(net339),
    .A2(net341),
    .Y(_1460_),
    .B1(_1459_));
 sg13g2_o21ai_1 _2312_ (.B1(_1456_),
    .Y(_1461_),
    .A1(_1423_),
    .A2(_1460_));
 sg13g2_nand3_1 _2313_ (.B(net338),
    .C(net340),
    .A(net336),
    .Y(_1462_));
 sg13g2_nand3_1 _2314_ (.B(_1454_),
    .C(_1461_),
    .A(_1429_),
    .Y(_1463_));
 sg13g2_nand2_1 _2315_ (.Y(_1464_),
    .A(\t[0] ),
    .B(net322));
 sg13g2_xor2_1 _2316_ (.B(net321),
    .A(\t[1] ),
    .X(_1465_));
 sg13g2_nor2b_1 _2317_ (.A(_1464_),
    .B_N(_1465_),
    .Y(_1466_));
 sg13g2_a21oi_1 _2318_ (.A1(\t[1] ),
    .A2(net321),
    .Y(_1467_),
    .B1(_1466_));
 sg13g2_xor2_1 _2319_ (.B(net320),
    .A(\t[2] ),
    .X(_1468_));
 sg13g2_xnor2_1 _2320_ (.Y(_1469_),
    .A(net337),
    .B(_1468_));
 sg13g2_xnor2_1 _2321_ (.Y(_1470_),
    .A(_1467_),
    .B(_1469_));
 sg13g2_nand2_1 _2322_ (.Y(_1471_),
    .A(_1372_),
    .B(net337));
 sg13g2_o21ai_1 _2323_ (.B1(_0032_),
    .Y(_1472_),
    .A1(_1443_),
    .A2(_1471_));
 sg13g2_xnor2_1 _2324_ (.Y(_1473_),
    .A(_1371_),
    .B(_1472_));
 sg13g2_nand2_1 _2325_ (.Y(_1474_),
    .A(net330),
    .B(net332));
 sg13g2_a21oi_1 _2326_ (.A1(_1431_),
    .A2(_1457_),
    .Y(_1475_),
    .B1(_1474_));
 sg13g2_or2_1 _2327_ (.X(_1476_),
    .B(_1475_),
    .A(net329));
 sg13g2_xor2_1 _2328_ (.B(net322),
    .A(net341),
    .X(_1477_));
 sg13g2_xnor2_1 _2329_ (.Y(_1478_),
    .A(\t[0] ),
    .B(_1477_));
 sg13g2_a221oi_1 _2330_ (.B2(_1429_),
    .C1(_1478_),
    .B1(_1476_),
    .A1(_1470_),
    .Y(_1479_),
    .A2(_1473_));
 sg13g2_nor2_1 _2331_ (.A(_1463_),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_nor2_1 _2332_ (.A(net323),
    .B(_1480_),
    .Y(_1481_));
 sg13g2_inv_1 _2333_ (.Y(_1482_),
    .A(_1481_));
 sg13g2_nor2b_1 _2334_ (.A(net311),
    .B_N(\px[9] ),
    .Y(_1483_));
 sg13g2_nor2_1 _2335_ (.A(net349),
    .B(_1390_),
    .Y(_1484_));
 sg13g2_nand2_1 _2336_ (.Y(_1485_),
    .A(net349),
    .B(_1390_));
 sg13g2_nor2b_1 _2337_ (.A(_1484_),
    .B_N(_1485_),
    .Y(_1486_));
 sg13g2_nor2b_1 _2338_ (.A(net351),
    .B_N(net315),
    .Y(_1487_));
 sg13g2_nand2b_2 _2339_ (.Y(_1488_),
    .B(net351),
    .A_N(net315));
 sg13g2_nor2b_1 _2340_ (.A(_1487_),
    .B_N(_1488_),
    .Y(_1489_));
 sg13g2_nand2b_1 _2341_ (.Y(_1490_),
    .B(net317),
    .A_N(net352));
 sg13g2_nor2b_1 _2342_ (.A(\px[2] ),
    .B_N(net320),
    .Y(_1491_));
 sg13g2_nor2b_2 _2343_ (.A(\px[3] ),
    .B_N(net319),
    .Y(_1492_));
 sg13g2_xnor2_1 _2344_ (.Y(_1493_),
    .A(\px[3] ),
    .B(net319));
 sg13g2_and2_1 _2345_ (.A(_1491_),
    .B(_1493_),
    .X(_1494_));
 sg13g2_nand2b_1 _2346_ (.Y(_1495_),
    .B(net321),
    .A_N(net353));
 sg13g2_xnor2_1 _2347_ (.Y(_1496_),
    .A(\px[2] ),
    .B(net320));
 sg13g2_nand2b_1 _2348_ (.Y(_1497_),
    .B(_1496_),
    .A_N(_1495_));
 sg13g2_nand2b_1 _2349_ (.Y(_1498_),
    .B(\px[1] ),
    .A_N(net321));
 sg13g2_xor2_1 _2350_ (.B(net321),
    .A(\px[1] ),
    .X(_1499_));
 sg13g2_nand2b_1 _2351_ (.Y(_1500_),
    .B(net354),
    .A_N(net322));
 sg13g2_nor2b_1 _2352_ (.A(_1499_),
    .B_N(_1500_),
    .Y(_1501_));
 sg13g2_xnor2_1 _2353_ (.Y(_1502_),
    .A(_1495_),
    .B(_1496_));
 sg13g2_nand4_1 _2354_ (.B(_1496_),
    .C(_1498_),
    .A(_1495_),
    .Y(_1503_),
    .D(_1500_));
 sg13g2_xnor2_1 _2355_ (.Y(_1504_),
    .A(_1491_),
    .B(_1493_));
 sg13g2_a21oi_2 _2356_ (.B1(_1504_),
    .Y(_1505_),
    .A2(_1503_),
    .A1(_1497_));
 sg13g2_nand2_1 _2357_ (.Y(_1506_),
    .A(\px[4] ),
    .B(_1392_));
 sg13g2_xnor2_1 _2358_ (.Y(_1507_),
    .A(\px[4] ),
    .B(net318));
 sg13g2_xor2_1 _2359_ (.B(_1507_),
    .A(_1492_),
    .X(_1508_));
 sg13g2_xnor2_1 _2360_ (.Y(_1509_),
    .A(_1492_),
    .B(_1507_));
 sg13g2_o21ai_1 _2361_ (.B1(_1508_),
    .Y(_1510_),
    .A1(_1494_),
    .A2(_1505_));
 sg13g2_o21ai_1 _2362_ (.B1(_1510_),
    .Y(_1511_),
    .A1(\px[4] ),
    .A2(_1392_));
 sg13g2_a21oi_2 _2363_ (.B1(_1511_),
    .Y(_1512_),
    .A2(_1507_),
    .A1(_1492_));
 sg13g2_nand2_1 _2364_ (.Y(_1513_),
    .A(net352),
    .B(net317));
 sg13g2_xor2_1 _2365_ (.B(net317),
    .A(net352),
    .X(_1514_));
 sg13g2_o21ai_1 _2366_ (.B1(_1490_),
    .Y(_1515_),
    .A1(_1512_),
    .A2(_1514_));
 sg13g2_a221oi_1 _2367_ (.B2(_1515_),
    .C1(_1487_),
    .B1(_1488_),
    .A1(_1384_),
    .Y(_1516_),
    .A2(net312));
 sg13g2_a21oi_1 _2368_ (.A1(net350),
    .A2(_1391_),
    .Y(_1517_),
    .B1(_1516_));
 sg13g2_nor2b_2 _2369_ (.A(\px[9] ),
    .B_N(net311),
    .Y(_1518_));
 sg13g2_inv_1 _2370_ (.Y(_1519_),
    .A(_1518_));
 sg13g2_a21oi_1 _2371_ (.A1(_1485_),
    .A2(_1517_),
    .Y(_1520_),
    .B1(_1484_));
 sg13g2_a21oi_2 _2372_ (.B1(_1483_),
    .Y(_1521_),
    .A2(_1520_),
    .A1(_1519_));
 sg13g2_xor2_1 _2373_ (.B(_1517_),
    .A(_1486_),
    .X(_1522_));
 sg13g2_xor2_1 _2374_ (.B(_1515_),
    .A(_1489_),
    .X(_1523_));
 sg13g2_or3_2 _2375_ (.A(_1494_),
    .B(_1505_),
    .C(_1508_),
    .X(_1524_));
 sg13g2_or3_1 _2376_ (.A(_1494_),
    .B(_1505_),
    .C(_1509_),
    .X(_1525_));
 sg13g2_o21ai_1 _2377_ (.B1(_1509_),
    .Y(_1526_),
    .A1(_1494_),
    .A2(_1505_));
 sg13g2_nand2_2 _2378_ (.Y(_1527_),
    .A(_1525_),
    .B(_1526_));
 sg13g2_nand2_2 _2379_ (.Y(_1528_),
    .A(_1441_),
    .B(_1444_));
 sg13g2_nand2_1 _2380_ (.Y(_1529_),
    .A(net327),
    .B(_1528_));
 sg13g2_nor2_1 _2381_ (.A(_0023_),
    .B(_1529_),
    .Y(_1530_));
 sg13g2_xnor2_1 _2382_ (.Y(_1531_),
    .A(_0057_),
    .B(_1530_));
 sg13g2_nor2_1 _2383_ (.A(_0022_),
    .B(_1531_),
    .Y(_1532_));
 sg13g2_nand2_1 _2384_ (.Y(_1533_),
    .A(net334),
    .B(\py[3] ));
 sg13g2_xnor2_1 _2385_ (.Y(_1534_),
    .A(net334),
    .B(net345));
 sg13g2_nand2_1 _2386_ (.Y(_1535_),
    .A(net336),
    .B(\py[2] ));
 sg13g2_xor2_1 _2387_ (.B(\py[2] ),
    .A(net336),
    .X(_1536_));
 sg13g2_nand2_1 _2388_ (.Y(_1537_),
    .A(net339),
    .B(\py[1] ));
 sg13g2_nand2_1 _2389_ (.Y(_1538_),
    .A(net341),
    .B(net347));
 sg13g2_nor2_1 _2390_ (.A(net338),
    .B(net346),
    .Y(_1539_));
 sg13g2_xor2_1 _2391_ (.B(net346),
    .A(net338),
    .X(_1540_));
 sg13g2_o21ai_1 _2392_ (.B1(_1537_),
    .Y(_1541_),
    .A1(_1538_),
    .A2(_1539_));
 sg13g2_nand2_1 _2393_ (.Y(_1542_),
    .A(_1536_),
    .B(_1541_));
 sg13g2_or2_1 _2394_ (.X(_1543_),
    .B(_1535_),
    .A(_1534_));
 sg13g2_xnor2_1 _2395_ (.Y(_1544_),
    .A(_1534_),
    .B(_1535_));
 sg13g2_nand3b_1 _2396_ (.B(_1536_),
    .C(_1541_),
    .Y(_1545_),
    .A_N(_1534_));
 sg13g2_xor2_1 _2397_ (.B(_1544_),
    .A(_1542_),
    .X(_1546_));
 sg13g2_xnor2_1 _2398_ (.Y(_1547_),
    .A(_1542_),
    .B(_1544_));
 sg13g2_xnor2_1 _2399_ (.Y(_1548_),
    .A(\px[0] ),
    .B(net322));
 sg13g2_xor2_1 _2400_ (.B(net322),
    .A(\px[0] ),
    .X(_1549_));
 sg13g2_xnor2_1 _2401_ (.Y(_1550_),
    .A(_1499_),
    .B(_1500_));
 sg13g2_inv_1 _2402_ (.Y(_1551_),
    .A(_1550_));
 sg13g2_nand2_2 _2403_ (.Y(_1552_),
    .A(net308),
    .B(_1550_));
 sg13g2_nor2_1 _2404_ (.A(_1499_),
    .B(net308),
    .Y(_1553_));
 sg13g2_a21oi_1 _2405_ (.A1(net308),
    .A2(_1550_),
    .Y(_1554_),
    .B1(_1553_));
 sg13g2_o21ai_1 _2406_ (.B1(_1552_),
    .Y(_1555_),
    .A1(_1499_),
    .A2(net308));
 sg13g2_xor2_1 _2407_ (.B(net347),
    .A(net340),
    .X(_1556_));
 sg13g2_xnor2_1 _2408_ (.Y(_1557_),
    .A(net340),
    .B(net347));
 sg13g2_xnor2_1 _2409_ (.Y(_1558_),
    .A(_1538_),
    .B(_1540_));
 sg13g2_inv_2 _2410_ (.Y(_1559_),
    .A(_1558_));
 sg13g2_nand2_2 _2411_ (.Y(_1560_),
    .A(_1540_),
    .B(net307));
 sg13g2_o21ai_1 _2412_ (.B1(_1560_),
    .Y(_1561_),
    .A1(net307),
    .A2(_1558_));
 sg13g2_xnor2_1 _2413_ (.Y(_1562_),
    .A(_1536_),
    .B(_1541_));
 sg13g2_xor2_1 _2414_ (.B(\py[4] ),
    .A(net332),
    .X(_1563_));
 sg13g2_xnor2_1 _2415_ (.Y(_1564_),
    .A(_1533_),
    .B(_1563_));
 sg13g2_xnor2_1 _2416_ (.Y(_1565_),
    .A(_1506_),
    .B(_1514_));
 sg13g2_or2_1 _2417_ (.X(_1566_),
    .B(_1518_),
    .A(_1483_));
 sg13g2_nor2_1 _2418_ (.A(_1485_),
    .B(_1566_),
    .Y(_1567_));
 sg13g2_nor4_1 _2419_ (.A(net323),
    .B(_1564_),
    .C(_1565_),
    .D(_1567_),
    .Y(_1568_));
 sg13g2_xor2_1 _2420_ (.B(net312),
    .A(net350),
    .X(_1569_));
 sg13g2_a22oi_1 _2421_ (.Y(_1570_),
    .B1(_1569_),
    .B2(_1488_),
    .A2(_1566_),
    .A1(_1485_));
 sg13g2_o21ai_1 _2422_ (.B1(_1570_),
    .Y(_1571_),
    .A1(_1488_),
    .A2(_1569_));
 sg13g2_a21oi_1 _2423_ (.A1(_1429_),
    .A2(_1528_),
    .Y(_1572_),
    .B1(_1571_));
 sg13g2_nand3_1 _2424_ (.B(_1568_),
    .C(_1572_),
    .A(_1562_),
    .Y(_1573_));
 sg13g2_a21o_1 _2425_ (.A2(_1561_),
    .A1(_1555_),
    .B1(_1573_),
    .X(_1574_));
 sg13g2_nor4_1 _2426_ (.A(_1527_),
    .B(_1532_),
    .C(_1547_),
    .D(_1574_),
    .Y(_1575_));
 sg13g2_nand2_1 _2427_ (.Y(_1576_),
    .A(_0026_),
    .B(_1445_));
 sg13g2_xnor2_1 _2428_ (.Y(_1577_),
    .A(_0026_),
    .B(_1445_));
 sg13g2_nor2b_1 _2429_ (.A(_0061_),
    .B_N(_1577_),
    .Y(_1578_));
 sg13g2_xor2_1 _2430_ (.B(_1576_),
    .A(net330),
    .X(_1579_));
 sg13g2_xnor2_1 _2431_ (.Y(_1580_),
    .A(\py[5] ),
    .B(_1579_));
 sg13g2_nor2_1 _2432_ (.A(_1578_),
    .B(_1580_),
    .Y(_1581_));
 sg13g2_xnor2_1 _2433_ (.Y(_1582_),
    .A(_1578_),
    .B(_1580_));
 sg13g2_xnor2_1 _2434_ (.Y(_1583_),
    .A(_1383_),
    .B(_1577_));
 sg13g2_xnor2_1 _2435_ (.Y(_1584_),
    .A(net334),
    .B(_1444_));
 sg13g2_xnor2_1 _2436_ (.Y(_1585_),
    .A(net336),
    .B(_1443_));
 sg13g2_nor2_1 _2437_ (.A(_0062_),
    .B(_1585_),
    .Y(_1586_));
 sg13g2_nand2_1 _2438_ (.Y(_1587_),
    .A(_1374_),
    .B(net348));
 sg13g2_nand3_1 _2439_ (.B(_1374_),
    .C(net347),
    .A(_1373_),
    .Y(_1588_));
 sg13g2_a22oi_1 _2440_ (.Y(_1589_),
    .B1(_1588_),
    .B2(_0063_),
    .A2(_1587_),
    .A1(_1427_));
 sg13g2_a22oi_1 _2441_ (.Y(_1590_),
    .B1(_1585_),
    .B2(_0062_),
    .A2(_1584_),
    .A1(_0027_));
 sg13g2_o21ai_1 _2442_ (.B1(_1590_),
    .Y(_1591_),
    .A1(_1586_),
    .A2(_1589_));
 sg13g2_o21ai_1 _2443_ (.B1(_1591_),
    .Y(_1592_),
    .A1(_0027_),
    .A2(_1584_));
 sg13g2_nor3_1 _2444_ (.A(_1582_),
    .B(_1583_),
    .C(_1592_),
    .Y(_1593_));
 sg13g2_and3_1 _2445_ (.X(_1594_),
    .A(_1582_),
    .B(_1583_),
    .C(_1592_));
 sg13g2_xor2_1 _2446_ (.B(_1529_),
    .A(net326),
    .X(_1595_));
 sg13g2_nor2_1 _2447_ (.A(_0024_),
    .B(_1595_),
    .Y(_1596_));
 sg13g2_xnor2_1 _2448_ (.Y(_1597_),
    .A(\py[9] ),
    .B(_1531_));
 sg13g2_nand2_1 _2449_ (.Y(_1598_),
    .A(_1596_),
    .B(_1597_));
 sg13g2_nand3_1 _2450_ (.B(_1503_),
    .C(_1504_),
    .A(_1497_),
    .Y(_1599_));
 sg13g2_nand2b_1 _2451_ (.Y(_1600_),
    .B(_1599_),
    .A_N(_1505_));
 sg13g2_xor2_1 _2452_ (.B(_1502_),
    .A(_1501_),
    .X(_1601_));
 sg13g2_inv_1 _2453_ (.Y(_1602_),
    .A(_1601_));
 sg13g2_a21oi_1 _2454_ (.A1(_1510_),
    .A2(_1524_),
    .Y(_1603_),
    .B1(_1601_));
 sg13g2_nor2b_1 _2455_ (.A(net304),
    .B_N(_1603_),
    .Y(_1604_));
 sg13g2_nor2_1 _2456_ (.A(_0060_),
    .B(_1579_),
    .Y(_1605_));
 sg13g2_a21oi_2 _2457_ (.B1(_1370_),
    .Y(_1606_),
    .A2(_1439_),
    .A1(_1372_));
 sg13g2_o21ai_1 _2458_ (.B1(_1528_),
    .Y(_1607_),
    .A1(_1370_),
    .A2(_1444_));
 sg13g2_nor2_2 _2459_ (.A(_1606_),
    .B(_1607_),
    .Y(_1608_));
 sg13g2_xnor2_1 _2460_ (.Y(_1609_),
    .A(\py[6] ),
    .B(_1608_));
 sg13g2_nand2_1 _2461_ (.Y(_1610_),
    .A(_1605_),
    .B(_1609_));
 sg13g2_nor2_1 _2462_ (.A(_0059_),
    .B(_1608_),
    .Y(_1611_));
 sg13g2_xor2_1 _2463_ (.B(_1528_),
    .A(_0025_),
    .X(_1612_));
 sg13g2_xnor2_1 _2464_ (.Y(_1613_),
    .A(\py[7] ),
    .B(_1612_));
 sg13g2_nand2_1 _2465_ (.Y(_1614_),
    .A(_1611_),
    .B(_1613_));
 sg13g2_xor2_1 _2466_ (.B(_1613_),
    .A(_1611_),
    .X(_1615_));
 sg13g2_xnor2_1 _2467_ (.Y(_1616_),
    .A(_1610_),
    .B(_1615_));
 sg13g2_or2_1 _2468_ (.X(_1617_),
    .B(_1609_),
    .A(_1605_));
 sg13g2_nand2_1 _2469_ (.Y(_1618_),
    .A(_1610_),
    .B(_1617_));
 sg13g2_nor2_1 _2470_ (.A(_1581_),
    .B(_1593_),
    .Y(_1619_));
 sg13g2_nor2_1 _2471_ (.A(_1618_),
    .B(_1619_),
    .Y(_1620_));
 sg13g2_xnor2_1 _2472_ (.Y(_1621_),
    .A(_1618_),
    .B(_1619_));
 sg13g2_xor2_1 _2473_ (.B(_1595_),
    .A(\py[8] ),
    .X(_1622_));
 sg13g2_or3_1 _2474_ (.A(_0064_),
    .B(_1612_),
    .C(_1622_),
    .X(_1623_));
 sg13g2_or3_1 _2475_ (.A(_1596_),
    .B(_1597_),
    .C(_1623_),
    .X(_1624_));
 sg13g2_o21ai_1 _2476_ (.B1(_1623_),
    .Y(_1625_),
    .A1(_1596_),
    .A2(_1597_));
 sg13g2_and2_1 _2477_ (.A(_1624_),
    .B(_1625_),
    .X(_1626_));
 sg13g2_o21ai_1 _2478_ (.B1(_1617_),
    .Y(_1627_),
    .A1(_1611_),
    .A2(_1613_));
 sg13g2_o21ai_1 _2479_ (.B1(_1614_),
    .Y(_1628_),
    .A1(_1620_),
    .A2(_1627_));
 sg13g2_o21ai_1 _2480_ (.B1(_1622_),
    .Y(_1629_),
    .A1(_0064_),
    .A2(_1612_));
 sg13g2_a21oi_1 _2481_ (.A1(_1623_),
    .A2(_1629_),
    .Y(_1630_),
    .B1(_1628_));
 sg13g2_nand3_1 _2482_ (.B(_1628_),
    .C(_1629_),
    .A(_1624_),
    .Y(_1631_));
 sg13g2_o21ai_1 _2483_ (.B1(_1604_),
    .Y(_1632_),
    .A1(_1593_),
    .A2(_1594_));
 sg13g2_nand3_1 _2484_ (.B(_1598_),
    .C(_1616_),
    .A(_1575_),
    .Y(_1633_));
 sg13g2_nor4_1 _2485_ (.A(_1523_),
    .B(_1626_),
    .C(_1632_),
    .D(_1633_),
    .Y(_1634_));
 sg13g2_nand3_1 _2486_ (.B(_1631_),
    .C(_1634_),
    .A(_1621_),
    .Y(_1635_));
 sg13g2_nor3_1 _2487_ (.A(_1522_),
    .B(_1630_),
    .C(_1635_),
    .Y(_1636_));
 sg13g2_and2_2 _2488_ (.A(_1521_),
    .B(_1636_),
    .X(_1637_));
 sg13g2_nand2b_1 _2489_ (.Y(_1638_),
    .B(_1481_),
    .A_N(_1637_));
 sg13g2_nor2_2 _2490_ (.A(net323),
    .B(_1429_),
    .Y(_1639_));
 sg13g2_nand2_2 _2491_ (.Y(_1640_),
    .A(_1368_),
    .B(_1430_));
 sg13g2_nand2_1 _2492_ (.Y(_1641_),
    .A(_1502_),
    .B(_1550_));
 sg13g2_a21oi_2 _2493_ (.B1(net308),
    .Y(_1642_),
    .A2(_1524_),
    .A1(_1510_));
 sg13g2_a21oi_2 _2494_ (.B1(_1564_),
    .Y(_1643_),
    .A2(_1545_),
    .A1(_1543_));
 sg13g2_and3_1 _2495_ (.X(_1644_),
    .A(_1543_),
    .B(_1545_),
    .C(_1564_));
 sg13g2_or2_2 _2496_ (.X(_1645_),
    .B(_1644_),
    .A(_1643_));
 sg13g2_nor2_2 _2497_ (.A(_1643_),
    .B(_1644_),
    .Y(_1646_));
 sg13g2_xnor2_1 _2498_ (.Y(_1647_),
    .A(_1641_),
    .B(_1646_));
 sg13g2_xnor2_1 _2499_ (.Y(_1648_),
    .A(_1642_),
    .B(_1647_));
 sg13g2_o21ai_1 _2500_ (.B1(_1641_),
    .Y(_1649_),
    .A1(_1602_),
    .A2(_1648_));
 sg13g2_a21oi_2 _2501_ (.B1(_1527_),
    .Y(_1650_),
    .A2(_1645_),
    .A1(_1548_));
 sg13g2_nor2_1 _2502_ (.A(net304),
    .B(_1602_),
    .Y(_1651_));
 sg13g2_nand2b_2 _2503_ (.Y(_1652_),
    .B(_1601_),
    .A_N(net304));
 sg13g2_a21oi_1 _2504_ (.A1(_1510_),
    .A2(_1524_),
    .Y(_1653_),
    .B1(_1555_));
 sg13g2_xnor2_1 _2505_ (.Y(_1654_),
    .A(_1652_),
    .B(_1653_));
 sg13g2_and2_1 _2506_ (.A(_1650_),
    .B(_1654_),
    .X(_1655_));
 sg13g2_or2_1 _2507_ (.X(_1656_),
    .B(_1654_),
    .A(_1650_));
 sg13g2_xnor2_1 _2508_ (.Y(_1657_),
    .A(_1650_),
    .B(_1654_));
 sg13g2_nor3_2 _2509_ (.A(_1557_),
    .B(_1643_),
    .C(_1644_),
    .Y(_1658_));
 sg13g2_nand2_2 _2510_ (.Y(_1659_),
    .A(net307),
    .B(_1646_));
 sg13g2_a21oi_1 _2511_ (.A1(_1510_),
    .A2(_1524_),
    .Y(_1660_),
    .B1(_1550_));
 sg13g2_and2_1 _2512_ (.A(_1651_),
    .B(_1660_),
    .X(_1661_));
 sg13g2_xnor2_1 _2513_ (.Y(_1662_),
    .A(_1652_),
    .B(_1660_));
 sg13g2_xnor2_1 _2514_ (.Y(_1663_),
    .A(_1659_),
    .B(_1662_));
 sg13g2_xnor2_1 _2515_ (.Y(_1664_),
    .A(_1657_),
    .B(_1663_));
 sg13g2_nand2_1 _2516_ (.Y(_1665_),
    .A(_1649_),
    .B(_1664_));
 sg13g2_xnor2_1 _2517_ (.Y(_1666_),
    .A(_1649_),
    .B(_1664_));
 sg13g2_nand2b_2 _2518_ (.Y(_1667_),
    .B(_1658_),
    .A_N(_1527_));
 sg13g2_nor2_2 _2519_ (.A(_1547_),
    .B(_1559_),
    .Y(_1668_));
 sg13g2_xor2_1 _2520_ (.B(_1658_),
    .A(_1642_),
    .X(_1669_));
 sg13g2_nand2_1 _2521_ (.Y(_1670_),
    .A(_1668_),
    .B(_1669_));
 sg13g2_o21ai_1 _2522_ (.B1(_1670_),
    .Y(_1671_),
    .A1(net308),
    .A2(_1667_));
 sg13g2_nor2_1 _2523_ (.A(_1551_),
    .B(_1600_),
    .Y(_1672_));
 sg13g2_nand3_1 _2524_ (.B(_1646_),
    .C(_1672_),
    .A(_1558_),
    .Y(_1673_));
 sg13g2_a21o_1 _2525_ (.A2(_1646_),
    .A1(_1558_),
    .B1(_1672_),
    .X(_1674_));
 sg13g2_and2_1 _2526_ (.A(_1673_),
    .B(_1674_),
    .X(_1675_));
 sg13g2_nand2_1 _2527_ (.Y(_1676_),
    .A(_1671_),
    .B(_1675_));
 sg13g2_xnor2_1 _2528_ (.Y(_1677_),
    .A(_1671_),
    .B(_1675_));
 sg13g2_o21ai_1 _2529_ (.B1(_1665_),
    .Y(_1678_),
    .A1(_1666_),
    .A2(_1677_));
 sg13g2_a21oi_1 _2530_ (.A1(_1656_),
    .A2(_1663_),
    .Y(_1679_),
    .B1(_1655_));
 sg13g2_xnor2_1 _2531_ (.Y(_1680_),
    .A(net304),
    .B(_1603_));
 sg13g2_xnor2_1 _2532_ (.Y(_1681_),
    .A(_1659_),
    .B(_1680_));
 sg13g2_a21oi_1 _2533_ (.A1(_1510_),
    .A2(_1524_),
    .Y(_1682_),
    .B1(_1552_));
 sg13g2_and2_2 _2534_ (.A(_1601_),
    .B(_1682_),
    .X(_1683_));
 sg13g2_a22oi_1 _2535_ (.Y(_1684_),
    .B1(_1555_),
    .B2(_1602_),
    .A2(_1524_),
    .A1(_1510_));
 sg13g2_nand4_1 _2536_ (.B(_1526_),
    .C(_1554_),
    .A(_1525_),
    .Y(_1685_),
    .D(_1601_));
 sg13g2_a221oi_1 _2537_ (.B2(_1685_),
    .C1(_1682_),
    .B1(_1684_),
    .A1(_1651_),
    .Y(_1686_),
    .A2(_1653_));
 sg13g2_nor2_1 _2538_ (.A(_1683_),
    .B(_1686_),
    .Y(_1687_));
 sg13g2_xor2_1 _2539_ (.B(_1687_),
    .A(_1681_),
    .X(_1688_));
 sg13g2_nor2b_1 _2540_ (.A(_1679_),
    .B_N(_1688_),
    .Y(_1689_));
 sg13g2_xnor2_1 _2541_ (.Y(_1690_),
    .A(_1679_),
    .B(_1688_));
 sg13g2_nor2_1 _2542_ (.A(_1544_),
    .B(_1562_),
    .Y(_1691_));
 sg13g2_a21o_1 _2543_ (.A2(_1662_),
    .A1(_1658_),
    .B1(_1661_),
    .X(_1692_));
 sg13g2_nor2_2 _2544_ (.A(_1559_),
    .B(_1562_),
    .Y(_1693_));
 sg13g2_and2_1 _2545_ (.A(_1559_),
    .B(_1562_),
    .X(_1694_));
 sg13g2_nor2_1 _2546_ (.A(_1693_),
    .B(_1694_),
    .Y(_1695_));
 sg13g2_and2_1 _2547_ (.A(_1646_),
    .B(_1695_),
    .X(_1696_));
 sg13g2_xnor2_1 _2548_ (.Y(_1697_),
    .A(net305),
    .B(_1696_));
 sg13g2_nor2b_1 _2549_ (.A(_1697_),
    .B_N(_1692_),
    .Y(_1698_));
 sg13g2_xnor2_1 _2550_ (.Y(_1699_),
    .A(_1692_),
    .B(_1697_));
 sg13g2_xor2_1 _2551_ (.B(_1699_),
    .A(_1691_),
    .X(_1700_));
 sg13g2_xor2_1 _2552_ (.B(_1700_),
    .A(_1690_),
    .X(_1701_));
 sg13g2_and2_1 _2553_ (.A(_1678_),
    .B(_1701_),
    .X(_1702_));
 sg13g2_nand2_1 _2554_ (.Y(_1703_),
    .A(_1562_),
    .B(_1646_));
 sg13g2_a21oi_2 _2555_ (.B1(_1703_),
    .Y(_1704_),
    .A2(_1676_),
    .A1(_1673_));
 sg13g2_nand3_1 _2556_ (.B(_1676_),
    .C(_1703_),
    .A(_1673_),
    .Y(_1705_));
 sg13g2_nor2b_1 _2557_ (.A(_1704_),
    .B_N(_1705_),
    .Y(_1706_));
 sg13g2_or2_1 _2558_ (.X(_1707_),
    .B(_1701_),
    .A(_1678_));
 sg13g2_xnor2_1 _2559_ (.Y(_1708_),
    .A(_1678_),
    .B(_1701_));
 sg13g2_a21oi_1 _2560_ (.A1(_1706_),
    .A2(_1707_),
    .Y(_1709_),
    .B1(_1702_));
 sg13g2_a21oi_1 _2561_ (.A1(_1691_),
    .A2(_1699_),
    .Y(_1710_),
    .B1(_1698_));
 sg13g2_nand2_1 _2562_ (.Y(_1711_),
    .A(_1547_),
    .B(_1646_));
 sg13g2_nor2_1 _2563_ (.A(_1710_),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_xor2_1 _2564_ (.B(_1711_),
    .A(_1710_),
    .X(_1713_));
 sg13g2_a21oi_1 _2565_ (.A1(_1690_),
    .A2(_1700_),
    .Y(_1714_),
    .B1(_1689_));
 sg13g2_a21oi_1 _2566_ (.A1(_1681_),
    .A2(_1687_),
    .Y(_1715_),
    .B1(_1683_));
 sg13g2_nor2_1 _2567_ (.A(_1682_),
    .B(_1684_),
    .Y(_1716_));
 sg13g2_nor2_2 _2568_ (.A(_1683_),
    .B(_1716_),
    .Y(_1717_));
 sg13g2_xnor2_1 _2569_ (.Y(_1718_),
    .A(_1527_),
    .B(_1658_));
 sg13g2_xnor2_1 _2570_ (.Y(_1719_),
    .A(_1717_),
    .B(_1718_));
 sg13g2_nor2_1 _2571_ (.A(_1715_),
    .B(_1719_),
    .Y(_1720_));
 sg13g2_xnor2_1 _2572_ (.Y(_1721_),
    .A(_1715_),
    .B(_1719_));
 sg13g2_nor2_1 _2573_ (.A(net305),
    .B(_1693_),
    .Y(_1722_));
 sg13g2_nor3_2 _2574_ (.A(_1645_),
    .B(_1694_),
    .C(_1722_),
    .Y(_1723_));
 sg13g2_nor2_1 _2575_ (.A(_1645_),
    .B(_1695_),
    .Y(_1724_));
 sg13g2_mux2_2 _2576_ (.A0(_1696_),
    .A1(_1724_),
    .S(net305),
    .X(_1725_));
 sg13g2_a21oi_1 _2577_ (.A1(_1658_),
    .A2(_1680_),
    .Y(_1726_),
    .B1(_1604_));
 sg13g2_nor2b_1 _2578_ (.A(_1726_),
    .B_N(_1725_),
    .Y(_1727_));
 sg13g2_xnor2_1 _2579_ (.Y(_1728_),
    .A(_1725_),
    .B(_1726_));
 sg13g2_xnor2_1 _2580_ (.Y(_1729_),
    .A(_1723_),
    .B(_1728_));
 sg13g2_nor2_1 _2581_ (.A(_1721_),
    .B(_1729_),
    .Y(_1730_));
 sg13g2_xnor2_1 _2582_ (.Y(_1731_),
    .A(_1721_),
    .B(_1729_));
 sg13g2_nor2_1 _2583_ (.A(_1714_),
    .B(_1731_),
    .Y(_1732_));
 sg13g2_xor2_1 _2584_ (.B(_1731_),
    .A(_1714_),
    .X(_1733_));
 sg13g2_xnor2_1 _2585_ (.Y(_1734_),
    .A(_1713_),
    .B(_1733_));
 sg13g2_nor2_1 _2586_ (.A(_1709_),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_xor2_1 _2587_ (.B(_1734_),
    .A(_1709_),
    .X(_1736_));
 sg13g2_a21oi_2 _2588_ (.B1(_1735_),
    .Y(_1737_),
    .A2(_1736_),
    .A1(_1704_));
 sg13g2_a21oi_1 _2589_ (.A1(_1713_),
    .A2(_1733_),
    .Y(_1738_),
    .B1(_1732_));
 sg13g2_a21oi_1 _2590_ (.A1(_1723_),
    .A2(_1728_),
    .Y(_1739_),
    .B1(_1727_));
 sg13g2_inv_1 _2591_ (.Y(_1740_),
    .A(_1739_));
 sg13g2_nor2_1 _2592_ (.A(_1720_),
    .B(_1730_),
    .Y(_1741_));
 sg13g2_or2_1 _2593_ (.X(_1742_),
    .B(_1667_),
    .A(net304));
 sg13g2_o21ai_1 _2594_ (.B1(_1659_),
    .Y(_1743_),
    .A1(_1527_),
    .A2(net304));
 sg13g2_nand2_1 _2595_ (.Y(_1744_),
    .A(_1742_),
    .B(_1743_));
 sg13g2_a21oi_1 _2596_ (.A1(_1742_),
    .A2(_1743_),
    .Y(_1745_),
    .B1(_1717_));
 sg13g2_xor2_1 _2597_ (.B(_1744_),
    .A(_1717_),
    .X(_1746_));
 sg13g2_a21oi_1 _2598_ (.A1(_1717_),
    .A2(_1718_),
    .Y(_1747_),
    .B1(_1683_));
 sg13g2_or2_1 _2599_ (.X(_1748_),
    .B(_1747_),
    .A(_1746_));
 sg13g2_xnor2_1 _2600_ (.Y(_1749_),
    .A(_1746_),
    .B(_1747_));
 sg13g2_nor2b_1 _2601_ (.A(_1667_),
    .B_N(_1725_),
    .Y(_1750_));
 sg13g2_xnor2_1 _2602_ (.Y(_1751_),
    .A(_1667_),
    .B(_1725_));
 sg13g2_xnor2_1 _2603_ (.Y(_1752_),
    .A(_1723_),
    .B(_1751_));
 sg13g2_xor2_1 _2604_ (.B(_1752_),
    .A(_1749_),
    .X(_1753_));
 sg13g2_nor2b_1 _2605_ (.A(_1741_),
    .B_N(_1753_),
    .Y(_1754_));
 sg13g2_xnor2_1 _2606_ (.Y(_1755_),
    .A(_1741_),
    .B(_1753_));
 sg13g2_xnor2_1 _2607_ (.Y(_1756_),
    .A(_1739_),
    .B(_1755_));
 sg13g2_nor2b_1 _2608_ (.A(_1738_),
    .B_N(_1756_),
    .Y(_1757_));
 sg13g2_xnor2_1 _2609_ (.Y(_1758_),
    .A(_1738_),
    .B(_1756_));
 sg13g2_xor2_1 _2610_ (.B(_1758_),
    .A(_1712_),
    .X(_1759_));
 sg13g2_nand2b_1 _2611_ (.Y(_1760_),
    .B(_1759_),
    .A_N(_1737_));
 sg13g2_nor2b_1 _2612_ (.A(_1759_),
    .B_N(_1737_),
    .Y(_1761_));
 sg13g2_xnor2_1 _2613_ (.Y(_1762_),
    .A(_1737_),
    .B(_1759_));
 sg13g2_nand2_1 _2614_ (.Y(_1763_),
    .A(net304),
    .B(_1602_));
 sg13g2_nand3_1 _2615_ (.B(_1652_),
    .C(_1763_),
    .A(net308),
    .Y(_1764_));
 sg13g2_nor2_1 _2616_ (.A(_1548_),
    .B(net304),
    .Y(_1765_));
 sg13g2_nand2_1 _2617_ (.Y(_1766_),
    .A(net305),
    .B(net307));
 sg13g2_nand3_1 _2618_ (.B(net307),
    .C(_1765_),
    .A(net305),
    .Y(_1767_));
 sg13g2_xnor2_1 _2619_ (.Y(_1768_),
    .A(_1765_),
    .B(_1766_));
 sg13g2_nand2b_1 _2620_ (.Y(_1769_),
    .B(_1768_),
    .A_N(_1764_));
 sg13g2_o21ai_1 _2621_ (.B1(_1769_),
    .Y(_1770_),
    .A1(_1548_),
    .A2(_1652_));
 sg13g2_xnor2_1 _2622_ (.Y(_1771_),
    .A(_1601_),
    .B(_1648_));
 sg13g2_and2_1 _2623_ (.A(_1770_),
    .B(_1771_),
    .X(_1772_));
 sg13g2_or2_1 _2624_ (.X(_1773_),
    .B(_1771_),
    .A(_1770_));
 sg13g2_xnor2_1 _2625_ (.Y(_1774_),
    .A(_1770_),
    .B(_1771_));
 sg13g2_xnor2_1 _2626_ (.Y(_1775_),
    .A(_1668_),
    .B(_1669_));
 sg13g2_nor2_1 _2627_ (.A(_1767_),
    .B(_1775_),
    .Y(_1776_));
 sg13g2_xor2_1 _2628_ (.B(_1775_),
    .A(_1767_),
    .X(_1777_));
 sg13g2_xor2_1 _2629_ (.B(_1777_),
    .A(_1693_),
    .X(_1778_));
 sg13g2_a21oi_1 _2630_ (.A1(_1773_),
    .A2(_1778_),
    .Y(_1779_),
    .B1(_1772_));
 sg13g2_xor2_1 _2631_ (.B(_1677_),
    .A(_1666_),
    .X(_1780_));
 sg13g2_nand2b_1 _2632_ (.Y(_1781_),
    .B(_1780_),
    .A_N(_1779_));
 sg13g2_xor2_1 _2633_ (.B(_1780_),
    .A(_1779_),
    .X(_1782_));
 sg13g2_nor2_1 _2634_ (.A(net307),
    .B(_1645_),
    .Y(_1783_));
 sg13g2_xnor2_1 _2635_ (.Y(_1784_),
    .A(_1562_),
    .B(_1668_));
 sg13g2_a22oi_1 _2636_ (.Y(_1785_),
    .B1(_1783_),
    .B2(_1784_),
    .A2(_1693_),
    .A1(_1546_));
 sg13g2_inv_1 _2637_ (.Y(_1786_),
    .A(_1785_));
 sg13g2_nor4_1 _2638_ (.A(_1558_),
    .B(_1645_),
    .C(_1767_),
    .D(_1775_),
    .Y(_1787_));
 sg13g2_a221oi_1 _2639_ (.B2(_1777_),
    .C1(_1776_),
    .B1(_1693_),
    .A1(_1559_),
    .Y(_1788_),
    .A2(_1646_));
 sg13g2_nor2_1 _2640_ (.A(_1787_),
    .B(_1788_),
    .Y(_1789_));
 sg13g2_xnor2_1 _2641_ (.Y(_1790_),
    .A(_1786_),
    .B(_1789_));
 sg13g2_o21ai_1 _2642_ (.B1(_1781_),
    .Y(_1791_),
    .A1(_1782_),
    .A2(_1790_));
 sg13g2_xnor2_1 _2643_ (.Y(_1792_),
    .A(_1706_),
    .B(_1708_));
 sg13g2_nand2_1 _2644_ (.Y(_1793_),
    .A(_1791_),
    .B(_1792_));
 sg13g2_a21oi_1 _2645_ (.A1(_1786_),
    .A2(_1789_),
    .Y(_1794_),
    .B1(_1787_));
 sg13g2_nor2_1 _2646_ (.A(_1791_),
    .B(_1792_),
    .Y(_1795_));
 sg13g2_xor2_1 _2647_ (.B(_1792_),
    .A(_1791_),
    .X(_1796_));
 sg13g2_o21ai_1 _2648_ (.B1(_1793_),
    .Y(_1797_),
    .A1(_1794_),
    .A2(_1795_));
 sg13g2_xnor2_1 _2649_ (.Y(_1798_),
    .A(_1704_),
    .B(_1736_));
 sg13g2_nor2b_1 _2650_ (.A(_1798_),
    .B_N(_1797_),
    .Y(_1799_));
 sg13g2_xnor2_1 _2651_ (.Y(_1800_),
    .A(_1794_),
    .B(_1796_));
 sg13g2_nand2_1 _2652_ (.Y(_1801_),
    .A(_1499_),
    .B(_1548_));
 sg13g2_nor2_1 _2653_ (.A(_1557_),
    .B(_1562_),
    .Y(_1802_));
 sg13g2_nand2b_1 _2654_ (.Y(_1803_),
    .B(_1802_),
    .A_N(_1801_));
 sg13g2_nand2_1 _2655_ (.Y(_1804_),
    .A(_1552_),
    .B(_1803_));
 sg13g2_xnor2_1 _2656_ (.Y(_1805_),
    .A(_1764_),
    .B(_1768_));
 sg13g2_and2_1 _2657_ (.A(_1804_),
    .B(_1805_),
    .X(_1806_));
 sg13g2_o21ai_1 _2658_ (.B1(_1556_),
    .Y(_1807_),
    .A1(net305),
    .A2(_1693_));
 sg13g2_a21oi_1 _2659_ (.A1(net305),
    .A2(_1693_),
    .Y(_1808_),
    .B1(_1807_));
 sg13g2_xor2_1 _2660_ (.B(_1805_),
    .A(_1804_),
    .X(_1809_));
 sg13g2_a21oi_1 _2661_ (.A1(_1808_),
    .A2(_1809_),
    .Y(_1810_),
    .B1(_1806_));
 sg13g2_xnor2_1 _2662_ (.Y(_1811_),
    .A(_1774_),
    .B(_1778_));
 sg13g2_nor2b_1 _2663_ (.A(_1810_),
    .B_N(_1811_),
    .Y(_1812_));
 sg13g2_xor2_1 _2664_ (.B(_1784_),
    .A(_1783_),
    .X(_1813_));
 sg13g2_nor2_1 _2665_ (.A(_1560_),
    .B(_1562_),
    .Y(_1814_));
 sg13g2_a21oi_1 _2666_ (.A1(net305),
    .A2(_1814_),
    .Y(_1815_),
    .B1(_1813_));
 sg13g2_inv_1 _2667_ (.Y(_1816_),
    .A(_1815_));
 sg13g2_xnor2_1 _2668_ (.Y(_1817_),
    .A(_1810_),
    .B(_1811_));
 sg13g2_a21oi_1 _2669_ (.A1(_1816_),
    .A2(_1817_),
    .Y(_1818_),
    .B1(_1812_));
 sg13g2_xnor2_1 _2670_ (.Y(_1819_),
    .A(_1782_),
    .B(_1790_));
 sg13g2_or2_1 _2671_ (.X(_1820_),
    .B(_1819_),
    .A(_1818_));
 sg13g2_xnor2_1 _2672_ (.Y(_1821_),
    .A(_1815_),
    .B(_1817_));
 sg13g2_a221oi_1 _2673_ (.B2(_1540_),
    .C1(_1694_),
    .B1(_1802_),
    .A1(_1557_),
    .Y(_1822_),
    .A2(_1559_));
 sg13g2_xnor2_1 _2674_ (.Y(_1823_),
    .A(_1801_),
    .B(_1802_));
 sg13g2_and2_1 _2675_ (.A(_1822_),
    .B(_1823_),
    .X(_1824_));
 sg13g2_inv_1 _2676_ (.Y(_1825_),
    .A(_1824_));
 sg13g2_xnor2_1 _2677_ (.Y(_1826_),
    .A(_1808_),
    .B(_1809_));
 sg13g2_xnor2_1 _2678_ (.Y(_1827_),
    .A(_1822_),
    .B(_1823_));
 sg13g2_xnor2_1 _2679_ (.Y(_1828_),
    .A(_1825_),
    .B(_1826_));
 sg13g2_or3_1 _2680_ (.A(_1560_),
    .B(_1827_),
    .C(_1828_),
    .X(_1829_));
 sg13g2_o21ai_1 _2681_ (.B1(_1829_),
    .Y(_1830_),
    .A1(_1825_),
    .A2(_1826_));
 sg13g2_nand2_1 _2682_ (.Y(_1831_),
    .A(_1821_),
    .B(_1830_));
 sg13g2_xnor2_1 _2683_ (.Y(_1832_),
    .A(_1818_),
    .B(_1819_));
 sg13g2_o21ai_1 _2684_ (.B1(_1820_),
    .Y(_1833_),
    .A1(_1831_),
    .A2(_1832_));
 sg13g2_and2_1 _2685_ (.A(_1800_),
    .B(_1833_),
    .X(_1834_));
 sg13g2_nand2b_1 _2686_ (.Y(_1835_),
    .B(_1798_),
    .A_N(_1797_));
 sg13g2_xor2_1 _2687_ (.B(_1798_),
    .A(_1797_),
    .X(_1836_));
 sg13g2_a21oi_1 _2688_ (.A1(_1834_),
    .A2(_1835_),
    .Y(_1837_),
    .B1(_1799_));
 sg13g2_o21ai_1 _2689_ (.B1(_1760_),
    .Y(_1838_),
    .A1(_1761_),
    .A2(_1837_));
 sg13g2_a21oi_1 _2690_ (.A1(_1740_),
    .A2(_1755_),
    .Y(_1839_),
    .B1(_1754_));
 sg13g2_o21ai_1 _2691_ (.B1(_1748_),
    .Y(_1840_),
    .A1(_1749_),
    .A2(_1752_));
 sg13g2_nand2_1 _2692_ (.Y(_1841_),
    .A(_1683_),
    .B(_1744_));
 sg13g2_o21ai_1 _2693_ (.B1(_1841_),
    .Y(_1842_),
    .A1(_1683_),
    .A2(_1745_));
 sg13g2_a21oi_1 _2694_ (.A1(_1723_),
    .A2(_1751_),
    .Y(_1843_),
    .B1(_1750_));
 sg13g2_xor2_1 _2695_ (.B(_1742_),
    .A(_1725_),
    .X(_1844_));
 sg13g2_xnor2_1 _2696_ (.Y(_1845_),
    .A(_1723_),
    .B(_1844_));
 sg13g2_xnor2_1 _2697_ (.Y(_1846_),
    .A(_1843_),
    .B(_1845_));
 sg13g2_xnor2_1 _2698_ (.Y(_1847_),
    .A(_1842_),
    .B(_1846_));
 sg13g2_xnor2_1 _2699_ (.Y(_1848_),
    .A(_1840_),
    .B(_1847_));
 sg13g2_xnor2_1 _2700_ (.Y(_0255_),
    .A(_1839_),
    .B(_1848_));
 sg13g2_a21oi_1 _2701_ (.A1(_1712_),
    .A2(_1758_),
    .Y(_0256_),
    .B1(_1757_));
 sg13g2_nand2_2 _2702_ (.Y(_0257_),
    .A(_0255_),
    .B(_0256_));
 sg13g2_nand2_1 _2703_ (.Y(_0258_),
    .A(_1838_),
    .B(_0257_));
 sg13g2_nand3_1 _2704_ (.B(_1838_),
    .C(_0257_),
    .A(\product_comp[9] ),
    .Y(_0259_));
 sg13g2_a21o_1 _2705_ (.A2(_0257_),
    .A1(_1838_),
    .B1(\product_comp[9] ),
    .X(_0260_));
 sg13g2_nand2_1 _2706_ (.Y(_0261_),
    .A(_0259_),
    .B(_0260_));
 sg13g2_xnor2_1 _2707_ (.Y(_0262_),
    .A(_1762_),
    .B(_1837_));
 sg13g2_xnor2_1 _2708_ (.Y(_0263_),
    .A(_0034_),
    .B(_0262_));
 sg13g2_a21oi_1 _2709_ (.A1(_0259_),
    .A2(_0260_),
    .Y(_0264_),
    .B1(_0263_));
 sg13g2_xnor2_1 _2710_ (.Y(_0265_),
    .A(_1834_),
    .B(_1836_));
 sg13g2_nand2b_1 _2711_ (.Y(_0266_),
    .B(_0265_),
    .A_N(net344));
 sg13g2_nand2b_1 _2712_ (.Y(_0267_),
    .B(net344),
    .A_N(_0265_));
 sg13g2_xor2_1 _2713_ (.B(_1833_),
    .A(_1800_),
    .X(_0268_));
 sg13g2_xnor2_1 _2714_ (.Y(_0269_),
    .A(_0035_),
    .B(_0268_));
 sg13g2_xor2_1 _2715_ (.B(_1832_),
    .A(_1831_),
    .X(_0270_));
 sg13g2_inv_1 _2716_ (.Y(_0271_),
    .A(_0270_));
 sg13g2_xor2_1 _2717_ (.B(_0270_),
    .A(_0036_),
    .X(_0272_));
 sg13g2_xor2_1 _2718_ (.B(_1830_),
    .A(_1821_),
    .X(_0273_));
 sg13g2_and2_1 _2719_ (.A(_0037_),
    .B(_0273_),
    .X(_0274_));
 sg13g2_nor2_1 _2720_ (.A(_0037_),
    .B(_0273_),
    .Y(_0275_));
 sg13g2_o21ai_1 _2721_ (.B1(_0272_),
    .Y(_0276_),
    .A1(_0037_),
    .A2(_0273_));
 sg13g2_nor3_1 _2722_ (.A(_0269_),
    .B(_0274_),
    .C(_0276_),
    .Y(_0277_));
 sg13g2_nand3_1 _2723_ (.B(_0267_),
    .C(_0277_),
    .A(_0266_),
    .Y(_0278_));
 sg13g2_o21ai_1 _2724_ (.B1(_1828_),
    .Y(_0279_),
    .A1(_1560_),
    .A2(_1827_));
 sg13g2_nand2_1 _2725_ (.Y(_0280_),
    .A(_1829_),
    .B(_0279_));
 sg13g2_nor2_1 _2726_ (.A(\product_comp[3] ),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_xnor2_1 _2727_ (.Y(_0282_),
    .A(_1560_),
    .B(_1827_));
 sg13g2_nor2_1 _2728_ (.A(_1548_),
    .B(_1557_),
    .Y(_0283_));
 sg13g2_nand2_1 _2729_ (.Y(_0284_),
    .A(_1549_),
    .B(net307));
 sg13g2_nor2_1 _2730_ (.A(net308),
    .B(net307),
    .Y(_0285_));
 sg13g2_o21ai_1 _2731_ (.B1(_0284_),
    .Y(_0286_),
    .A1(\product_comp[0] ),
    .A2(_0285_));
 sg13g2_nand2b_1 _2732_ (.Y(_0287_),
    .B(_0286_),
    .A_N(\product_comp[1] ));
 sg13g2_o21ai_1 _2733_ (.B1(_0287_),
    .Y(_0288_),
    .A1(\product_comp[2] ),
    .A2(_0282_));
 sg13g2_nor2_1 _2734_ (.A(_0281_),
    .B(_0288_),
    .Y(_0289_));
 sg13g2_a22oi_1 _2735_ (.Y(_0290_),
    .B1(_0282_),
    .B2(\product_comp[2] ),
    .A2(_0280_),
    .A1(\product_comp[3] ));
 sg13g2_a21oi_1 _2736_ (.A1(_0288_),
    .A2(_0290_),
    .Y(_0291_),
    .B1(_0281_));
 sg13g2_nand4_1 _2737_ (.B(_0267_),
    .C(_0277_),
    .A(_0266_),
    .Y(_0292_),
    .D(_0291_));
 sg13g2_nand2b_1 _2738_ (.Y(_0293_),
    .B(\product_comp[6] ),
    .A_N(_0268_));
 sg13g2_a22oi_1 _2739_ (.Y(_0294_),
    .B1(_0272_),
    .B2(_0275_),
    .A2(_0271_),
    .A1(\product_comp[5] ));
 sg13g2_o21ai_1 _2740_ (.B1(_0293_),
    .Y(_0295_),
    .A1(_0269_),
    .A2(_0294_));
 sg13g2_nand2_1 _2741_ (.Y(_0296_),
    .A(_0266_),
    .B(_0295_));
 sg13g2_nand3_1 _2742_ (.B(_0292_),
    .C(_0296_),
    .A(_0267_),
    .Y(_0297_));
 sg13g2_nor2b_1 _2743_ (.A(_0262_),
    .B_N(\product_comp[8] ),
    .Y(_0298_));
 sg13g2_a21oi_1 _2744_ (.A1(_1838_),
    .A2(_0257_),
    .Y(_0299_),
    .B1(_0033_));
 sg13g2_a221oi_1 _2745_ (.B2(_0261_),
    .C1(_0299_),
    .B1(_0298_),
    .A1(_0264_),
    .Y(_0300_),
    .A2(_0297_));
 sg13g2_o21ai_1 _2746_ (.B1(_1376_),
    .Y(_0301_),
    .A1(_1397_),
    .A2(_0300_));
 sg13g2_nor3_2 _2747_ (.A(\py[2] ),
    .B(\py[1] ),
    .C(net347),
    .Y(_0302_));
 sg13g2_nor2b_1 _2748_ (.A(net345),
    .B_N(_0302_),
    .Y(_0303_));
 sg13g2_and2_1 _2749_ (.A(_1383_),
    .B(_0303_),
    .X(_0304_));
 sg13g2_nor2b_1 _2750_ (.A(\py[5] ),
    .B_N(_0304_),
    .Y(_0305_));
 sg13g2_and2_1 _2751_ (.A(_1382_),
    .B(_0305_),
    .X(_0306_));
 sg13g2_nand2b_2 _2752_ (.Y(_0307_),
    .B(\py[7] ),
    .A_N(_0306_));
 sg13g2_inv_1 _2753_ (.Y(_0308_),
    .A(_0307_));
 sg13g2_xor2_1 _2754_ (.B(_0307_),
    .A(\py[8] ),
    .X(_0309_));
 sg13g2_xnor2_1 _2755_ (.Y(_0310_),
    .A(_0064_),
    .B(_0306_));
 sg13g2_xnor2_1 _2756_ (.Y(_0311_),
    .A(\py[6] ),
    .B(_0305_));
 sg13g2_xnor2_1 _2757_ (.Y(_0312_),
    .A(\py[5] ),
    .B(_0304_));
 sg13g2_inv_1 _2758_ (.Y(_0313_),
    .A(_0312_));
 sg13g2_nor2_1 _2759_ (.A(_0311_),
    .B(_0312_),
    .Y(_0314_));
 sg13g2_nor2b_2 _2760_ (.A(_0310_),
    .B_N(_0314_),
    .Y(_0315_));
 sg13g2_nand2b_2 _2761_ (.Y(_0316_),
    .B(_0315_),
    .A_N(_0309_));
 sg13g2_xor2_1 _2762_ (.B(_0315_),
    .A(_0309_),
    .X(_0317_));
 sg13g2_xnor2_1 _2763_ (.Y(_0318_),
    .A(\py[4] ),
    .B(_0303_));
 sg13g2_o21ai_1 _2764_ (.B1(\py[2] ),
    .Y(_0319_),
    .A1(net346),
    .A2(net347));
 sg13g2_nand2b_1 _2765_ (.Y(_0320_),
    .B(_0319_),
    .A_N(_0302_));
 sg13g2_xor2_1 _2766_ (.B(net347),
    .A(net346),
    .X(_0321_));
 sg13g2_a22oi_1 _2767_ (.Y(_0322_),
    .B1(_0031_),
    .B2(_0321_),
    .A2(net347),
    .A1(_1374_));
 sg13g2_o21ai_1 _2768_ (.B1(_0322_),
    .Y(_0323_),
    .A1(_0031_),
    .A2(_0321_));
 sg13g2_o21ai_1 _2769_ (.B1(_0323_),
    .Y(_0324_),
    .A1(_1373_),
    .A2(_0321_));
 sg13g2_xnor2_1 _2770_ (.Y(_0325_),
    .A(_0030_),
    .B(_0320_));
 sg13g2_a22oi_1 _2771_ (.Y(_0326_),
    .B1(_0324_),
    .B2(_0325_),
    .A2(_0320_),
    .A1(net336));
 sg13g2_xnor2_1 _2772_ (.Y(_0327_),
    .A(net345),
    .B(_0302_));
 sg13g2_xnor2_1 _2773_ (.Y(_0328_),
    .A(_1372_),
    .B(_0327_));
 sg13g2_nor2_1 _2774_ (.A(_0326_),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_nor2_1 _2775_ (.A(_0032_),
    .B(_0327_),
    .Y(_0330_));
 sg13g2_nor2_1 _2776_ (.A(_0026_),
    .B(_0318_),
    .Y(_0331_));
 sg13g2_nor3_1 _2777_ (.A(_0329_),
    .B(_0330_),
    .C(_0331_),
    .Y(_0332_));
 sg13g2_a21oi_2 _2778_ (.B1(_0332_),
    .Y(_0333_),
    .A2(_0318_),
    .A1(_0026_));
 sg13g2_xor2_1 _2779_ (.B(_0312_),
    .A(net330),
    .X(_0334_));
 sg13g2_a22oi_1 _2780_ (.Y(_0335_),
    .B1(_0333_),
    .B2(_0334_),
    .A2(_0312_),
    .A1(_1402_));
 sg13g2_a21oi_1 _2781_ (.A1(_1382_),
    .A2(_0312_),
    .Y(_0336_),
    .B1(_0314_));
 sg13g2_xor2_1 _2782_ (.B(_0336_),
    .A(_0029_),
    .X(_0337_));
 sg13g2_xnor2_1 _2783_ (.Y(_0338_),
    .A(_0310_),
    .B(_0314_));
 sg13g2_a22oi_1 _2784_ (.Y(_0339_),
    .B1(_0338_),
    .B2(net327),
    .A2(_0336_),
    .A1(net329));
 sg13g2_o21ai_1 _2785_ (.B1(_0339_),
    .Y(_0340_),
    .A1(_0335_),
    .A2(_0337_));
 sg13g2_nor2_1 _2786_ (.A(net327),
    .B(_0338_),
    .Y(_0341_));
 sg13g2_a21oi_1 _2787_ (.A1(_0023_),
    .A2(_0317_),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_nand2_1 _2788_ (.Y(_0343_),
    .A(_0340_),
    .B(_0342_));
 sg13g2_o21ai_1 _2789_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0023_),
    .A2(_0317_));
 sg13g2_nor2_1 _2790_ (.A(_0024_),
    .B(_0307_),
    .Y(_0345_));
 sg13g2_xnor2_1 _2791_ (.Y(_0346_),
    .A(_0022_),
    .B(_0345_));
 sg13g2_xor2_1 _2792_ (.B(_0346_),
    .A(_0057_),
    .X(_0347_));
 sg13g2_xnor2_1 _2793_ (.Y(_0348_),
    .A(_0316_),
    .B(_0347_));
 sg13g2_o21ai_1 _2794_ (.B1(net323),
    .Y(_0349_),
    .A1(_0316_),
    .A2(_0346_));
 sg13g2_a21oi_1 _2795_ (.A1(_0316_),
    .A2(_0346_),
    .Y(_0350_),
    .B1(_0349_));
 sg13g2_a21oi_1 _2796_ (.A1(_0344_),
    .A2(_0348_),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_nand2b_1 _2797_ (.Y(_0352_),
    .B(net329),
    .A_N(_0311_));
 sg13g2_xnor2_1 _2798_ (.Y(_0353_),
    .A(_1402_),
    .B(_0312_));
 sg13g2_a22oi_1 _2799_ (.Y(_0354_),
    .B1(_0333_),
    .B2(_0353_),
    .A2(_0313_),
    .A1(net330));
 sg13g2_xor2_1 _2800_ (.B(_0311_),
    .A(_0029_),
    .X(_0355_));
 sg13g2_nand2b_1 _2801_ (.Y(_0356_),
    .B(_0355_),
    .A_N(_0354_));
 sg13g2_a22oi_1 _2802_ (.Y(_0357_),
    .B1(_0352_),
    .B2(_0356_),
    .A2(_0310_),
    .A1(_1369_));
 sg13g2_nand2b_1 _2803_ (.Y(_0358_),
    .B(net327),
    .A_N(_0310_));
 sg13g2_o21ai_1 _2804_ (.B1(_0358_),
    .Y(_0359_),
    .A1(_0023_),
    .A2(_0309_));
 sg13g2_o21ai_1 _2805_ (.B1(_0347_),
    .Y(_0360_),
    .A1(_0357_),
    .A2(_0359_));
 sg13g2_a21oi_1 _2806_ (.A1(_0023_),
    .A2(_0309_),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_nand2_1 _2807_ (.Y(_0362_),
    .A(net351),
    .B(net352));
 sg13g2_nor2_1 _2808_ (.A(_0028_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_xor2_1 _2809_ (.B(_0363_),
    .A(net349),
    .X(_0364_));
 sg13g2_xnor2_1 _2810_ (.Y(_0365_),
    .A(net351),
    .B(net352));
 sg13g2_xnor2_1 _2811_ (.Y(_0366_),
    .A(\matt_venn_vga.digit_0.char[0] ),
    .B(_0365_));
 sg13g2_o21ai_1 _2812_ (.B1(_0366_),
    .Y(_0367_),
    .A1(net352),
    .A2(net317));
 sg13g2_a21oi_1 _2813_ (.A1(_1512_),
    .A2(_1513_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_xnor2_1 _2814_ (.Y(_0369_),
    .A(_0028_),
    .B(_0362_));
 sg13g2_a221oi_1 _2815_ (.B2(net312),
    .C1(_0368_),
    .B1(_0369_),
    .A1(net315),
    .Y(_0370_),
    .A2(_0365_));
 sg13g2_xnor2_1 _2816_ (.Y(_0371_),
    .A(_0055_),
    .B(_0364_));
 sg13g2_nor2_1 _2817_ (.A(_0370_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_o21ai_1 _2818_ (.B1(_0372_),
    .Y(_0373_),
    .A1(net312),
    .A2(_0369_));
 sg13g2_o21ai_1 _2819_ (.B1(_0373_),
    .Y(_0374_),
    .A1(_1390_),
    .A2(_0364_));
 sg13g2_nand4_1 _2820_ (.B(net350),
    .C(net351),
    .A(net349),
    .Y(_0375_),
    .D(net352));
 sg13g2_nor2b_1 _2821_ (.A(_1483_),
    .B_N(_0375_),
    .Y(_0376_));
 sg13g2_o21ai_1 _2822_ (.B1(_0374_),
    .Y(_0377_),
    .A1(_1518_),
    .A2(_0376_));
 sg13g2_a221oi_1 _2823_ (.B2(_1518_),
    .C1(\py[9] ),
    .B1(_0375_),
    .A1(\py[8] ),
    .Y(_0378_),
    .A2(_0308_));
 sg13g2_a21o_1 _2824_ (.A2(_0316_),
    .A1(_1368_),
    .B1(_0346_),
    .X(_0379_));
 sg13g2_nand4_1 _2825_ (.B(_0377_),
    .C(_0378_),
    .A(_1521_),
    .Y(_0380_),
    .D(_0379_));
 sg13g2_or3_2 _2826_ (.A(_0351_),
    .B(_0361_),
    .C(_0380_),
    .X(_0381_));
 sg13g2_o21ai_1 _2827_ (.B1(\product_comp[0] ),
    .Y(_0382_),
    .A1(_0283_),
    .A2(_0285_));
 sg13g2_a21oi_1 _2828_ (.A1(\product_comp[1] ),
    .A2(_0284_),
    .Y(_0383_),
    .B1(_1397_));
 sg13g2_nand4_1 _2829_ (.B(_0290_),
    .C(_0382_),
    .A(_0289_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_nor2_1 _2830_ (.A(_0278_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_a21oi_2 _2831_ (.B1(_0381_),
    .Y(_0386_),
    .A2(_0385_),
    .A1(_0264_));
 sg13g2_and2_2 _2832_ (.A(_0301_),
    .B(_0386_),
    .X(_0387_));
 sg13g2_nand3_1 _2833_ (.B(_0282_),
    .C(_0285_),
    .A(_1828_),
    .Y(_0388_));
 sg13g2_and4_1 _2834_ (.A(_0268_),
    .B(_0270_),
    .C(_0273_),
    .D(_0388_),
    .X(_0389_));
 sg13g2_a21oi_1 _2835_ (.A1(_0265_),
    .A2(_0389_),
    .Y(_0390_),
    .B1(_0262_));
 sg13g2_nand3b_1 _2836_ (.B(_0390_),
    .C(_0258_),
    .Y(_0391_),
    .A_N(_0381_));
 sg13g2_inv_1 _2837_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_a21oi_2 _2838_ (.B1(_0392_),
    .Y(_0393_),
    .A2(_0386_),
    .A1(_0301_));
 sg13g2_nand3_1 _2839_ (.B(net5),
    .C(\matt_venn_vga.activevideo ),
    .A(\matt_venn_vga.draw ),
    .Y(_0394_));
 sg13g2_nor2_1 _2840_ (.A(\matt_venn_vga.color[5] ),
    .B(\matt_venn_vga.color[0] ),
    .Y(_0395_));
 sg13g2_nor4_1 _2841_ (.A(\matt_venn_vga.color[1] ),
    .B(\matt_venn_vga.color[2] ),
    .C(\matt_venn_vga.color[3] ),
    .D(\matt_venn_vga.color[4] ),
    .Y(_0396_));
 sg13g2_a21oi_2 _2842_ (.B1(_0394_),
    .Y(_0397_),
    .A2(_0396_),
    .A1(_0395_));
 sg13g2_nor2_1 _2843_ (.A(\matt_venn_vga_shadow.color[0] ),
    .B(\matt_venn_vga_shadow.color[1] ),
    .Y(_0398_));
 sg13g2_nor4_1 _2844_ (.A(\matt_venn_vga_shadow.color[2] ),
    .B(\matt_venn_vga_shadow.color[3] ),
    .C(\matt_venn_vga_shadow.color[4] ),
    .D(\matt_venn_vga_shadow.color[5] ),
    .Y(_0399_));
 sg13g2_nand2_1 _2845_ (.Y(_0400_),
    .A(_0398_),
    .B(_0399_));
 sg13g2_nand4_1 _2846_ (.B(\matt_venn_vga_shadow.draw ),
    .C(\matt_venn_vga.activevideo ),
    .A(net5),
    .Y(_0401_),
    .D(_0400_));
 sg13g2_nand3b_1 _2847_ (.B(_0397_),
    .C(_0401_),
    .Y(_0402_),
    .A_N(_1477_));
 sg13g2_inv_1 _2848_ (.Y(_0403_),
    .A(_0402_));
 sg13g2_nand4_1 _2849_ (.B(\matt_venn_vga.color[5] ),
    .C(net5),
    .A(\matt_venn_vga.draw ),
    .Y(_0404_),
    .D(\matt_venn_vga.activevideo ));
 sg13g2_nand3_1 _2850_ (.B(_0402_),
    .C(_0404_),
    .A(_0393_),
    .Y(_0405_));
 sg13g2_a21oi_1 _2851_ (.A1(_1639_),
    .A2(_0405_),
    .Y(_0406_),
    .B1(_1638_));
 sg13g2_o21ai_1 _2852_ (.B1(_1451_),
    .Y(uo_out[0]),
    .A1(_1452_),
    .A2(_0406_));
 sg13g2_xnor2_1 _2853_ (.Y(_0407_),
    .A(net6),
    .B(\vga_sync.vsync ));
 sg13g2_nand2_1 _2854_ (.Y(_0408_),
    .A(net361),
    .B(_0407_));
 sg13g2_nor2b_1 _2855_ (.A(\matt_venn_vga.color[3] ),
    .B_N(_0397_),
    .Y(_0409_));
 sg13g2_nor2_1 _2856_ (.A(_0397_),
    .B(_0401_),
    .Y(_0410_));
 sg13g2_nand2_1 _2857_ (.Y(_0411_),
    .A(\t[1] ),
    .B(net322));
 sg13g2_xor2_1 _2858_ (.B(net321),
    .A(\t[2] ),
    .X(_0412_));
 sg13g2_nand2b_1 _2859_ (.Y(_0413_),
    .B(_0412_),
    .A_N(_0411_));
 sg13g2_o21ai_1 _2860_ (.B1(_0413_),
    .Y(_0414_),
    .A1(_1379_),
    .A2(_1394_));
 sg13g2_xnor2_1 _2861_ (.Y(_0415_),
    .A(net320),
    .B(_0030_));
 sg13g2_xnor2_1 _2862_ (.Y(_0416_),
    .A(\t[3] ),
    .B(_0415_));
 sg13g2_o21ai_1 _2863_ (.B1(net331),
    .Y(_0417_),
    .A1(_0414_),
    .A2(_0416_));
 sg13g2_a21o_1 _2864_ (.A2(_0416_),
    .A1(_0414_),
    .B1(_0417_),
    .X(_0418_));
 sg13g2_xnor2_1 _2865_ (.Y(_0419_),
    .A(net339),
    .B(_0032_));
 sg13g2_xnor2_1 _2866_ (.Y(_0420_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_xnor2_1 _2867_ (.Y(_0421_),
    .A(_0419_),
    .B(_0420_));
 sg13g2_xnor2_1 _2868_ (.Y(_0422_),
    .A(\t[1] ),
    .B(_1477_));
 sg13g2_xnor2_1 _2869_ (.Y(_0423_),
    .A(_0030_),
    .B(_0422_));
 sg13g2_nand3_1 _2870_ (.B(_0421_),
    .C(_0423_),
    .A(_0418_),
    .Y(_0424_));
 sg13g2_nand3_1 _2871_ (.B(_1431_),
    .C(_1439_),
    .A(_0029_),
    .Y(_0425_));
 sg13g2_o21ai_1 _2872_ (.B1(_0424_),
    .Y(_0426_),
    .A1(_0422_),
    .A2(_0425_));
 sg13g2_nor4_2 _2873_ (.A(net324),
    .B(net325),
    .C(net328),
    .Y(_0427_),
    .D(\matt_venn_vga.y_px[6] ));
 sg13g2_nand3b_1 _2874_ (.B(_0426_),
    .C(_0427_),
    .Y(_0428_),
    .A_N(_0397_));
 sg13g2_nand2b_1 _2875_ (.Y(_0429_),
    .B(_0428_),
    .A_N(_0410_));
 sg13g2_o21ai_1 _2876_ (.B1(_0402_),
    .Y(_0430_),
    .A1(_0409_),
    .A2(_0429_));
 sg13g2_nor2_1 _2877_ (.A(\product_comp[1] ),
    .B(\product_comp[0] ),
    .Y(_0431_));
 sg13g2_o21ai_1 _2878_ (.B1(\product_comp[2] ),
    .Y(_0432_),
    .A1(\product_comp[1] ),
    .A2(\product_comp[0] ));
 sg13g2_nand2_2 _2879_ (.Y(_0433_),
    .A(_1377_),
    .B(_0432_));
 sg13g2_nand4_1 _2880_ (.B(\product_comp[5] ),
    .C(\product_comp[4] ),
    .A(net344),
    .Y(_0434_),
    .D(_0433_));
 sg13g2_nand2_1 _2881_ (.Y(_0435_),
    .A(net344),
    .B(\product_comp[6] ));
 sg13g2_inv_1 _2882_ (.Y(_0436_),
    .A(_0435_));
 sg13g2_nand3_1 _2883_ (.B(_0434_),
    .C(_0435_),
    .A(_0065_),
    .Y(_0437_));
 sg13g2_nor3_2 _2884_ (.A(\product_comp[10] ),
    .B(\product_comp[9] ),
    .C(\product_comp[8] ),
    .Y(_0438_));
 sg13g2_nand2b_1 _2885_ (.Y(_0439_),
    .B(_0431_),
    .A_N(\product_comp[2] ));
 sg13g2_nand3_1 _2886_ (.B(_0436_),
    .C(_0439_),
    .A(\product_comp[3] ),
    .Y(_0440_));
 sg13g2_nand4_1 _2887_ (.B(_0434_),
    .C(_0435_),
    .A(_0065_),
    .Y(_0441_),
    .D(_0438_));
 sg13g2_a22oi_1 _2888_ (.Y(_0442_),
    .B1(_0441_),
    .B2(_0387_),
    .A2(_0430_),
    .A1(_0393_));
 sg13g2_a21oi_1 _2889_ (.A1(_1429_),
    .A2(_1454_),
    .Y(_0443_),
    .B1(net324));
 sg13g2_nor2_1 _2890_ (.A(net334),
    .B(_1458_),
    .Y(_0444_));
 sg13g2_a21o_1 _2891_ (.A2(_0444_),
    .A1(_1456_),
    .B1(_0443_),
    .X(_0445_));
 sg13g2_a21oi_1 _2892_ (.A1(_1441_),
    .A2(_1462_),
    .Y(_0446_),
    .B1(_1430_));
 sg13g2_nor4_1 _2893_ (.A(_1426_),
    .B(_1454_),
    .C(_1458_),
    .D(_1471_),
    .Y(_0447_));
 sg13g2_or3_1 _2894_ (.A(net323),
    .B(_0446_),
    .C(_0447_),
    .X(_0448_));
 sg13g2_inv_1 _2895_ (.Y(_0449_),
    .A(_0448_));
 sg13g2_xnor2_1 _2896_ (.Y(_0450_),
    .A(_1464_),
    .B(_1465_));
 sg13g2_xnor2_1 _2897_ (.Y(_0451_),
    .A(_0419_),
    .B(_0450_));
 sg13g2_xor2_1 _2898_ (.B(_1478_),
    .A(net337),
    .X(_0452_));
 sg13g2_nand3_1 _2899_ (.B(_0451_),
    .C(_0452_),
    .A(_0448_),
    .Y(_0453_));
 sg13g2_nand2_1 _2900_ (.Y(_0454_),
    .A(_0445_),
    .B(_0453_));
 sg13g2_a21oi_1 _2901_ (.A1(_1639_),
    .A2(_0442_),
    .Y(_0455_),
    .B1(_0454_));
 sg13g2_o21ai_1 _2902_ (.B1(_1453_),
    .Y(_0456_),
    .A1(_1637_),
    .A2(_0455_));
 sg13g2_nand2_2 _2903_ (.Y(uo_out[1]),
    .A(_0408_),
    .B(_0456_));
 sg13g2_o21ai_1 _2904_ (.B1(_0436_),
    .Y(_0457_),
    .A1(\product_comp[5] ),
    .A2(\product_comp[4] ));
 sg13g2_and2_1 _2905_ (.A(\product_comp[1] ),
    .B(\product_comp[0] ),
    .X(_0458_));
 sg13g2_nor4_1 _2906_ (.A(\product_comp[5] ),
    .B(\product_comp[3] ),
    .C(\product_comp[2] ),
    .D(_0458_),
    .Y(_0459_));
 sg13g2_or2_1 _2907_ (.X(_0460_),
    .B(_0459_),
    .A(_0457_));
 sg13g2_nor3_1 _2908_ (.A(\product_comp[9] ),
    .B(\product_comp[8] ),
    .C(_1397_),
    .Y(_0461_));
 sg13g2_nand4_1 _2909_ (.B(_0440_),
    .C(_0457_),
    .A(_0438_),
    .Y(_0462_),
    .D(_0461_));
 sg13g2_nor2b_1 _2910_ (.A(\matt_venn_vga.color[0] ),
    .B_N(_0397_),
    .Y(_0463_));
 sg13g2_nor4_1 _2911_ (.A(_0392_),
    .B(_0403_),
    .C(_0410_),
    .D(_0463_),
    .Y(_0464_));
 sg13g2_mux2_1 _2912_ (.A0(_0464_),
    .A1(_0462_),
    .S(_0387_),
    .X(_0465_));
 sg13g2_a21oi_1 _2913_ (.A1(_1639_),
    .A2(_0465_),
    .Y(_0466_),
    .B1(_1637_));
 sg13g2_nand2b_1 _2914_ (.Y(_0467_),
    .B(net4),
    .A_N(_0466_));
 sg13g2_nand3_1 _2915_ (.B(_0460_),
    .C(_0461_),
    .A(_0387_),
    .Y(_0468_));
 sg13g2_nor2b_1 _2916_ (.A(\matt_venn_vga.color[1] ),
    .B_N(_0397_),
    .Y(_0469_));
 sg13g2_o21ai_1 _2917_ (.B1(_0402_),
    .Y(_0470_),
    .A1(_0410_),
    .A2(_0469_));
 sg13g2_a21oi_1 _2918_ (.A1(_0391_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(_0387_));
 sg13g2_nor2_1 _2919_ (.A(_1640_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_a21oi_1 _2920_ (.A1(_0468_),
    .A2(_0472_),
    .Y(_0473_),
    .B1(_1637_));
 sg13g2_o21ai_1 _2921_ (.B1(_0467_),
    .Y(uo_out[2]),
    .A1(_1452_),
    .A2(_0473_));
 sg13g2_nor2_1 _2922_ (.A(net361),
    .B(_0407_),
    .Y(_0474_));
 sg13g2_a21oi_2 _2923_ (.B1(_0474_),
    .Y(uo_out[3]),
    .A2(_0473_),
    .A1(net361));
 sg13g2_a21oi_1 _2924_ (.A1(\matt_venn_vga.color[2] ),
    .A2(_0397_),
    .Y(_0475_),
    .B1(_0403_));
 sg13g2_a21oi_1 _2925_ (.A1(_0428_),
    .A2(_0475_),
    .Y(_0476_),
    .B1(_0410_));
 sg13g2_or2_1 _2926_ (.X(_0477_),
    .B(_0432_),
    .A(_1377_));
 sg13g2_nor3_2 _2927_ (.A(\product_comp[6] ),
    .B(\product_comp[5] ),
    .C(\product_comp[4] ),
    .Y(_0478_));
 sg13g2_a21oi_1 _2928_ (.A1(_0477_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(_0437_));
 sg13g2_a21o_1 _2929_ (.A2(_0479_),
    .A1(\product_comp[7] ),
    .B1(_0462_),
    .X(_0480_));
 sg13g2_a221oi_1 _2930_ (.B2(_0387_),
    .C1(_1640_),
    .B1(_0480_),
    .A1(_0393_),
    .Y(_0481_),
    .A2(_0476_));
 sg13g2_nor2b_1 _2931_ (.A(_1470_),
    .B_N(_0032_),
    .Y(_0482_));
 sg13g2_nor2b_1 _2932_ (.A(_0032_),
    .B_N(_1470_),
    .Y(_0483_));
 sg13g2_xor2_1 _2933_ (.B(_1478_),
    .A(_0031_),
    .X(_0484_));
 sg13g2_xor2_1 _2934_ (.B(_0030_),
    .A(net339),
    .X(_0485_));
 sg13g2_xnor2_1 _2935_ (.Y(_0486_),
    .A(_0450_),
    .B(_0485_));
 sg13g2_nor4_1 _2936_ (.A(_0482_),
    .B(_0483_),
    .C(_0484_),
    .D(_0486_),
    .Y(_0487_));
 sg13g2_o21ai_1 _2937_ (.B1(_0449_),
    .Y(_0488_),
    .A1(_1639_),
    .A2(_0487_));
 sg13g2_o21ai_1 _2938_ (.B1(_0453_),
    .Y(_0489_),
    .A1(_0481_),
    .A2(_0488_));
 sg13g2_a21oi_1 _2939_ (.A1(_0445_),
    .A2(_0489_),
    .Y(_0490_),
    .B1(_1638_));
 sg13g2_nor2b_1 _2940_ (.A(\matt_venn_vga.color[4] ),
    .B_N(_0397_),
    .Y(_0491_));
 sg13g2_o21ai_1 _2941_ (.B1(_0402_),
    .Y(_0492_),
    .A1(_0429_),
    .A2(_0491_));
 sg13g2_a21o_1 _2942_ (.A2(_0492_),
    .A1(_0391_),
    .B1(_1640_),
    .X(_0493_));
 sg13g2_o21ai_1 _2943_ (.B1(_0449_),
    .Y(_0494_),
    .A1(_0387_),
    .A2(_0493_));
 sg13g2_a21oi_1 _2944_ (.A1(_0445_),
    .A2(_0494_),
    .Y(_0495_),
    .B1(_1482_));
 sg13g2_o21ai_1 _2945_ (.B1(_1453_),
    .Y(_0496_),
    .A1(_1637_),
    .A2(_0495_));
 sg13g2_o21ai_1 _2946_ (.B1(_0496_),
    .Y(uo_out[4]),
    .A1(_1403_),
    .A2(_0490_));
 sg13g2_o21ai_1 _2947_ (.B1(net4),
    .Y(_0497_),
    .A1(_1637_),
    .A2(_0455_));
 sg13g2_o21ai_1 _2948_ (.B1(_0497_),
    .Y(uo_out[5]),
    .A1(_1452_),
    .A2(_0490_));
 sg13g2_o21ai_1 _2949_ (.B1(net361),
    .Y(_0498_),
    .A1(_1637_),
    .A2(_0495_));
 sg13g2_o21ai_1 _2950_ (.B1(_0498_),
    .Y(uo_out[6]),
    .A1(_1452_),
    .A2(_0466_));
 sg13g2_nor2_1 _2951_ (.A(_0070_),
    .B(net361),
    .Y(_0499_));
 sg13g2_a21oi_2 _2952_ (.B1(_0499_),
    .Y(uo_out[7]),
    .A2(_0406_),
    .A1(net361));
 sg13g2_xnor2_1 _2953_ (.Y(_0500_),
    .A(_0055_),
    .B(_1416_));
 sg13g2_xor2_1 _2954_ (.B(net309),
    .A(\matt_venn_vga.x_px[8] ),
    .X(_0501_));
 sg13g2_nor2_1 _2955_ (.A(net309),
    .B(_1416_),
    .Y(_0502_));
 sg13g2_a21oi_2 _2956_ (.B1(_0502_),
    .Y(_0503_),
    .A2(_0501_),
    .A1(_1416_));
 sg13g2_nor2_2 _2957_ (.A(_0500_),
    .B(net306),
    .Y(_0504_));
 sg13g2_or2_1 _2958_ (.X(_0505_),
    .B(net306),
    .A(_0500_));
 sg13g2_nor2_1 _2959_ (.A(net319),
    .B(net320),
    .Y(_0506_));
 sg13g2_nand2_2 _2960_ (.Y(_0507_),
    .A(_1392_),
    .B(_0506_));
 sg13g2_nor3_2 _2961_ (.A(net313),
    .B(net316),
    .C(_0507_),
    .Y(_0508_));
 sg13g2_o21ai_1 _2962_ (.B1(net313),
    .Y(_0509_),
    .A1(net316),
    .A2(_0507_));
 sg13g2_and2_2 _2963_ (.A(_1391_),
    .B(_0509_),
    .X(_0510_));
 sg13g2_inv_1 _2964_ (.Y(_0511_),
    .A(_0510_));
 sg13g2_o21ai_1 _2965_ (.B1(_0504_),
    .Y(_0512_),
    .A1(_0508_),
    .A2(_0511_));
 sg13g2_xnor2_1 _2966_ (.Y(_0513_),
    .A(_1391_),
    .B(_0509_));
 sg13g2_nor2_1 _2967_ (.A(net309),
    .B(_0510_),
    .Y(_0514_));
 sg13g2_nor2_1 _2968_ (.A(net309),
    .B(_0513_),
    .Y(_0515_));
 sg13g2_or2_1 _2969_ (.X(_0516_),
    .B(_0513_),
    .A(net309));
 sg13g2_nor2b_2 _2970_ (.A(_0508_),
    .B_N(_0509_),
    .Y(_0517_));
 sg13g2_nor2b_1 _2971_ (.A(net306),
    .B_N(_0500_),
    .Y(_0518_));
 sg13g2_nor2b_2 _2972_ (.A(_0517_),
    .B_N(_0518_),
    .Y(_0519_));
 sg13g2_a21o_2 _2973_ (.A2(_0510_),
    .A1(_0501_),
    .B1(_0514_),
    .X(_0520_));
 sg13g2_a21oi_2 _2974_ (.B1(_0514_),
    .Y(_0521_),
    .A2(_0510_),
    .A1(_0501_));
 sg13g2_a21o_1 _2975_ (.A2(_0520_),
    .A1(_0041_),
    .B1(_0519_),
    .X(_0522_));
 sg13g2_xnor2_1 _2976_ (.Y(_0523_),
    .A(_0055_),
    .B(_0510_));
 sg13g2_or2_2 _2977_ (.X(_0524_),
    .B(_0523_),
    .A(_0521_));
 sg13g2_nor2_2 _2978_ (.A(_0516_),
    .B(_0517_),
    .Y(_0525_));
 sg13g2_a22oi_1 _2979_ (.Y(_0526_),
    .B1(_0525_),
    .B2(_0040_),
    .A2(_0522_),
    .A1(_0516_));
 sg13g2_nand2_1 _2980_ (.Y(_0527_),
    .A(_0524_),
    .B(_0526_));
 sg13g2_nand2_2 _2981_ (.Y(_0528_),
    .A(net313),
    .B(_1391_));
 sg13g2_nor2_1 _2982_ (.A(net303),
    .B(_0528_),
    .Y(_0529_));
 sg13g2_or2_2 _2983_ (.X(_0530_),
    .B(_0528_),
    .A(net303));
 sg13g2_or2_1 _2984_ (.X(_0246_),
    .B(_0503_),
    .A(net382));
 sg13g2_nand2b_1 _2985_ (.Y(_0531_),
    .B(net312),
    .A_N(net314));
 sg13g2_nor2_1 _2986_ (.A(net316),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nand2_1 _2987_ (.Y(_0533_),
    .A(_0055_),
    .B(_0532_));
 sg13g2_or2_1 _2988_ (.X(_0534_),
    .B(_0533_),
    .A(_0246_));
 sg13g2_a21o_2 _2989_ (.A2(_0534_),
    .A1(_0530_),
    .B1(_0517_),
    .X(_0535_));
 sg13g2_nor2_1 _2990_ (.A(net303),
    .B(_0513_),
    .Y(_0536_));
 sg13g2_a22oi_1 _2991_ (.Y(_0537_),
    .B1(_0536_),
    .B2(_0039_),
    .A2(_0527_),
    .A1(_0512_));
 sg13g2_nand2_1 _2992_ (.Y(_0538_),
    .A(_0535_),
    .B(_0537_));
 sg13g2_nor3_1 _2993_ (.A(_0042_),
    .B(net303),
    .C(_0513_),
    .Y(_0539_));
 sg13g2_nor2_1 _2994_ (.A(_0046_),
    .B(_0521_),
    .Y(_0540_));
 sg13g2_o21ai_1 _2995_ (.B1(_0516_),
    .Y(_0541_),
    .A1(_0519_),
    .A2(_0540_));
 sg13g2_a21oi_1 _2996_ (.A1(_0045_),
    .A2(_0519_),
    .Y(_0542_),
    .B1(_0541_));
 sg13g2_a21oi_1 _2997_ (.A1(_1404_),
    .A2(_0525_),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_o21ai_1 _2998_ (.B1(_0512_),
    .Y(_0544_),
    .A1(_1405_),
    .A2(_0524_));
 sg13g2_a21oi_1 _2999_ (.A1(_0524_),
    .A2(_0543_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_or2_2 _3000_ (.X(_0546_),
    .B(_0545_),
    .A(_0539_));
 sg13g2_nand2b_1 _3001_ (.Y(_0547_),
    .B(_0546_),
    .A_N(_0538_));
 sg13g2_nand3b_1 _3002_ (.B(_0520_),
    .C(_0038_),
    .Y(_0548_),
    .A_N(_0519_));
 sg13g2_a21oi_1 _3003_ (.A1(_0072_),
    .A2(_0519_),
    .Y(_0549_),
    .B1(_0515_));
 sg13g2_a22oi_1 _3004_ (.Y(_0550_),
    .B1(_0548_),
    .B2(_0549_),
    .A2(_0525_),
    .A1(\clock_min_u[0] ));
 sg13g2_o21ai_1 _3005_ (.B1(_0512_),
    .Y(_0551_),
    .A1(\clock_min_d[0] ),
    .A2(_0524_));
 sg13g2_a21oi_1 _3006_ (.A1(_0524_),
    .A2(_0550_),
    .Y(_0552_),
    .B1(_0551_));
 sg13g2_a21oi_1 _3007_ (.A1(\clock_hrs_u[0] ),
    .A2(_0536_),
    .Y(_0553_),
    .B1(_0552_));
 sg13g2_nand2_1 _3008_ (.Y(_0554_),
    .A(_0535_),
    .B(_0553_));
 sg13g2_o21ai_1 _3009_ (.B1(_0554_),
    .Y(_0555_),
    .A1(\clock_hrs_d[0] ),
    .A2(_0535_));
 sg13g2_nor2b_1 _3010_ (.A(_0555_),
    .B_N(_0547_),
    .Y(_0011_));
 sg13g2_nor2b_1 _3011_ (.A(\clock_sec_d[1] ),
    .B_N(_0519_),
    .Y(_0556_));
 sg13g2_nor3_1 _3012_ (.A(\clock_sec_u[1] ),
    .B(_0519_),
    .C(_0521_),
    .Y(_0557_));
 sg13g2_o21ai_1 _3013_ (.B1(_0516_),
    .Y(_0558_),
    .A1(_0556_),
    .A2(_0557_));
 sg13g2_nand2b_1 _3014_ (.Y(_0559_),
    .B(_0525_),
    .A_N(\clock_min_u[1] ));
 sg13g2_nand3_1 _3015_ (.B(_0558_),
    .C(_0559_),
    .A(_0524_),
    .Y(_0560_));
 sg13g2_o21ai_1 _3016_ (.B1(_0512_),
    .Y(_0561_),
    .A1(_1350_),
    .A2(_0524_));
 sg13g2_nand2b_1 _3017_ (.Y(_0562_),
    .B(_0560_),
    .A_N(_0561_));
 sg13g2_nand2_1 _3018_ (.Y(_0563_),
    .A(_0048_),
    .B(_0536_));
 sg13g2_nand3_1 _3019_ (.B(_0562_),
    .C(_0563_),
    .A(_0535_),
    .Y(_0564_));
 sg13g2_o21ai_1 _3020_ (.B1(_0564_),
    .Y(_0565_),
    .A1(_0047_),
    .A2(_0535_));
 sg13g2_and2_1 _3021_ (.A(_0547_),
    .B(_0565_),
    .X(_0012_));
 sg13g2_nand2_1 _3022_ (.Y(_0566_),
    .A(_0535_),
    .B(_0546_));
 sg13g2_nor2_1 _3023_ (.A(_0555_),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_nand3_1 _3024_ (.B(_0538_),
    .C(_0546_),
    .A(_0535_),
    .Y(_0568_));
 sg13g2_inv_1 _3025_ (.Y(_0569_),
    .A(_0568_));
 sg13g2_a21oi_1 _3026_ (.A1(_0555_),
    .A2(_0568_),
    .Y(_0013_),
    .B1(_0567_));
 sg13g2_o21ai_1 _3027_ (.B1(_0538_),
    .Y(_0570_),
    .A1(_0555_),
    .A2(_0566_));
 sg13g2_nor2_1 _3028_ (.A(_0565_),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_nand2b_1 _3029_ (.Y(_0572_),
    .B(_0547_),
    .A_N(_0565_));
 sg13g2_a21oi_1 _3030_ (.A1(_0570_),
    .A2(_0572_),
    .Y(_0014_),
    .B1(_0571_));
 sg13g2_nor2_1 _3031_ (.A(_0538_),
    .B(_0546_),
    .Y(_0573_));
 sg13g2_nand2_1 _3032_ (.Y(_0574_),
    .A(_0565_),
    .B(_0573_));
 sg13g2_nor2b_1 _3033_ (.A(_0555_),
    .B_N(_0565_),
    .Y(_0575_));
 sg13g2_o21ai_1 _3034_ (.B1(_0574_),
    .Y(_0015_),
    .A1(_0568_),
    .A2(_0575_));
 sg13g2_a21o_1 _3035_ (.A2(_0575_),
    .A1(_0569_),
    .B1(_0573_),
    .X(_0016_));
 sg13g2_nand2_1 _3036_ (.Y(_0576_),
    .A(net555),
    .B(_1606_));
 sg13g2_xnor2_1 _3037_ (.Y(_0577_),
    .A(_1369_),
    .B(_1606_));
 sg13g2_nor2_1 _3038_ (.A(_1441_),
    .B(_1606_),
    .Y(_0578_));
 sg13g2_xnor2_1 _3039_ (.Y(_0579_),
    .A(_0069_),
    .B(_1440_));
 sg13g2_xnor2_1 _3040_ (.Y(_0580_),
    .A(net333),
    .B(net334));
 sg13g2_nand2_1 _3041_ (.Y(_0581_),
    .A(\matt_venn_vga.digit_0.digit_index[0] ),
    .B(_0580_));
 sg13g2_xor2_1 _3042_ (.B(_0579_),
    .A(\matt_venn_vga.digit_0.digit_index[1] ),
    .X(_0582_));
 sg13g2_nor2b_1 _3043_ (.A(_0581_),
    .B_N(_0582_),
    .Y(_0583_));
 sg13g2_a21o_1 _3044_ (.A2(_0579_),
    .A1(\matt_venn_vga.digit_0.digit_index[1] ),
    .B1(_0583_),
    .X(_0584_));
 sg13g2_xnor2_1 _3045_ (.Y(_0585_),
    .A(\matt_venn_vga.digit_0.digit_index[2] ),
    .B(_0578_));
 sg13g2_nor2b_1 _3046_ (.A(_0585_),
    .B_N(_0584_),
    .Y(_0586_));
 sg13g2_a21o_1 _3047_ (.A2(_0578_),
    .A1(\matt_venn_vga.digit_0.digit_index[2] ),
    .B1(_0586_),
    .X(_0587_));
 sg13g2_xnor2_1 _3048_ (.Y(_0588_),
    .A(\matt_venn_vga.digit_0.digit_index[3] ),
    .B(_0577_));
 sg13g2_nor2b_1 _3049_ (.A(_0588_),
    .B_N(_0587_),
    .Y(_0589_));
 sg13g2_a21oi_1 _3050_ (.A1(\matt_venn_vga.digit_0.digit_index[3] ),
    .A2(_0577_),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_xor2_1 _3051_ (.B(_0576_),
    .A(net325),
    .X(_0591_));
 sg13g2_nand2_1 _3052_ (.Y(_0592_),
    .A(\matt_venn_vga.digit_0.digit_index[4] ),
    .B(_0591_));
 sg13g2_xnor2_1 _3053_ (.Y(_0593_),
    .A(\matt_venn_vga.digit_0.digit_index[4] ),
    .B(_0591_));
 sg13g2_xor2_1 _3054_ (.B(_0593_),
    .A(_0590_),
    .X(_0594_));
 sg13g2_xnor2_1 _3055_ (.Y(_0595_),
    .A(_0581_),
    .B(_0582_));
 sg13g2_xor2_1 _3056_ (.B(_0580_),
    .A(\matt_venn_vga.digit_0.digit_index[0] ),
    .X(_0596_));
 sg13g2_nor2_1 _3057_ (.A(_0595_),
    .B(_0596_),
    .Y(_0597_));
 sg13g2_xor2_1 _3058_ (.B(_0588_),
    .A(_0587_),
    .X(_0598_));
 sg13g2_o21ai_1 _3059_ (.B1(_0592_),
    .Y(_0599_),
    .A1(_0590_),
    .A2(_0593_));
 sg13g2_o21ai_1 _3060_ (.B1(_0023_),
    .Y(_0600_),
    .A1(net325),
    .A2(_0576_));
 sg13g2_xor2_1 _3061_ (.B(_0600_),
    .A(_0057_),
    .X(_0601_));
 sg13g2_xnor2_1 _3062_ (.Y(_0602_),
    .A(\matt_venn_vga.digit_0.digit_index[5] ),
    .B(_0601_));
 sg13g2_xnor2_1 _3063_ (.Y(_0603_),
    .A(_0599_),
    .B(_0602_));
 sg13g2_o21ai_1 _3064_ (.B1(_0597_),
    .Y(_0604_),
    .A1(net287),
    .A2(_0603_));
 sg13g2_xnor2_1 _3065_ (.Y(_0605_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_xor2_1 _3066_ (.B(_0585_),
    .A(_0584_),
    .X(_0606_));
 sg13g2_nor2_1 _3067_ (.A(_0597_),
    .B(_0605_),
    .Y(_0607_));
 sg13g2_nand2b_1 _3068_ (.Y(_0608_),
    .B(_0605_),
    .A_N(net287));
 sg13g2_nor2b_2 _3069_ (.A(_0582_),
    .B_N(_0596_),
    .Y(_0609_));
 sg13g2_o21ai_1 _3070_ (.B1(_0604_),
    .Y(_0610_),
    .A1(_0608_),
    .A2(_0609_));
 sg13g2_nor2_1 _3071_ (.A(_0607_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_nand2_1 _3072_ (.Y(_0612_),
    .A(_0596_),
    .B(_0606_));
 sg13g2_nand2_1 _3073_ (.Y(_0613_),
    .A(_0595_),
    .B(_0612_));
 sg13g2_o21ai_1 _3074_ (.B1(_0594_),
    .Y(_0614_),
    .A1(net287),
    .A2(_0613_));
 sg13g2_nor2_1 _3075_ (.A(_0603_),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_nand2b_1 _3076_ (.Y(_0616_),
    .B(net287),
    .A_N(_0595_));
 sg13g2_o21ai_1 _3077_ (.B1(_0608_),
    .Y(_0617_),
    .A1(_0605_),
    .A2(_0616_));
 sg13g2_a21oi_1 _3078_ (.A1(_0603_),
    .A2(_0617_),
    .Y(_0618_),
    .B1(_0615_));
 sg13g2_o21ai_1 _3079_ (.B1(_0618_),
    .Y(_0008_),
    .A1(_0594_),
    .A2(_0611_));
 sg13g2_nand2b_1 _3080_ (.Y(_0619_),
    .B(_0612_),
    .A_N(_0609_));
 sg13g2_inv_1 _3081_ (.Y(_0620_),
    .A(_0619_));
 sg13g2_o21ai_1 _3082_ (.B1(_0619_),
    .Y(_0621_),
    .A1(_0582_),
    .A2(_0605_));
 sg13g2_nor2_1 _3083_ (.A(_0605_),
    .B(_0609_),
    .Y(_0622_));
 sg13g2_xnor2_1 _3084_ (.Y(_0623_),
    .A(_0606_),
    .B(_0609_));
 sg13g2_nand2b_1 _3085_ (.Y(_0624_),
    .B(_0595_),
    .A_N(_0596_));
 sg13g2_o21ai_1 _3086_ (.B1(_0612_),
    .Y(_0625_),
    .A1(_0606_),
    .A2(_0624_));
 sg13g2_mux4_1 _3087_ (.S0(_0594_),
    .A0(_0625_),
    .A1(_0606_),
    .A2(_0623_),
    .A3(_0621_),
    .S1(net288),
    .X(_0626_));
 sg13g2_a21oi_1 _3088_ (.A1(net288),
    .A2(_0607_),
    .Y(_0627_),
    .B1(_0594_));
 sg13g2_o21ai_1 _3089_ (.B1(_0627_),
    .Y(_0628_),
    .A1(net287),
    .A2(_0621_));
 sg13g2_nand2_1 _3090_ (.Y(_0629_),
    .A(net288),
    .B(_0625_));
 sg13g2_o21ai_1 _3091_ (.B1(_0629_),
    .Y(_0630_),
    .A1(net287),
    .A2(_0620_));
 sg13g2_a21oi_1 _3092_ (.A1(_0594_),
    .A2(_0630_),
    .Y(_0631_),
    .B1(_0603_));
 sg13g2_a22oi_1 _3093_ (.Y(_0009_),
    .B1(_0628_),
    .B2(_0631_),
    .A2(_0626_),
    .A1(_0603_));
 sg13g2_nor2_1 _3094_ (.A(_0606_),
    .B(_0616_),
    .Y(_0632_));
 sg13g2_a21oi_1 _3095_ (.A1(_0594_),
    .A2(_0608_),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_o21ai_1 _3096_ (.B1(_0620_),
    .Y(_0634_),
    .A1(_0596_),
    .A2(_0606_));
 sg13g2_o21ai_1 _3097_ (.B1(_0594_),
    .Y(_0635_),
    .A1(_0597_),
    .A2(net287));
 sg13g2_a21oi_1 _3098_ (.A1(net288),
    .A2(_0634_),
    .Y(_0636_),
    .B1(_0635_));
 sg13g2_nand3b_1 _3099_ (.B(_0622_),
    .C(_0624_),
    .Y(_0637_),
    .A_N(net288));
 sg13g2_nand3_1 _3100_ (.B(net287),
    .C(_0605_),
    .A(_0595_),
    .Y(_0638_));
 sg13g2_a21oi_1 _3101_ (.A1(_0637_),
    .A2(_0638_),
    .Y(_0639_),
    .B1(_0594_));
 sg13g2_nor3_1 _3102_ (.A(_0603_),
    .B(_0636_),
    .C(_0639_),
    .Y(_0640_));
 sg13g2_a21o_1 _3103_ (.A2(_0633_),
    .A1(_0603_),
    .B1(_0640_),
    .X(_0010_));
 sg13g2_nand2_1 _3104_ (.Y(_0641_),
    .A(_1423_),
    .B(_1439_));
 sg13g2_a21oi_2 _3105_ (.B1(_1370_),
    .Y(_0642_),
    .A2(_1439_),
    .A1(_1423_));
 sg13g2_xnor2_1 _3106_ (.Y(_0643_),
    .A(net517),
    .B(_0642_));
 sg13g2_nand2_1 _3107_ (.Y(_0644_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[3] ),
    .B(_0643_));
 sg13g2_xnor2_1 _3108_ (.Y(_0645_),
    .A(_1370_),
    .B(_0641_));
 sg13g2_nand2_1 _3109_ (.Y(_0646_),
    .A(_0026_),
    .B(_1423_));
 sg13g2_xnor2_1 _3110_ (.Y(_0647_),
    .A(_1402_),
    .B(_0646_));
 sg13g2_nand2_1 _3111_ (.Y(_0648_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[1] ),
    .B(_0647_));
 sg13g2_xnor2_1 _3112_ (.Y(_0649_),
    .A(net332),
    .B(_1422_));
 sg13g2_nand2_1 _3113_ (.Y(_0650_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[0] ),
    .B(_0649_));
 sg13g2_xnor2_1 _3114_ (.Y(_0651_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[1] ),
    .B(_0647_));
 sg13g2_inv_1 _3115_ (.Y(_0652_),
    .A(_0651_));
 sg13g2_o21ai_1 _3116_ (.B1(_0648_),
    .Y(_0653_),
    .A1(_0650_),
    .A2(_0651_));
 sg13g2_xnor2_1 _3117_ (.Y(_0654_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[2] ),
    .B(_0645_));
 sg13g2_nor2b_1 _3118_ (.A(_0654_),
    .B_N(_0653_),
    .Y(_0655_));
 sg13g2_a21oi_1 _3119_ (.A1(\matt_venn_vga_shadow.digit_0.digit_index[2] ),
    .A2(_0645_),
    .Y(_0656_),
    .B1(_0655_));
 sg13g2_xnor2_1 _3120_ (.Y(_0657_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[3] ),
    .B(_0643_));
 sg13g2_o21ai_1 _3121_ (.B1(_0644_),
    .Y(_0658_),
    .A1(_0656_),
    .A2(_0657_));
 sg13g2_nand2_1 _3122_ (.Y(_0659_),
    .A(net327),
    .B(_0642_));
 sg13g2_xor2_1 _3123_ (.B(_0659_),
    .A(_0023_),
    .X(_0660_));
 sg13g2_nor2b_1 _3124_ (.A(_0660_),
    .B_N(\matt_venn_vga_shadow.digit_0.digit_index[4] ),
    .Y(_0661_));
 sg13g2_xnor2_1 _3125_ (.Y(_0662_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[4] ),
    .B(_0660_));
 sg13g2_xor2_1 _3126_ (.B(_0662_),
    .A(_0658_),
    .X(_0663_));
 sg13g2_xor2_1 _3127_ (.B(_0651_),
    .A(_0650_),
    .X(_0664_));
 sg13g2_xor2_1 _3128_ (.B(_0649_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[0] ),
    .X(_0665_));
 sg13g2_xnor2_1 _3129_ (.Y(_0666_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[0] ),
    .B(_0649_));
 sg13g2_nor2_1 _3130_ (.A(_0664_),
    .B(_0665_),
    .Y(_0667_));
 sg13g2_xor2_1 _3131_ (.B(_0657_),
    .A(_0656_),
    .X(_0668_));
 sg13g2_a21oi_1 _3132_ (.A1(_0658_),
    .A2(_0662_),
    .Y(_0669_),
    .B1(_0661_));
 sg13g2_a21oi_1 _3133_ (.A1(net327),
    .A2(_0642_),
    .Y(_0670_),
    .B1(net326));
 sg13g2_xnor2_1 _3134_ (.Y(_0671_),
    .A(_0057_),
    .B(_0670_));
 sg13g2_xor2_1 _3135_ (.B(_0671_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[5] ),
    .X(_0672_));
 sg13g2_xnor2_1 _3136_ (.Y(_0673_),
    .A(_0669_),
    .B(_0672_));
 sg13g2_inv_1 _3137_ (.Y(_0674_),
    .A(_0673_));
 sg13g2_nand2_1 _3138_ (.Y(_0675_),
    .A(_0668_),
    .B(_0674_));
 sg13g2_xnor2_1 _3139_ (.Y(_0676_),
    .A(_0653_),
    .B(_0654_));
 sg13g2_or2_1 _3140_ (.X(_0677_),
    .B(net298),
    .A(_0667_));
 sg13g2_and2_1 _3141_ (.A(_0668_),
    .B(net298),
    .X(_0678_));
 sg13g2_nand2_2 _3142_ (.Y(_0679_),
    .A(_0651_),
    .B(_0665_));
 sg13g2_a22oi_1 _3143_ (.Y(_0680_),
    .B1(_0678_),
    .B2(_0679_),
    .A2(_0675_),
    .A1(_0667_));
 sg13g2_and2_1 _3144_ (.A(_0677_),
    .B(_0680_),
    .X(_0681_));
 sg13g2_nor2_1 _3145_ (.A(_0666_),
    .B(net298),
    .Y(_0682_));
 sg13g2_nand2_1 _3146_ (.Y(_0683_),
    .A(_0664_),
    .B(_0668_));
 sg13g2_o21ai_1 _3147_ (.B1(_0663_),
    .Y(_0684_),
    .A1(_0682_),
    .A2(_0683_));
 sg13g2_or2_1 _3148_ (.X(_0685_),
    .B(_0668_),
    .A(_0664_));
 sg13g2_inv_1 _3149_ (.Y(_0686_),
    .A(_0685_));
 sg13g2_o21ai_1 _3150_ (.B1(_0673_),
    .Y(_0687_),
    .A1(net299),
    .A2(_0685_));
 sg13g2_nor2_1 _3151_ (.A(_0678_),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_a21o_1 _3152_ (.A2(_0684_),
    .A1(_0674_),
    .B1(_0688_),
    .X(_0689_));
 sg13g2_o21ai_1 _3153_ (.B1(_0689_),
    .Y(_0019_),
    .A1(_0663_),
    .A2(_0681_));
 sg13g2_a21oi_1 _3154_ (.A1(_0652_),
    .A2(net299),
    .Y(_0690_),
    .B1(_0666_));
 sg13g2_o21ai_1 _3155_ (.B1(_0690_),
    .Y(_0691_),
    .A1(_0652_),
    .A2(net298));
 sg13g2_and2_1 _3156_ (.A(_0664_),
    .B(_0666_),
    .X(_0692_));
 sg13g2_a21o_1 _3157_ (.A2(_0692_),
    .A1(net298),
    .B1(_0682_),
    .X(_0693_));
 sg13g2_mux4_1 _3158_ (.S0(_0668_),
    .A0(_0677_),
    .A1(_0691_),
    .A2(_0693_),
    .A3(_0690_),
    .S1(_0663_),
    .X(_0694_));
 sg13g2_inv_1 _3159_ (.Y(_0695_),
    .A(_0694_));
 sg13g2_nor2b_1 _3160_ (.A(_0678_),
    .B_N(_0663_),
    .Y(_0696_));
 sg13g2_o21ai_1 _3161_ (.B1(_0696_),
    .Y(_0697_),
    .A1(_0668_),
    .A2(_0691_));
 sg13g2_nand2b_1 _3162_ (.Y(_0698_),
    .B(_0679_),
    .A_N(net298));
 sg13g2_xnor2_1 _3163_ (.Y(_0699_),
    .A(net298),
    .B(_0679_));
 sg13g2_mux2_1 _3164_ (.A0(_0699_),
    .A1(_0693_),
    .S(_0668_),
    .X(_0700_));
 sg13g2_nand2b_1 _3165_ (.Y(_0701_),
    .B(_0700_),
    .A_N(_0663_));
 sg13g2_nand3_1 _3166_ (.B(_0697_),
    .C(_0701_),
    .A(_0673_),
    .Y(_0702_));
 sg13g2_o21ai_1 _3167_ (.B1(_0702_),
    .Y(_0020_),
    .A1(_0673_),
    .A2(_0695_));
 sg13g2_a21oi_1 _3168_ (.A1(_0666_),
    .A2(net299),
    .Y(_0703_),
    .B1(_0690_));
 sg13g2_and2_1 _3169_ (.A(_0664_),
    .B(net298),
    .X(_0704_));
 sg13g2_nor2_1 _3170_ (.A(_0692_),
    .B(_0698_),
    .Y(_0705_));
 sg13g2_a21oi_1 _3171_ (.A1(net299),
    .A2(_0686_),
    .Y(_0706_),
    .B1(_0696_));
 sg13g2_mux4_1 _3172_ (.S0(_0668_),
    .A0(_0704_),
    .A1(_0705_),
    .A2(_0703_),
    .A3(_0667_),
    .S1(_0663_),
    .X(_0707_));
 sg13g2_nand2_1 _3173_ (.Y(_0708_),
    .A(_0673_),
    .B(_0706_));
 sg13g2_o21ai_1 _3174_ (.B1(_0708_),
    .Y(_0021_),
    .A1(_0673_),
    .A2(_0707_));
 sg13g2_and2_1 _3175_ (.A(\clock_color_offset[0] ),
    .B(_0517_),
    .X(_0709_));
 sg13g2_xor2_1 _3176_ (.B(_0517_),
    .A(\clock_color_offset[0] ),
    .X(_0710_));
 sg13g2_xor2_1 _3177_ (.B(_0513_),
    .A(net563),
    .X(_0711_));
 sg13g2_nand2_1 _3178_ (.Y(_0712_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_inv_1 _3179_ (.Y(_0713_),
    .A(_0712_));
 sg13g2_a22oi_1 _3180_ (.Y(_0714_),
    .B1(_0709_),
    .B2(_0711_),
    .A2(_0513_),
    .A1(_1393_));
 sg13g2_xnor2_1 _3181_ (.Y(_0715_),
    .A(_1351_),
    .B(_0523_));
 sg13g2_xnor2_1 _3182_ (.Y(_0716_),
    .A(_0714_),
    .B(_0715_));
 sg13g2_inv_1 _3183_ (.Y(_0717_),
    .A(_0716_));
 sg13g2_xnor2_1 _3184_ (.Y(_0718_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_a21oi_1 _3185_ (.A1(_0716_),
    .A2(_0718_),
    .Y(_0017_),
    .B1(_0713_));
 sg13g2_nand2_1 _3186_ (.Y(_0719_),
    .A(_0710_),
    .B(_0716_));
 sg13g2_o21ai_1 _3187_ (.B1(_0719_),
    .Y(_0018_),
    .A1(_0713_),
    .A2(_0716_));
 sg13g2_nand2_2 _3188_ (.Y(_0720_),
    .A(_0055_),
    .B(_0502_));
 sg13g2_nor2b_2 _3189_ (.A(_0720_),
    .B_N(_1417_),
    .Y(_0721_));
 sg13g2_nand2b_1 _3190_ (.Y(_0722_),
    .B(_0721_),
    .A_N(_0042_));
 sg13g2_and2_1 _3191_ (.A(net314),
    .B(_0518_),
    .X(_0723_));
 sg13g2_nand2_1 _3192_ (.Y(_0724_),
    .A(net313),
    .B(_0518_));
 sg13g2_o21ai_1 _3193_ (.B1(_0724_),
    .Y(_0725_),
    .A1(_0046_),
    .A2(net306));
 sg13g2_a21oi_2 _3194_ (.B1(net306),
    .Y(_0726_),
    .A2(_0500_),
    .A1(_1418_));
 sg13g2_a21oi_1 _3195_ (.A1(_0045_),
    .A2(_0723_),
    .Y(_0727_),
    .B1(_0726_));
 sg13g2_o21ai_1 _3196_ (.B1(_0505_),
    .Y(_0728_),
    .A1(net309),
    .A2(_0528_));
 sg13g2_a221oi_1 _3197_ (.B2(_1404_),
    .C1(_0504_),
    .B1(_0728_),
    .A1(_0725_),
    .Y(_0729_),
    .A2(_0727_));
 sg13g2_o21ai_1 _3198_ (.B1(_0720_),
    .Y(_0730_),
    .A1(_1405_),
    .A2(net303));
 sg13g2_o21ai_1 _3199_ (.B1(_0722_),
    .Y(_0731_),
    .A1(_0729_),
    .A2(_0730_));
 sg13g2_nand2b_1 _3200_ (.Y(_0732_),
    .B(_0041_),
    .A_N(net306));
 sg13g2_a21oi_1 _3201_ (.A1(_0724_),
    .A2(_0732_),
    .Y(_0733_),
    .B1(_0726_));
 sg13g2_a21oi_1 _3202_ (.A1(_0040_),
    .A2(_0728_),
    .Y(_0734_),
    .B1(_0733_));
 sg13g2_nand2_1 _3203_ (.Y(_0735_),
    .A(net303),
    .B(_0734_));
 sg13g2_a22oi_1 _3204_ (.Y(_0736_),
    .B1(_0735_),
    .B2(_0720_),
    .A2(_0721_),
    .A1(_0039_));
 sg13g2_nand2_1 _3205_ (.Y(_0737_),
    .A(_0530_),
    .B(_0736_));
 sg13g2_nand3_1 _3206_ (.B(_0731_),
    .C(_0736_),
    .A(_0530_),
    .Y(_0738_));
 sg13g2_inv_1 _3207_ (.Y(_0739_),
    .A(_0738_));
 sg13g2_nand3b_1 _3208_ (.B(_0724_),
    .C(_0038_),
    .Y(_0740_),
    .A_N(net306));
 sg13g2_a21oi_1 _3209_ (.A1(_0072_),
    .A2(_0723_),
    .Y(_0741_),
    .B1(_0726_));
 sg13g2_a22oi_1 _3210_ (.Y(_0742_),
    .B1(_0740_),
    .B2(_0741_),
    .A2(_0728_),
    .A1(\clock_min_u[0] ));
 sg13g2_o21ai_1 _3211_ (.B1(_0720_),
    .Y(_0743_),
    .A1(\clock_min_d[0] ),
    .A2(net303));
 sg13g2_a21oi_1 _3212_ (.A1(net303),
    .A2(_0742_),
    .Y(_0744_),
    .B1(_0743_));
 sg13g2_a21oi_1 _3213_ (.A1(\clock_hrs_u[0] ),
    .A2(_0721_),
    .Y(_0745_),
    .B1(_0744_));
 sg13g2_nor2_1 _3214_ (.A(_0529_),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_a21oi_2 _3215_ (.B1(_0746_),
    .Y(_0747_),
    .A2(_0529_),
    .A1(net508));
 sg13g2_nor2_1 _3216_ (.A(_0739_),
    .B(_0747_),
    .Y(_0000_));
 sg13g2_o21ai_1 _3217_ (.B1(_0724_),
    .Y(_0748_),
    .A1(\clock_sec_u[1] ),
    .A2(net306));
 sg13g2_a21oi_1 _3218_ (.A1(\clock_sec_d[1] ),
    .A2(_0723_),
    .Y(_0749_),
    .B1(_0726_));
 sg13g2_nand2_1 _3219_ (.Y(_0750_),
    .A(\clock_min_u[1] ),
    .B(_0505_));
 sg13g2_a22oi_1 _3220_ (.Y(_0751_),
    .B1(_0750_),
    .B2(_0728_),
    .A2(_0749_),
    .A1(_0748_));
 sg13g2_a21oi_1 _3221_ (.A1(\clock_min_d[1] ),
    .A2(_0504_),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_a221oi_1 _3222_ (.B2(_0720_),
    .C1(_0529_),
    .B1(_0752_),
    .A1(_0048_),
    .Y(_0753_),
    .A2(_0721_));
 sg13g2_inv_1 _3223_ (.Y(_0754_),
    .A(_0753_));
 sg13g2_o21ai_1 _3224_ (.B1(_0754_),
    .Y(_0755_),
    .A1(net543),
    .A2(_0530_));
 sg13g2_and2_1 _3225_ (.A(_0738_),
    .B(_0755_),
    .X(_0001_));
 sg13g2_and2_1 _3226_ (.A(_0731_),
    .B(_0746_),
    .X(_0756_));
 sg13g2_nand3_1 _3227_ (.B(_0731_),
    .C(_0737_),
    .A(_0530_),
    .Y(_0757_));
 sg13g2_a21oi_1 _3228_ (.A1(_0747_),
    .A2(_0757_),
    .Y(_0002_),
    .B1(_0756_));
 sg13g2_xor2_1 _3229_ (.B(_0756_),
    .A(_0755_),
    .X(_0758_));
 sg13g2_nor2_1 _3230_ (.A(_0731_),
    .B(_0737_),
    .Y(_0759_));
 sg13g2_inv_1 _3231_ (.Y(_0760_),
    .A(_0759_));
 sg13g2_nand2_1 _3232_ (.Y(_0761_),
    .A(_0737_),
    .B(_0758_));
 sg13g2_o21ai_1 _3233_ (.B1(_0761_),
    .Y(_0003_),
    .A1(_0758_),
    .A2(_0760_));
 sg13g2_nand2_1 _3234_ (.Y(_0762_),
    .A(_0755_),
    .B(_0759_));
 sg13g2_nor2b_1 _3235_ (.A(_0747_),
    .B_N(_0755_),
    .Y(_0763_));
 sg13g2_o21ai_1 _3236_ (.B1(_0762_),
    .Y(_0004_),
    .A1(_0757_),
    .A2(_0763_));
 sg13g2_nand2b_1 _3237_ (.Y(_0764_),
    .B(_0763_),
    .A_N(_0757_));
 sg13g2_nand2_1 _3238_ (.Y(_0005_),
    .A(_0760_),
    .B(_0764_));
 sg13g2_nor2b_1 _3239_ (.A(net313),
    .B_N(\clock_color_offset[0] ),
    .Y(_0765_));
 sg13g2_xnor2_1 _3240_ (.Y(_0766_),
    .A(\clock_color_offset[0] ),
    .B(net313));
 sg13g2_xor2_1 _3241_ (.B(_1418_),
    .A(net562),
    .X(_0767_));
 sg13g2_and2_1 _3242_ (.A(_0766_),
    .B(_0767_),
    .X(_0768_));
 sg13g2_nand2_1 _3243_ (.Y(_0769_),
    .A(_0766_),
    .B(_0767_));
 sg13g2_xnor2_1 _3244_ (.Y(_0770_),
    .A(_0765_),
    .B(_0767_));
 sg13g2_a22oi_1 _3245_ (.Y(_0771_),
    .B1(_0765_),
    .B2(_0767_),
    .A2(_1418_),
    .A1(_1393_));
 sg13g2_xnor2_1 _3246_ (.Y(_0772_),
    .A(\clock_color_offset[2] ),
    .B(_0500_));
 sg13g2_xnor2_1 _3247_ (.Y(_0773_),
    .A(_0771_),
    .B(_0772_));
 sg13g2_xor2_1 _3248_ (.B(_0772_),
    .A(_0771_),
    .X(_0774_));
 sg13g2_a21oi_1 _3249_ (.A1(_0770_),
    .A2(_0774_),
    .Y(_0006_),
    .B1(_0768_));
 sg13g2_nor2_1 _3250_ (.A(_0766_),
    .B(_0773_),
    .Y(_0775_));
 sg13g2_a21oi_1 _3251_ (.A1(_0768_),
    .A2(_0773_),
    .Y(_0007_),
    .B1(_0775_));
 sg13g2_nand2b_1 _3252_ (.Y(_0776_),
    .B(_0770_),
    .A_N(_0766_));
 sg13g2_a21oi_1 _3253_ (.A1(_0769_),
    .A2(_0776_),
    .Y(_0079_),
    .B1(_0773_));
 sg13g2_nor2_1 _3254_ (.A(_0768_),
    .B(_0773_),
    .Y(_0080_));
 sg13g2_nor2_2 _3255_ (.A(_1421_),
    .B(_1434_),
    .Y(_0777_));
 sg13g2_nand2_2 _3256_ (.Y(_0778_),
    .A(hmax),
    .B(\vga_sync.o_vmax ));
 sg13g2_nand4_1 _3257_ (.B(_1415_),
    .C(_1418_),
    .A(_1413_),
    .Y(_0779_),
    .D(_1420_));
 sg13g2_nor2_2 _3258_ (.A(_1434_),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_or2_1 _3259_ (.X(_0781_),
    .B(_0779_),
    .A(_1434_));
 sg13g2_a21oi_1 _3260_ (.A1(\ydelta[0] ),
    .A2(net300),
    .Y(_0782_),
    .B1(net360));
 sg13g2_nor3_2 _3261_ (.A(\ydelta[2] ),
    .B(\ydelta[1] ),
    .C(\ydelta[0] ),
    .Y(_0783_));
 sg13g2_nor2b_1 _3262_ (.A(\ydelta[3] ),
    .B_N(_0783_),
    .Y(_0784_));
 sg13g2_and2_1 _3263_ (.A(_1388_),
    .B(_0784_),
    .X(_0785_));
 sg13g2_nor2b_1 _3264_ (.A(\ydelta[5] ),
    .B_N(_0785_),
    .Y(_0786_));
 sg13g2_nor2b_2 _3265_ (.A(\ydelta[6] ),
    .B_N(_0786_),
    .Y(_0787_));
 sg13g2_o21ai_1 _3266_ (.B1(_0064_),
    .Y(_0788_),
    .A1(_1387_),
    .A2(_0787_));
 sg13g2_xnor2_1 _3267_ (.Y(_0789_),
    .A(\ydelta[6] ),
    .B(_0786_));
 sg13g2_xnor2_1 _3268_ (.Y(_0790_),
    .A(\ydelta[5] ),
    .B(_0785_));
 sg13g2_nand2b_1 _3269_ (.Y(_0791_),
    .B(_0790_),
    .A_N(\py[5] ));
 sg13g2_xnor2_1 _3270_ (.Y(_0792_),
    .A(\ydelta[3] ),
    .B(_0783_));
 sg13g2_nor2b_1 _3271_ (.A(net345),
    .B_N(_0792_),
    .Y(_0793_));
 sg13g2_nand2b_1 _3272_ (.Y(_0794_),
    .B(net345),
    .A_N(_0792_));
 sg13g2_o21ai_1 _3273_ (.B1(\ydelta[2] ),
    .Y(_0795_),
    .A1(\ydelta[1] ),
    .A2(\ydelta[0] ));
 sg13g2_nor2b_1 _3274_ (.A(_0783_),
    .B_N(_0795_),
    .Y(_0796_));
 sg13g2_nor2b_1 _3275_ (.A(\py[2] ),
    .B_N(_0796_),
    .Y(_0797_));
 sg13g2_a21oi_1 _3276_ (.A1(_0794_),
    .A2(_0797_),
    .Y(_0798_),
    .B1(_0793_));
 sg13g2_xor2_1 _3277_ (.B(\ydelta[0] ),
    .A(\ydelta[1] ),
    .X(_0799_));
 sg13g2_nor2b_1 _3278_ (.A(\ydelta[0] ),
    .B_N(net348),
    .Y(_0800_));
 sg13g2_nor3_1 _3279_ (.A(_1396_),
    .B(_0799_),
    .C(_0800_),
    .Y(_0801_));
 sg13g2_o21ai_1 _3280_ (.B1(net346),
    .Y(_0802_),
    .A1(_0063_),
    .A2(_0800_));
 sg13g2_a21o_1 _3281_ (.A2(_0802_),
    .A1(_0799_),
    .B1(_0801_),
    .X(_0803_));
 sg13g2_xor2_1 _3282_ (.B(_0796_),
    .A(_0062_),
    .X(_0804_));
 sg13g2_nand3_1 _3283_ (.B(_0803_),
    .C(_0804_),
    .A(_0794_),
    .Y(_0805_));
 sg13g2_xnor2_1 _3284_ (.Y(_0806_),
    .A(net475),
    .B(_0784_));
 sg13g2_nand2_1 _3285_ (.Y(_0807_),
    .A(_0061_),
    .B(_0806_));
 sg13g2_nand3_1 _3286_ (.B(_0805_),
    .C(_0807_),
    .A(_0798_),
    .Y(_0808_));
 sg13g2_xnor2_1 _3287_ (.Y(_0809_),
    .A(_0060_),
    .B(_0790_));
 sg13g2_o21ai_1 _3288_ (.B1(_0808_),
    .Y(_0810_),
    .A1(_0061_),
    .A2(_0806_));
 sg13g2_o21ai_1 _3289_ (.B1(_0791_),
    .Y(_0811_),
    .A1(_0809_),
    .A2(_0810_));
 sg13g2_xor2_1 _3290_ (.B(_0789_),
    .A(_0059_),
    .X(_0812_));
 sg13g2_a22oi_1 _3291_ (.Y(_0813_),
    .B1(_0811_),
    .B2(_0812_),
    .A2(_0789_),
    .A1(_1382_));
 sg13g2_nor2_1 _3292_ (.A(\py[7] ),
    .B(net355),
    .Y(_0814_));
 sg13g2_xor2_1 _3293_ (.B(net355),
    .A(\py[7] ),
    .X(_0815_));
 sg13g2_xnor2_1 _3294_ (.Y(_0816_),
    .A(_0787_),
    .B(_0815_));
 sg13g2_o21ai_1 _3295_ (.B1(_0788_),
    .Y(_0817_),
    .A1(_0813_),
    .A2(_0816_));
 sg13g2_nor2_1 _3296_ (.A(\pym[11] ),
    .B(\pym[10] ),
    .Y(_0818_));
 sg13g2_nor3_1 _3297_ (.A(\py[9] ),
    .B(\py[8] ),
    .C(_0058_),
    .Y(_0819_));
 sg13g2_nand3_1 _3298_ (.B(_0818_),
    .C(_0819_),
    .A(_0817_),
    .Y(_0820_));
 sg13g2_a21oi_2 _3299_ (.B1(_0820_),
    .Y(_0821_),
    .A2(_0787_),
    .A1(_1387_));
 sg13g2_nor2b_1 _3300_ (.A(_0050_),
    .B_N(net286),
    .Y(_0822_));
 sg13g2_o21ai_1 _3301_ (.B1(_0777_),
    .Y(_0823_),
    .A1(net268),
    .A2(net286));
 sg13g2_o21ai_1 _3302_ (.B1(_0782_),
    .Y(_0081_),
    .A1(_0822_),
    .A2(_0823_));
 sg13g2_nor2_2 _3303_ (.A(net358),
    .B(net301),
    .Y(_0824_));
 sg13g2_nand2_2 _3304_ (.Y(_0825_),
    .A(net364),
    .B(net300));
 sg13g2_nand2_1 _3305_ (.Y(_0826_),
    .A(net481),
    .B(net293));
 sg13g2_nor2_2 _3306_ (.A(net357),
    .B(_0778_),
    .Y(_0827_));
 sg13g2_nand2_1 _3307_ (.Y(_0828_),
    .A(net364),
    .B(_0777_));
 sg13g2_nand2b_1 _3308_ (.Y(_0829_),
    .B(_0827_),
    .A_N(net286));
 sg13g2_nor2_1 _3309_ (.A(\px[1] ),
    .B(\px[0] ),
    .Y(_0830_));
 sg13g2_xnor2_1 _3310_ (.Y(_0831_),
    .A(net353),
    .B(net354));
 sg13g2_nor3_2 _3311_ (.A(net360),
    .B(net300),
    .C(net286),
    .Y(_0832_));
 sg13g2_mux2_1 _3312_ (.A0(_0799_),
    .A1(_0831_),
    .S(net286),
    .X(_0833_));
 sg13g2_o21ai_1 _3313_ (.B1(_0826_),
    .Y(_0082_),
    .A1(net289),
    .A2(_0833_));
 sg13g2_a21o_1 _3314_ (.A2(net354),
    .A1(net353),
    .B1(\px[2] ),
    .X(_0834_));
 sg13g2_nand4_1 _3315_ (.B(net353),
    .C(net354),
    .A(\px[2] ),
    .Y(_0835_),
    .D(_0827_));
 sg13g2_and2_1 _3316_ (.A(net285),
    .B(_0835_),
    .X(_0836_));
 sg13g2_o21ai_1 _3317_ (.B1(_0836_),
    .Y(_0837_),
    .A1(net289),
    .A2(_0834_));
 sg13g2_o21ai_1 _3318_ (.B1(_0837_),
    .Y(_0838_),
    .A1(_0796_),
    .A2(net286));
 sg13g2_o21ai_1 _3319_ (.B1(_0838_),
    .Y(_0839_),
    .A1(net531),
    .A2(_0825_));
 sg13g2_inv_1 _3320_ (.Y(_0083_),
    .A(_0839_));
 sg13g2_nand2_1 _3321_ (.Y(_0840_),
    .A(net381),
    .B(net291));
 sg13g2_nor2b_1 _3322_ (.A(net286),
    .B_N(_0792_),
    .Y(_0841_));
 sg13g2_o21ai_1 _3323_ (.B1(_0840_),
    .Y(_0084_),
    .A1(_0836_),
    .A2(_0841_));
 sg13g2_a22oi_1 _3324_ (.Y(_0085_),
    .B1(_0832_),
    .B2(_0806_),
    .A2(net291),
    .A1(_1388_));
 sg13g2_nand2_1 _3325_ (.Y(_0842_),
    .A(net446),
    .B(net290));
 sg13g2_o21ai_1 _3326_ (.B1(_0842_),
    .Y(_0086_),
    .A1(_0790_),
    .A2(net284));
 sg13g2_nand2_1 _3327_ (.Y(_0843_),
    .A(net441),
    .B(net290));
 sg13g2_o21ai_1 _3328_ (.B1(_0843_),
    .Y(_0087_),
    .A1(_0789_),
    .A2(net284));
 sg13g2_nand2_1 _3329_ (.Y(_0844_),
    .A(net355),
    .B(net290));
 sg13g2_xor2_1 _3330_ (.B(_0787_),
    .A(net407),
    .X(_0845_));
 sg13g2_o21ai_1 _3331_ (.B1(_0844_),
    .Y(_0088_),
    .A1(net284),
    .A2(_0845_));
 sg13g2_a22oi_1 _3332_ (.Y(_0846_),
    .B1(_0827_),
    .B2(net233),
    .A2(net293),
    .A1(\pxm[0] ));
 sg13g2_inv_1 _3333_ (.Y(_0089_),
    .A(net234));
 sg13g2_nand2_1 _3334_ (.Y(_0847_),
    .A(net245),
    .B(net293));
 sg13g2_nor2b_1 _3335_ (.A(net342),
    .B_N(\pxm[1] ),
    .Y(_0848_));
 sg13g2_nand2b_1 _3336_ (.Y(_0849_),
    .B(net342),
    .A_N(\pxm[1] ));
 sg13g2_nand2b_1 _3337_ (.Y(_0850_),
    .B(_0849_),
    .A_N(_0848_));
 sg13g2_xnor2_1 _3338_ (.Y(_0851_),
    .A(net233),
    .B(_0850_));
 sg13g2_o21ai_1 _3339_ (.B1(_0847_),
    .Y(_0090_),
    .A1(net289),
    .A2(_0851_));
 sg13g2_nand2_1 _3340_ (.Y(_0852_),
    .A(net354),
    .B(net293));
 sg13g2_xor2_1 _3341_ (.B(net354),
    .A(net342),
    .X(_0853_));
 sg13g2_o21ai_1 _3342_ (.B1(_0849_),
    .Y(_0854_),
    .A1(net557),
    .A2(_0848_));
 sg13g2_or2_1 _3343_ (.X(_0855_),
    .B(_0854_),
    .A(_0853_));
 sg13g2_xnor2_1 _3344_ (.Y(_0856_),
    .A(_0853_),
    .B(_0854_));
 sg13g2_o21ai_1 _3345_ (.B1(_0852_),
    .Y(_0091_),
    .A1(net289),
    .A2(_0856_));
 sg13g2_nand2_1 _3346_ (.Y(_0857_),
    .A(net353),
    .B(net293));
 sg13g2_xor2_1 _3347_ (.B(net353),
    .A(net342),
    .X(_0858_));
 sg13g2_o21ai_1 _3348_ (.B1(_0855_),
    .Y(_0859_),
    .A1(net342),
    .A2(_1386_));
 sg13g2_xnor2_1 _3349_ (.Y(_0860_),
    .A(_0858_),
    .B(_0859_));
 sg13g2_o21ai_1 _3350_ (.B1(_0857_),
    .Y(_0092_),
    .A1(net289),
    .A2(_0860_));
 sg13g2_nand2_1 _3351_ (.Y(_0861_),
    .A(net521),
    .B(net293));
 sg13g2_xor2_1 _3352_ (.B(\px[2] ),
    .A(net342),
    .X(_0862_));
 sg13g2_o21ai_1 _3353_ (.B1(net353),
    .Y(_0863_),
    .A1(net342),
    .A2(net354));
 sg13g2_nand2_1 _3354_ (.Y(_0864_),
    .A(_0855_),
    .B(_0863_));
 sg13g2_o21ai_1 _3355_ (.B1(_0864_),
    .Y(_0865_),
    .A1(net342),
    .A2(net353));
 sg13g2_or2_1 _3356_ (.X(_0866_),
    .B(_0865_),
    .A(_0862_));
 sg13g2_xnor2_1 _3357_ (.Y(_0867_),
    .A(_0862_),
    .B(_0865_));
 sg13g2_o21ai_1 _3358_ (.B1(_0861_),
    .Y(_0093_),
    .A1(net289),
    .A2(_0867_));
 sg13g2_nand2_1 _3359_ (.Y(_0868_),
    .A(net422),
    .B(net294));
 sg13g2_o21ai_1 _3360_ (.B1(_0866_),
    .Y(_0869_),
    .A1(net343),
    .A2(_1385_));
 sg13g2_xnor2_1 _3361_ (.Y(_0870_),
    .A(net343),
    .B(\px[3] ));
 sg13g2_xnor2_1 _3362_ (.Y(_0871_),
    .A(_0869_),
    .B(_0870_));
 sg13g2_o21ai_1 _3363_ (.B1(_0868_),
    .Y(_0094_),
    .A1(net289),
    .A2(_0871_));
 sg13g2_nand2_1 _3364_ (.Y(_0872_),
    .A(net491),
    .B(net294));
 sg13g2_xor2_1 _3365_ (.B(\px[4] ),
    .A(dx),
    .X(_0873_));
 sg13g2_nand2b_2 _3366_ (.Y(_0874_),
    .B(_0870_),
    .A_N(_0866_));
 sg13g2_nor2_1 _3367_ (.A(\px[3] ),
    .B(\px[2] ),
    .Y(_0875_));
 sg13g2_or2_1 _3368_ (.X(_0876_),
    .B(_0875_),
    .A(dx));
 sg13g2_nand3_1 _3369_ (.B(_0874_),
    .C(_0876_),
    .A(_0873_),
    .Y(_0877_));
 sg13g2_a21oi_1 _3370_ (.A1(_0874_),
    .A2(_0876_),
    .Y(_0878_),
    .B1(_0873_));
 sg13g2_nand2_1 _3371_ (.Y(_0879_),
    .A(_0827_),
    .B(_0877_));
 sg13g2_o21ai_1 _3372_ (.B1(_0872_),
    .Y(_0095_),
    .A1(_0878_),
    .A2(_0879_));
 sg13g2_nand2_1 _3373_ (.Y(_0880_),
    .A(net267),
    .B(net297));
 sg13g2_xor2_1 _3374_ (.B(net352),
    .A(net343),
    .X(_0881_));
 sg13g2_a21oi_1 _3375_ (.A1(_1375_),
    .A2(\px[4] ),
    .Y(_0882_),
    .B1(_0878_));
 sg13g2_xnor2_1 _3376_ (.Y(_0883_),
    .A(_0881_),
    .B(_0882_));
 sg13g2_o21ai_1 _3377_ (.B1(_0880_),
    .Y(_0096_),
    .A1(_0828_),
    .A2(_0883_));
 sg13g2_nand2_1 _3378_ (.Y(_0884_),
    .A(net263),
    .B(net297));
 sg13g2_xor2_1 _3379_ (.B(\px[6] ),
    .A(net343),
    .X(_0885_));
 sg13g2_nor3_1 _3380_ (.A(_0873_),
    .B(_0874_),
    .C(_0881_),
    .Y(_0886_));
 sg13g2_o21ai_1 _3381_ (.B1(_1375_),
    .Y(_0887_),
    .A1(\px[5] ),
    .A2(\px[4] ));
 sg13g2_nand2_1 _3382_ (.Y(_0888_),
    .A(_0876_),
    .B(_0887_));
 sg13g2_nor2_1 _3383_ (.A(_0886_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_nor2_1 _3384_ (.A(_0885_),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_a21o_1 _3385_ (.A2(_0889_),
    .A1(_0885_),
    .B1(net289),
    .X(_0891_));
 sg13g2_o21ai_1 _3386_ (.B1(_0884_),
    .Y(_0097_),
    .A1(_0890_),
    .A2(_0891_));
 sg13g2_nand2_1 _3387_ (.Y(_0892_),
    .A(net237),
    .B(net297));
 sg13g2_xor2_1 _3388_ (.B(net350),
    .A(net343),
    .X(_0893_));
 sg13g2_a21oi_1 _3389_ (.A1(_1375_),
    .A2(net351),
    .Y(_0894_),
    .B1(_0890_));
 sg13g2_xnor2_1 _3390_ (.Y(_0895_),
    .A(_0893_),
    .B(_0894_));
 sg13g2_o21ai_1 _3391_ (.B1(_0892_),
    .Y(_0098_),
    .A1(_0828_),
    .A2(_0895_));
 sg13g2_o21ai_1 _3392_ (.B1(_0890_),
    .Y(_0896_),
    .A1(_1375_),
    .A2(net350));
 sg13g2_o21ai_1 _3393_ (.B1(_1375_),
    .Y(_0897_),
    .A1(net350),
    .A2(net351));
 sg13g2_and2_1 _3394_ (.A(_0896_),
    .B(_0897_),
    .X(_0898_));
 sg13g2_xor2_1 _3395_ (.B(net547),
    .A(net343),
    .X(_0899_));
 sg13g2_o21ai_1 _3396_ (.B1(_0827_),
    .Y(_0900_),
    .A1(_0898_),
    .A2(_0899_));
 sg13g2_a21oi_1 _3397_ (.A1(_0898_),
    .A2(_0899_),
    .Y(_0901_),
    .B1(_0900_));
 sg13g2_a21o_1 _3398_ (.A2(net297),
    .A1(net349),
    .B1(_0901_),
    .X(_0099_));
 sg13g2_nor2_1 _3399_ (.A(net349),
    .B(_0898_),
    .Y(_0902_));
 sg13g2_a21oi_1 _3400_ (.A1(_1375_),
    .A2(net349),
    .Y(_0903_),
    .B1(_0778_));
 sg13g2_a21oi_1 _3401_ (.A1(net343),
    .A2(_0896_),
    .Y(_0904_),
    .B1(_0902_));
 sg13g2_and2_1 _3402_ (.A(_0903_),
    .B(_0904_),
    .X(_0905_));
 sg13g2_o21ai_1 _3403_ (.B1(net364),
    .Y(_0906_),
    .A1(net490),
    .A2(_0905_));
 sg13g2_a21oi_1 _3404_ (.A1(net490),
    .A2(_0905_),
    .Y(_0100_),
    .B1(_0906_));
 sg13g2_nand2_1 _3405_ (.Y(_0907_),
    .A(net348),
    .B(net293));
 sg13g2_nand2_1 _3406_ (.Y(_0908_),
    .A(net348),
    .B(\ydelta[0] ));
 sg13g2_xnor2_1 _3407_ (.Y(_0909_),
    .A(net348),
    .B(net500));
 sg13g2_o21ai_1 _3408_ (.B1(_0907_),
    .Y(_0101_),
    .A1(net285),
    .A2(net501));
 sg13g2_nand2_1 _3409_ (.Y(_0910_),
    .A(net346),
    .B(net291));
 sg13g2_nand2_1 _3410_ (.Y(_0911_),
    .A(net346),
    .B(\ydelta[1] ));
 sg13g2_xnor2_1 _3411_ (.Y(_0912_),
    .A(net346),
    .B(\ydelta[1] ));
 sg13g2_xnor2_1 _3412_ (.Y(_0913_),
    .A(_0908_),
    .B(_0912_));
 sg13g2_o21ai_1 _3413_ (.B1(_0910_),
    .Y(_0102_),
    .A1(net285),
    .A2(_0913_));
 sg13g2_nand2_1 _3414_ (.Y(_0914_),
    .A(net541),
    .B(net291));
 sg13g2_o21ai_1 _3415_ (.B1(_0911_),
    .Y(_0915_),
    .A1(_0908_),
    .A2(_0912_));
 sg13g2_and2_1 _3416_ (.A(\py[2] ),
    .B(\ydelta[2] ),
    .X(_0916_));
 sg13g2_xor2_1 _3417_ (.B(\ydelta[2] ),
    .A(\py[2] ),
    .X(_0917_));
 sg13g2_xnor2_1 _3418_ (.Y(_0918_),
    .A(_0915_),
    .B(_0917_));
 sg13g2_o21ai_1 _3419_ (.B1(_0914_),
    .Y(_0103_),
    .A1(net285),
    .A2(_0918_));
 sg13g2_nand2_1 _3420_ (.Y(_0919_),
    .A(net345),
    .B(net292));
 sg13g2_a21oi_1 _3421_ (.A1(_0915_),
    .A2(_0917_),
    .Y(_0920_),
    .B1(_0916_));
 sg13g2_and2_1 _3422_ (.A(net345),
    .B(\ydelta[3] ),
    .X(_0921_));
 sg13g2_or2_1 _3423_ (.X(_0922_),
    .B(\ydelta[3] ),
    .A(net345));
 sg13g2_nand2b_1 _3424_ (.Y(_0923_),
    .B(_0922_),
    .A_N(_0921_));
 sg13g2_xnor2_1 _3425_ (.Y(_0924_),
    .A(_0920_),
    .B(_0923_));
 sg13g2_o21ai_1 _3426_ (.B1(_0919_),
    .Y(_0104_),
    .A1(net285),
    .A2(_0924_));
 sg13g2_nand2_1 _3427_ (.Y(_0925_),
    .A(\py[4] ),
    .B(\ydelta[4] ));
 sg13g2_xor2_1 _3428_ (.B(\ydelta[4] ),
    .A(\py[4] ),
    .X(_0926_));
 sg13g2_a221oi_1 _3429_ (.B2(_0922_),
    .C1(_0921_),
    .B1(_0916_),
    .A1(_0798_),
    .Y(_0927_),
    .A2(_0915_));
 sg13g2_nand2b_1 _3430_ (.Y(_0928_),
    .B(_0926_),
    .A_N(_0927_));
 sg13g2_xnor2_1 _3431_ (.Y(_0929_),
    .A(_0926_),
    .B(_0927_));
 sg13g2_nand2_1 _3432_ (.Y(_0930_),
    .A(_0832_),
    .B(_0929_));
 sg13g2_o21ai_1 _3433_ (.B1(_0930_),
    .Y(_0105_),
    .A1(_1383_),
    .A2(_0825_));
 sg13g2_nand2_1 _3434_ (.Y(_0931_),
    .A(net503),
    .B(net290));
 sg13g2_nand2_1 _3435_ (.Y(_0932_),
    .A(_0925_),
    .B(_0928_));
 sg13g2_nor2_1 _3436_ (.A(\py[5] ),
    .B(\ydelta[5] ),
    .Y(_0933_));
 sg13g2_a21oi_1 _3437_ (.A1(_0925_),
    .A2(_0928_),
    .Y(_0934_),
    .B1(_0933_));
 sg13g2_xor2_1 _3438_ (.B(\ydelta[5] ),
    .A(\py[5] ),
    .X(_0935_));
 sg13g2_xnor2_1 _3439_ (.Y(_0936_),
    .A(_0932_),
    .B(_0935_));
 sg13g2_o21ai_1 _3440_ (.B1(_0931_),
    .Y(_0106_),
    .A1(net284),
    .A2(_0936_));
 sg13g2_nand2_1 _3441_ (.Y(_0937_),
    .A(net453),
    .B(net292));
 sg13g2_nand2_1 _3442_ (.Y(_0938_),
    .A(\py[6] ),
    .B(\ydelta[6] ));
 sg13g2_xnor2_1 _3443_ (.Y(_0939_),
    .A(\py[6] ),
    .B(\ydelta[6] ));
 sg13g2_a21oi_1 _3444_ (.A1(\py[5] ),
    .A2(\ydelta[5] ),
    .Y(_0940_),
    .B1(_0934_));
 sg13g2_xnor2_1 _3445_ (.Y(_0941_),
    .A(_0939_),
    .B(_0940_));
 sg13g2_o21ai_1 _3446_ (.B1(_0937_),
    .Y(_0107_),
    .A1(net285),
    .A2(_0941_));
 sg13g2_nand2_1 _3447_ (.Y(_0942_),
    .A(net447),
    .B(net290));
 sg13g2_o21ai_1 _3448_ (.B1(_0938_),
    .Y(_0943_),
    .A1(_0939_),
    .A2(_0940_));
 sg13g2_xnor2_1 _3449_ (.Y(_0944_),
    .A(_0815_),
    .B(_0943_));
 sg13g2_o21ai_1 _3450_ (.B1(_0942_),
    .Y(_0108_),
    .A1(net284),
    .A2(_0944_));
 sg13g2_xnor2_1 _3451_ (.Y(_0945_),
    .A(\py[8] ),
    .B(net356));
 sg13g2_a21oi_1 _3452_ (.A1(\py[7] ),
    .A2(net355),
    .Y(_0946_),
    .B1(_0943_));
 sg13g2_o21ai_1 _3453_ (.B1(_0945_),
    .Y(_0947_),
    .A1(_0814_),
    .A2(_0946_));
 sg13g2_nor3_1 _3454_ (.A(_0814_),
    .B(_0945_),
    .C(_0946_),
    .Y(_0948_));
 sg13g2_nor2_1 _3455_ (.A(net284),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_a22oi_1 _3456_ (.Y(_0950_),
    .B1(_0947_),
    .B2(_0949_),
    .A2(net290),
    .A1(net528));
 sg13g2_inv_1 _3457_ (.Y(_0109_),
    .A(_0950_));
 sg13g2_a21oi_1 _3458_ (.A1(\py[8] ),
    .A2(net356),
    .Y(_0951_),
    .B1(_0948_));
 sg13g2_nand2_1 _3459_ (.Y(_0952_),
    .A(\py[9] ),
    .B(net356));
 sg13g2_nor2_1 _3460_ (.A(\py[9] ),
    .B(net356),
    .Y(_0953_));
 sg13g2_xnor2_1 _3461_ (.Y(_0954_),
    .A(\py[9] ),
    .B(net355));
 sg13g2_a21oi_1 _3462_ (.A1(_0951_),
    .A2(_0954_),
    .Y(_0955_),
    .B1(net284));
 sg13g2_o21ai_1 _3463_ (.B1(_0955_),
    .Y(_0956_),
    .A1(_0951_),
    .A2(_0954_));
 sg13g2_o21ai_1 _3464_ (.B1(_0956_),
    .Y(_0110_),
    .A1(_1381_),
    .A2(_0825_));
 sg13g2_xor2_1 _3465_ (.B(net355),
    .A(\pym[10] ),
    .X(_0957_));
 sg13g2_o21ai_1 _3466_ (.B1(_0952_),
    .Y(_0958_),
    .A1(_0951_),
    .A2(_0953_));
 sg13g2_nand2_1 _3467_ (.Y(_0959_),
    .A(_0957_),
    .B(_0958_));
 sg13g2_nor2_1 _3468_ (.A(_0957_),
    .B(_0958_),
    .Y(_0960_));
 sg13g2_nor2_1 _3469_ (.A(net284),
    .B(_0960_),
    .Y(_0961_));
 sg13g2_a22oi_1 _3470_ (.Y(_0962_),
    .B1(_0959_),
    .B2(_0961_),
    .A2(net290),
    .A1(net396));
 sg13g2_inv_1 _3471_ (.Y(_0111_),
    .A(_0962_));
 sg13g2_o21ai_1 _3472_ (.B1(_0959_),
    .Y(_0963_),
    .A1(_1380_),
    .A2(_1387_));
 sg13g2_xnor2_1 _3473_ (.Y(_0964_),
    .A(net377),
    .B(net355));
 sg13g2_xnor2_1 _3474_ (.Y(_0965_),
    .A(_0963_),
    .B(_0964_));
 sg13g2_a22oi_1 _3475_ (.Y(_0966_),
    .B1(_0832_),
    .B2(_0965_),
    .A2(net290),
    .A1(net377));
 sg13g2_inv_1 _3476_ (.Y(_0112_),
    .A(_0966_));
 sg13g2_a22oi_1 _3477_ (.Y(_0967_),
    .B1(_0827_),
    .B2(net226),
    .A2(net297),
    .A1(\t[0] ));
 sg13g2_inv_1 _3478_ (.Y(_0113_),
    .A(net227));
 sg13g2_a21oi_1 _3479_ (.A1(net463),
    .A2(net302),
    .Y(_0968_),
    .B1(\t[1] ));
 sg13g2_nand3_1 _3480_ (.B(\t[0] ),
    .C(net302),
    .A(\t[1] ),
    .Y(_0969_));
 sg13g2_nand2_1 _3481_ (.Y(_0970_),
    .A(net367),
    .B(_0969_));
 sg13g2_nor2_1 _3482_ (.A(net464),
    .B(_0970_),
    .Y(_0114_));
 sg13g2_or2_1 _3483_ (.X(_0971_),
    .B(_0969_),
    .A(_1379_));
 sg13g2_nand2_1 _3484_ (.Y(_0972_),
    .A(net367),
    .B(_0971_));
 sg13g2_a21oi_1 _3485_ (.A1(_1379_),
    .A2(_0969_),
    .Y(_0115_),
    .B1(_0972_));
 sg13g2_o21ai_1 _3486_ (.B1(net367),
    .Y(_0973_),
    .A1(_1378_),
    .A2(_0971_));
 sg13g2_a21oi_1 _3487_ (.A1(_1378_),
    .A2(_0971_),
    .Y(_0116_),
    .B1(_0973_));
 sg13g2_nor2_1 _3488_ (.A(net349),
    .B(net350),
    .Y(_0974_));
 sg13g2_nor4_1 _3489_ (.A(\px[9] ),
    .B(net351),
    .C(\px[5] ),
    .D(\px[4] ),
    .Y(_0975_));
 sg13g2_nand4_1 _3490_ (.B(_0875_),
    .C(_0974_),
    .A(_0830_),
    .Y(_0976_),
    .D(_0975_));
 sg13g2_nand2_1 _3491_ (.Y(_0977_),
    .A(_0362_),
    .B(_0974_));
 sg13g2_nand2_1 _3492_ (.Y(_0978_),
    .A(\px[9] ),
    .B(_0977_));
 sg13g2_nand2_2 _3493_ (.Y(_0979_),
    .A(_0976_),
    .B(_0978_));
 sg13g2_nor2_1 _3494_ (.A(_0821_),
    .B(_0979_),
    .Y(_0980_));
 sg13g2_nor2_1 _3495_ (.A(_1397_),
    .B(_0432_),
    .Y(_0981_));
 sg13g2_and2_1 _3496_ (.A(\product_comp[2] ),
    .B(\product_comp[1] ),
    .X(_0982_));
 sg13g2_nand3b_1 _3497_ (.B(_0438_),
    .C(_0478_),
    .Y(_0983_),
    .A_N(\product_comp[7] ));
 sg13g2_nor4_1 _3498_ (.A(\product_comp[3] ),
    .B(_0981_),
    .C(_0982_),
    .D(_0983_),
    .Y(_0984_));
 sg13g2_nor4_2 _3499_ (.A(_0778_),
    .B(net286),
    .C(_0979_),
    .Y(_0985_),
    .D(_0984_));
 sg13g2_nor4_1 _3500_ (.A(net344),
    .B(\product_comp[3] ),
    .C(_0981_),
    .D(_0982_),
    .Y(_0986_));
 sg13g2_nand4_1 _3501_ (.B(_0478_),
    .C(_0980_),
    .A(_0438_),
    .Y(_0987_),
    .D(_0986_));
 sg13g2_and2_2 _3502_ (.A(_0780_),
    .B(_0987_),
    .X(_0988_));
 sg13g2_inv_1 _3503_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_o21ai_1 _3504_ (.B1(net368),
    .Y(_0990_),
    .A1(net489),
    .A2(net283));
 sg13g2_a21oi_1 _3505_ (.A1(net489),
    .A2(_0988_),
    .Y(_0117_),
    .B1(_0990_));
 sg13g2_o21ai_1 _3506_ (.B1(net283),
    .Y(_0991_),
    .A1(_0431_),
    .A2(_0458_));
 sg13g2_nand2_1 _3507_ (.Y(_0992_),
    .A(net514),
    .B(_0989_));
 sg13g2_nand3_1 _3508_ (.B(_0991_),
    .C(_0992_),
    .A(net368),
    .Y(_0118_));
 sg13g2_nand2_1 _3509_ (.Y(_0993_),
    .A(_0432_),
    .B(_0439_));
 sg13g2_o21ai_1 _3510_ (.B1(net368),
    .Y(_0994_),
    .A1(net523),
    .A2(_0988_));
 sg13g2_a21oi_1 _3511_ (.A1(net283),
    .A2(_0993_),
    .Y(_0119_),
    .B1(_0994_));
 sg13g2_nand3_1 _3512_ (.B(_0477_),
    .C(net283),
    .A(_0433_),
    .Y(_0995_));
 sg13g2_o21ai_1 _3513_ (.B1(_0995_),
    .Y(_0996_),
    .A1(net549),
    .A2(_0988_));
 sg13g2_nand2_1 _3514_ (.Y(_0120_),
    .A(net368),
    .B(_0996_));
 sg13g2_xnor2_1 _3515_ (.Y(_0997_),
    .A(net485),
    .B(_0433_));
 sg13g2_o21ai_1 _3516_ (.B1(net368),
    .Y(_0998_),
    .A1(\product_comp[4] ),
    .A2(_0988_));
 sg13g2_a21oi_1 _3517_ (.A1(_0985_),
    .A2(_0997_),
    .Y(_0121_),
    .B1(_0998_));
 sg13g2_nor2_1 _3518_ (.A(\product_comp[4] ),
    .B(_0433_),
    .Y(_0999_));
 sg13g2_xnor2_1 _3519_ (.Y(_1000_),
    .A(net429),
    .B(_0999_));
 sg13g2_a22oi_1 _3520_ (.Y(_1001_),
    .B1(net283),
    .B2(_1000_),
    .A2(net300),
    .A1(\product_comp[5] ));
 sg13g2_nor2_1 _3521_ (.A(net357),
    .B(net430),
    .Y(_0122_));
 sg13g2_nor3_1 _3522_ (.A(\product_comp[5] ),
    .B(\product_comp[4] ),
    .C(_0433_),
    .Y(_1002_));
 sg13g2_xor2_1 _3523_ (.B(_1002_),
    .A(net439),
    .X(_1003_));
 sg13g2_o21ai_1 _3524_ (.B1(net367),
    .Y(_1004_),
    .A1(\product_comp[6] ),
    .A2(_0988_));
 sg13g2_a21oi_1 _3525_ (.A1(net283),
    .A2(_1003_),
    .Y(_0123_),
    .B1(_1004_));
 sg13g2_nand3_1 _3526_ (.B(_0432_),
    .C(_0478_),
    .A(_1377_),
    .Y(_1005_));
 sg13g2_or2_1 _3527_ (.X(_1006_),
    .B(_1005_),
    .A(net344));
 sg13g2_xor2_1 _3528_ (.B(_1005_),
    .A(net344),
    .X(_1007_));
 sg13g2_o21ai_1 _3529_ (.B1(net367),
    .Y(_1008_),
    .A1(net344),
    .A2(_0988_));
 sg13g2_a21oi_1 _3530_ (.A1(_0985_),
    .A2(_1007_),
    .Y(_0124_),
    .B1(_1008_));
 sg13g2_xor2_1 _3531_ (.B(_1006_),
    .A(net437),
    .X(_1009_));
 sg13g2_a22oi_1 _3532_ (.Y(_1010_),
    .B1(_1009_),
    .B2(net283),
    .A2(_0989_),
    .A1(\product_comp[8] ));
 sg13g2_nor2_1 _3533_ (.A(net357),
    .B(net438),
    .Y(_0125_));
 sg13g2_nor2_1 _3534_ (.A(\product_comp[8] ),
    .B(_1006_),
    .Y(_1011_));
 sg13g2_xnor2_1 _3535_ (.Y(_1012_),
    .A(net435),
    .B(_1011_));
 sg13g2_a22oi_1 _3536_ (.Y(_1013_),
    .B1(_1012_),
    .B2(net283),
    .A2(_0989_),
    .A1(\product_comp[9] ));
 sg13g2_nor2_1 _3537_ (.A(net357),
    .B(net436),
    .Y(_0126_));
 sg13g2_nor3_1 _3538_ (.A(\product_comp[9] ),
    .B(\product_comp[8] ),
    .C(_1006_),
    .Y(_1014_));
 sg13g2_xnor2_1 _3539_ (.Y(_1015_),
    .A(_0065_),
    .B(_1014_));
 sg13g2_a22oi_1 _3540_ (.Y(_1016_),
    .B1(_1015_),
    .B2(_0985_),
    .A2(_0989_),
    .A1(net388));
 sg13g2_nor2_1 _3541_ (.A(net357),
    .B(net389),
    .Y(_0127_));
 sg13g2_a22oi_1 _3542_ (.Y(_1017_),
    .B1(_0977_),
    .B2(net490),
    .A2(_0976_),
    .A1(_1375_));
 sg13g2_nand2b_1 _3543_ (.Y(_0128_),
    .B(net364),
    .A_N(_1017_));
 sg13g2_nor3_1 _3544_ (.A(_0766_),
    .B(_0770_),
    .C(_0774_),
    .Y(_0129_));
 sg13g2_nand2b_1 _3545_ (.Y(_1018_),
    .B(_0718_),
    .A_N(_0710_));
 sg13g2_a21oi_1 _3546_ (.A1(_0712_),
    .A2(_1018_),
    .Y(_0130_),
    .B1(_0717_));
 sg13g2_nor2_1 _3547_ (.A(_0713_),
    .B(_0717_),
    .Y(_0131_));
 sg13g2_nor2b_1 _3548_ (.A(_0716_),
    .B_N(_1018_),
    .Y(_0132_));
 sg13g2_nand3b_1 _3549_ (.B(net6),
    .C(\matt_venn_vga.x_px[8] ),
    .Y(_1019_),
    .A_N(net309));
 sg13g2_nand4_1 _3550_ (.B(net318),
    .C(net319),
    .A(net316),
    .Y(_1020_),
    .D(\h[2] ));
 sg13g2_or2_1 _3551_ (.X(_1021_),
    .B(net321),
    .A(net322));
 sg13g2_nor4_1 _3552_ (.A(_0528_),
    .B(_1019_),
    .C(_1020_),
    .D(_1021_),
    .Y(_1022_));
 sg13g2_nor2_1 _3553_ (.A(net406),
    .B(_1022_),
    .Y(_1023_));
 sg13g2_xnor2_1 _3554_ (.Y(_1024_),
    .A(net318),
    .B(_0506_));
 sg13g2_nor3_1 _3555_ (.A(net319),
    .B(net320),
    .C(_1021_),
    .Y(_1025_));
 sg13g2_and4_1 _3556_ (.A(_1390_),
    .B(_1395_),
    .C(net309),
    .D(_1025_),
    .X(_1026_));
 sg13g2_nand3_1 _3557_ (.B(_1024_),
    .C(_1026_),
    .A(_0532_),
    .Y(_1027_));
 sg13g2_nand4_1 _3558_ (.B(net312),
    .C(net318),
    .A(net314),
    .Y(_1028_),
    .D(_1026_));
 sg13g2_or4_1 _3559_ (.A(net322),
    .B(_1394_),
    .C(_0507_),
    .D(_0531_),
    .X(_1029_));
 sg13g2_o21ai_1 _3560_ (.B1(_1028_),
    .Y(_1030_),
    .A1(_1019_),
    .A2(_1029_));
 sg13g2_a221oi_1 _3561_ (.B2(net316),
    .C1(net359),
    .B1(_1030_),
    .A1(_1023_),
    .Y(_0133_),
    .A2(_1027_));
 sg13g2_o21ai_1 _3562_ (.B1(net297),
    .Y(_1031_),
    .A1(_1374_),
    .A2(_0779_));
 sg13g2_a21oi_1 _3563_ (.A1(_1374_),
    .A2(_1421_),
    .Y(_0134_),
    .B1(_1031_));
 sg13g2_o21ai_1 _3564_ (.B1(_1373_),
    .Y(_1032_),
    .A1(_1374_),
    .A2(_1421_));
 sg13g2_or2_1 _3565_ (.X(_1033_),
    .B(_0779_),
    .A(_1457_));
 sg13g2_and3_1 _3566_ (.X(_0135_),
    .A(net364),
    .B(_1032_),
    .C(_1033_));
 sg13g2_xor2_1 _3567_ (.B(_1033_),
    .A(net336),
    .X(_1034_));
 sg13g2_nor2_1 _3568_ (.A(_0825_),
    .B(_1034_),
    .Y(_0136_));
 sg13g2_nor2_1 _3569_ (.A(_0030_),
    .B(_1033_),
    .Y(_1035_));
 sg13g2_xnor2_1 _3570_ (.Y(_1036_),
    .A(net334),
    .B(_1035_));
 sg13g2_nor2_1 _3571_ (.A(_0825_),
    .B(_1036_),
    .Y(_0137_));
 sg13g2_nor3_2 _3572_ (.A(_1372_),
    .B(_1462_),
    .C(_0779_),
    .Y(_1037_));
 sg13g2_or3_1 _3573_ (.A(_1372_),
    .B(_1421_),
    .C(_1462_),
    .X(_1038_));
 sg13g2_o21ai_1 _3574_ (.B1(net362),
    .Y(_1039_),
    .A1(net332),
    .A2(_1037_));
 sg13g2_a21oi_1 _3575_ (.A1(net332),
    .A2(_1037_),
    .Y(_0138_),
    .B1(_1039_));
 sg13g2_nor2_1 _3576_ (.A(_0026_),
    .B(_1038_),
    .Y(_1040_));
 sg13g2_o21ai_1 _3577_ (.B1(net294),
    .Y(_1041_),
    .A1(net330),
    .A2(_1040_));
 sg13g2_a21oi_1 _3578_ (.A1(net330),
    .A2(_1040_),
    .Y(_0139_),
    .B1(_1041_));
 sg13g2_nand3_1 _3579_ (.B(net332),
    .C(_1037_),
    .A(net330),
    .Y(_1042_));
 sg13g2_nor2_1 _3580_ (.A(_1474_),
    .B(_1038_),
    .Y(_1043_));
 sg13g2_xnor2_1 _3581_ (.Y(_1044_),
    .A(net329),
    .B(_1043_));
 sg13g2_nor2_1 _3582_ (.A(net360),
    .B(_1044_),
    .Y(_0140_));
 sg13g2_nor2_1 _3583_ (.A(net552),
    .B(_1042_),
    .Y(_1045_));
 sg13g2_o21ai_1 _3584_ (.B1(net294),
    .Y(_1046_),
    .A1(net327),
    .A2(_1045_));
 sg13g2_a21oi_1 _3585_ (.A1(net327),
    .A2(_1045_),
    .Y(_0141_),
    .B1(_1046_));
 sg13g2_nand3_1 _3586_ (.B(net329),
    .C(_1043_),
    .A(net328),
    .Y(_1047_));
 sg13g2_xor2_1 _3587_ (.B(_1047_),
    .A(net326),
    .X(_1048_));
 sg13g2_nor2_1 _3588_ (.A(_0825_),
    .B(_1048_),
    .Y(_0142_));
 sg13g2_nor2_1 _3589_ (.A(_0023_),
    .B(_1047_),
    .Y(_1049_));
 sg13g2_o21ai_1 _3590_ (.B1(net294),
    .Y(_1050_),
    .A1(net323),
    .A2(_1049_));
 sg13g2_a21oi_1 _3591_ (.A1(net323),
    .A2(_1049_),
    .Y(_0143_),
    .B1(_1050_));
 sg13g2_nand3_1 _3592_ (.B(net325),
    .C(_1455_),
    .A(net324),
    .Y(_1051_));
 sg13g2_nor2_1 _3593_ (.A(_1372_),
    .B(net337),
    .Y(_1052_));
 sg13g2_nand2_1 _3594_ (.Y(_1053_),
    .A(_1443_),
    .B(_1052_));
 sg13g2_o21ai_1 _3595_ (.B1(net364),
    .Y(_1054_),
    .A1(_1051_),
    .A2(_1053_));
 sg13g2_nor4_1 _3596_ (.A(net339),
    .B(_1374_),
    .C(_1471_),
    .D(_1051_),
    .Y(_1055_));
 sg13g2_nor3_1 _3597_ (.A(_1395_),
    .B(_1054_),
    .C(_1055_),
    .Y(_1056_));
 sg13g2_nand3_1 _3598_ (.B(_1459_),
    .C(_1052_),
    .A(_1447_),
    .Y(_1057_));
 sg13g2_nor4_1 _3599_ (.A(net339),
    .B(net341),
    .C(_1423_),
    .D(_1458_),
    .Y(_1058_));
 sg13g2_nand2_1 _3600_ (.Y(_1059_),
    .A(_1447_),
    .B(_1058_));
 sg13g2_nand4_1 _3601_ (.B(net362),
    .C(_1057_),
    .A(_1395_),
    .Y(_1060_),
    .D(_1059_));
 sg13g2_nand2b_1 _3602_ (.Y(_1061_),
    .B(_1060_),
    .A_N(_1056_));
 sg13g2_nor2b_1 _3603_ (.A(_1054_),
    .B_N(_1059_),
    .Y(_1062_));
 sg13g2_mux2_1 _3604_ (.A0(_1062_),
    .A1(net383),
    .S(_1061_),
    .X(_0144_));
 sg13g2_nand2_1 _3605_ (.Y(_0145_),
    .A(_0520_),
    .B(_1024_));
 sg13g2_xor2_1 _3606_ (.B(_0507_),
    .A(net317),
    .X(_1063_));
 sg13g2_nand2_1 _3607_ (.Y(_0146_),
    .A(_0520_),
    .B(_1063_));
 sg13g2_and2_1 _3608_ (.A(_0773_),
    .B(_0776_),
    .X(_0147_));
 sg13g2_nor3_1 _3609_ (.A(_0710_),
    .B(_0716_),
    .C(_0718_),
    .Y(_0148_));
 sg13g2_nand2_2 _3610_ (.Y(_1064_),
    .A(net367),
    .B(_1421_));
 sg13g2_and3_1 _3611_ (.X(_0149_),
    .A(net367),
    .B(net225),
    .C(_1421_));
 sg13g2_and3_1 _3612_ (.X(_0150_),
    .A(net367),
    .B(_1412_),
    .C(_1021_));
 sg13g2_and2_1 _3613_ (.A(net320),
    .B(_1411_),
    .X(_1065_));
 sg13g2_nor2_1 _3614_ (.A(net320),
    .B(net533),
    .Y(_1066_));
 sg13g2_nor3_1 _3615_ (.A(_1064_),
    .B(_1065_),
    .C(net534),
    .Y(_0151_));
 sg13g2_and2_1 _3616_ (.A(net319),
    .B(_1065_),
    .X(_1067_));
 sg13g2_nor2_1 _3617_ (.A(net319),
    .B(_1065_),
    .Y(_1068_));
 sg13g2_nor3_1 _3618_ (.A(_1064_),
    .B(_1067_),
    .C(_1068_),
    .Y(_0152_));
 sg13g2_nor2b_1 _3619_ (.A(_1410_),
    .B_N(_1065_),
    .Y(_1069_));
 sg13g2_nor2_1 _3620_ (.A(net318),
    .B(_1067_),
    .Y(_1070_));
 sg13g2_nor3_1 _3621_ (.A(_1064_),
    .B(_1069_),
    .C(_1070_),
    .Y(_0153_));
 sg13g2_nor2_2 _3622_ (.A(_1412_),
    .B(_1020_),
    .Y(_1071_));
 sg13g2_nor2_1 _3623_ (.A(net316),
    .B(_1069_),
    .Y(_1072_));
 sg13g2_nor3_1 _3624_ (.A(_1064_),
    .B(_1071_),
    .C(_1072_),
    .Y(_0154_));
 sg13g2_xnor2_1 _3625_ (.Y(_1073_),
    .A(net314),
    .B(net546));
 sg13g2_nor2_1 _3626_ (.A(_1064_),
    .B(_1073_),
    .Y(_0155_));
 sg13g2_nor3_1 _3627_ (.A(net518),
    .B(_1412_),
    .C(_1020_),
    .Y(_1074_));
 sg13g2_xnor2_1 _3628_ (.Y(_1075_),
    .A(net312),
    .B(net519));
 sg13g2_nor2_1 _3629_ (.A(_1064_),
    .B(net520),
    .Y(_0156_));
 sg13g2_nand2b_1 _3630_ (.Y(_1076_),
    .B(_1071_),
    .A_N(_1417_));
 sg13g2_xnor2_1 _3631_ (.Y(_1077_),
    .A(_1390_),
    .B(_1076_));
 sg13g2_nor2_1 _3632_ (.A(_1064_),
    .B(net551),
    .Y(_0157_));
 sg13g2_nor2_1 _3633_ (.A(_0055_),
    .B(_1076_),
    .Y(_1078_));
 sg13g2_xnor2_1 _3634_ (.Y(_1079_),
    .A(net310),
    .B(_1078_));
 sg13g2_nor2_1 _3635_ (.A(_1064_),
    .B(_1079_),
    .Y(_0158_));
 sg13g2_or2_1 _3636_ (.X(_1080_),
    .B(\matt_venn_clock.pulse_hrs.comp[2] ),
    .A(\matt_venn_clock.pulse_hrs.comp[3] ));
 sg13g2_nand2_1 _3637_ (.Y(_1081_),
    .A(_1364_),
    .B(_0068_));
 sg13g2_nor4_2 _3638_ (.A(\matt_venn_clock.pulse_hrs.count[3] ),
    .B(\matt_venn_clock.pulse_hrs.count[1] ),
    .C(\matt_venn_clock.pulse_hrs.count[0] ),
    .Y(_1082_),
    .D(_1081_));
 sg13g2_o21ai_1 _3639_ (.B1(_1082_),
    .Y(_1083_),
    .A1(\matt_venn_clock.pulse_hrs.comp[4] ),
    .A2(_1080_));
 sg13g2_or2_1 _3640_ (.X(_1084_),
    .B(_1083_),
    .A(net300));
 sg13g2_a21oi_1 _3641_ (.A1(net1),
    .A2(_1083_),
    .Y(_1085_),
    .B1(_0778_));
 sg13g2_o21ai_1 _3642_ (.B1(net492),
    .Y(_1086_),
    .A1(_1401_),
    .A2(_1084_));
 sg13g2_nand2b_1 _3643_ (.Y(_1087_),
    .B(_1085_),
    .A_N(net492));
 sg13g2_a21oi_1 _3644_ (.A1(net1),
    .A2(_1083_),
    .Y(_1088_),
    .B1(net300));
 sg13g2_nand3_1 _3645_ (.B(_1086_),
    .C(_1087_),
    .A(net369),
    .Y(_0159_));
 sg13g2_a21oi_2 _3646_ (.B1(net358),
    .Y(_1089_),
    .A2(net301),
    .A1(_1401_));
 sg13g2_nor2_1 _3647_ (.A(\matt_venn_clock.pulse_hrs.comp[1] ),
    .B(\matt_venn_clock.pulse_hrs.comp[0] ),
    .Y(_1090_));
 sg13g2_o21ai_1 _3648_ (.B1(_1089_),
    .Y(_1091_),
    .A1(net474),
    .A2(_1087_));
 sg13g2_a21o_1 _3649_ (.A2(_1087_),
    .A1(net474),
    .B1(_1091_),
    .X(_0160_));
 sg13g2_o21ai_1 _3650_ (.B1(net450),
    .Y(_1092_),
    .A1(\matt_venn_clock.pulse_hrs.comp[1] ),
    .A2(_1087_));
 sg13g2_nand3_1 _3651_ (.B(_1088_),
    .C(_1090_),
    .A(_1366_),
    .Y(_1093_));
 sg13g2_nand3_1 _3652_ (.B(net451),
    .C(_1093_),
    .A(_1089_),
    .Y(_0161_));
 sg13g2_or4_1 _3653_ (.A(\matt_venn_clock.pulse_hrs.comp[1] ),
    .B(\matt_venn_clock.pulse_hrs.comp[0] ),
    .C(_1080_),
    .D(_1084_),
    .X(_1094_));
 sg13g2_nand2_1 _3654_ (.Y(_1095_),
    .A(net432),
    .B(_1093_));
 sg13g2_nand3_1 _3655_ (.B(_1094_),
    .C(_1095_),
    .A(_1089_),
    .Y(_0162_));
 sg13g2_and3_1 _3656_ (.X(_0163_),
    .A(net254),
    .B(_1089_),
    .C(_1094_));
 sg13g2_xor2_1 _3657_ (.B(\matt_venn_clock.pulse_hrs.comp[4] ),
    .A(\matt_venn_clock.pulse_hrs.count[4] ),
    .X(_1096_));
 sg13g2_xnor2_1 _3658_ (.Y(_1097_),
    .A(\matt_venn_clock.pulse_hrs.count[3] ),
    .B(\matt_venn_clock.pulse_hrs.comp[3] ));
 sg13g2_a221oi_1 _3659_ (.B2(\matt_venn_clock.pulse_hrs.count[1] ),
    .C1(_1096_),
    .B1(_1367_),
    .A1(_1364_),
    .Y(_1098_),
    .A2(\matt_venn_clock.pulse_hrs.comp[2] ));
 sg13g2_xnor2_1 _3660_ (.Y(_1099_),
    .A(\matt_venn_clock.pulse_hrs.count[0] ),
    .B(\matt_venn_clock.pulse_hrs.comp[0] ));
 sg13g2_a22oi_1 _3661_ (.Y(_1100_),
    .B1(\matt_venn_clock.pulse_hrs.comp[1] ),
    .B2(_1365_),
    .A2(_1366_),
    .A1(\matt_venn_clock.pulse_hrs.count[2] ));
 sg13g2_nand4_1 _3662_ (.B(_1098_),
    .C(_1099_),
    .A(_1097_),
    .Y(_1101_),
    .D(_1100_));
 sg13g2_and3_1 _3663_ (.X(_1102_),
    .A(net1),
    .B(_0780_),
    .C(_1101_));
 sg13g2_nand2_1 _3664_ (.Y(_1103_),
    .A(net542),
    .B(net301));
 sg13g2_o21ai_1 _3665_ (.B1(_1103_),
    .Y(_1104_),
    .A1(net542),
    .A2(_1102_));
 sg13g2_nor2_1 _3666_ (.A(net357),
    .B(_1104_),
    .Y(_0164_));
 sg13g2_nand2_1 _3667_ (.Y(_1105_),
    .A(net496),
    .B(net295));
 sg13g2_nand2_2 _3668_ (.Y(_1106_),
    .A(net369),
    .B(_1102_));
 sg13g2_inv_1 _3669_ (.Y(_1107_),
    .A(_1106_));
 sg13g2_xnor2_1 _3670_ (.Y(_1108_),
    .A(net496),
    .B(\matt_venn_clock.pulse_hrs.count[0] ));
 sg13g2_o21ai_1 _3671_ (.B1(_1105_),
    .Y(_0165_),
    .A1(_1106_),
    .A2(_1108_));
 sg13g2_a21oi_1 _3672_ (.A1(\matt_venn_clock.pulse_hrs.count[1] ),
    .A2(\matt_venn_clock.pulse_hrs.count[0] ),
    .Y(_1109_),
    .B1(net399));
 sg13g2_nand3_1 _3673_ (.B(\matt_venn_clock.pulse_hrs.count[1] ),
    .C(\matt_venn_clock.pulse_hrs.count[0] ),
    .A(\matt_venn_clock.pulse_hrs.count[2] ),
    .Y(_1110_));
 sg13g2_a22oi_1 _3674_ (.Y(_1111_),
    .B1(_1107_),
    .B2(_1110_),
    .A2(net295),
    .A1(net399));
 sg13g2_nor2_1 _3675_ (.A(net400),
    .B(_1111_),
    .Y(_0166_));
 sg13g2_nand2_1 _3676_ (.Y(_1112_),
    .A(net444),
    .B(net295));
 sg13g2_nand4_1 _3677_ (.B(\matt_venn_clock.pulse_hrs.count[2] ),
    .C(\matt_venn_clock.pulse_hrs.count[1] ),
    .A(\matt_venn_clock.pulse_hrs.count[3] ),
    .Y(_1113_),
    .D(\matt_venn_clock.pulse_hrs.count[0] ));
 sg13g2_xor2_1 _3678_ (.B(_1110_),
    .A(net444),
    .X(_1114_));
 sg13g2_o21ai_1 _3679_ (.B1(_1112_),
    .Y(_0167_),
    .A1(_1106_),
    .A2(_1114_));
 sg13g2_nand2_1 _3680_ (.Y(_1115_),
    .A(net265),
    .B(net297));
 sg13g2_xnor2_1 _3681_ (.Y(_1116_),
    .A(_0068_),
    .B(_1113_));
 sg13g2_o21ai_1 _3682_ (.B1(_1115_),
    .Y(_0168_),
    .A1(_1106_),
    .A2(_1116_));
 sg13g2_or2_1 _3683_ (.X(_1117_),
    .B(\matt_venn_clock.pulse_min.comp[2] ),
    .A(\matt_venn_clock.pulse_min.comp[3] ));
 sg13g2_nand2b_1 _3684_ (.Y(_1118_),
    .B(_0067_),
    .A_N(\matt_venn_clock.pulse_min.count[2] ));
 sg13g2_nor4_2 _3685_ (.A(\matt_venn_clock.pulse_min.count[3] ),
    .B(\matt_venn_clock.pulse_min.count[1] ),
    .C(\matt_venn_clock.pulse_min.count[0] ),
    .Y(_1119_),
    .D(_1118_));
 sg13g2_o21ai_1 _3686_ (.B1(_1119_),
    .Y(_1120_),
    .A1(\matt_venn_clock.pulse_min.comp[4] ),
    .A2(_1117_));
 sg13g2_or2_1 _3687_ (.X(_1121_),
    .B(_1120_),
    .A(net300));
 sg13g2_a21oi_1 _3688_ (.A1(net2),
    .A2(_1120_),
    .Y(_1122_),
    .B1(_0778_));
 sg13g2_o21ai_1 _3689_ (.B1(net458),
    .Y(_1123_),
    .A1(_1400_),
    .A2(_1121_));
 sg13g2_nand2b_1 _3690_ (.Y(_1124_),
    .B(_1122_),
    .A_N(net458));
 sg13g2_nand3_1 _3691_ (.B(_1123_),
    .C(_1124_),
    .A(net369),
    .Y(_0169_));
 sg13g2_nand2_1 _3692_ (.Y(_1125_),
    .A(net418),
    .B(_1124_));
 sg13g2_a21oi_2 _3693_ (.B1(net358),
    .Y(_1126_),
    .A2(net301),
    .A1(_1400_));
 sg13g2_nand2b_1 _3694_ (.Y(_1127_),
    .B(_1363_),
    .A_N(_1124_));
 sg13g2_nand3_1 _3695_ (.B(_1126_),
    .C(_1127_),
    .A(net419),
    .Y(_0170_));
 sg13g2_o21ai_1 _3696_ (.B1(_1126_),
    .Y(_1128_),
    .A1(net434),
    .A2(_1127_));
 sg13g2_a21o_1 _3697_ (.A2(_1127_),
    .A1(net434),
    .B1(_1128_),
    .X(_0171_));
 sg13g2_or4_1 _3698_ (.A(net418),
    .B(net458),
    .C(_1117_),
    .D(_1121_),
    .X(_1129_));
 sg13g2_o21ai_1 _3699_ (.B1(net459),
    .Y(_1130_),
    .A1(net434),
    .A2(_1127_));
 sg13g2_nand3_1 _3700_ (.B(_1129_),
    .C(_1130_),
    .A(_1126_),
    .Y(_0172_));
 sg13g2_and3_1 _3701_ (.X(_0173_),
    .A(net255),
    .B(_1126_),
    .C(_1129_));
 sg13g2_a22oi_1 _3702_ (.Y(_1131_),
    .B1(\matt_venn_clock.pulse_min.comp[1] ),
    .B2(_1360_),
    .A2(_1361_),
    .A1(\matt_venn_clock.pulse_min.count[4] ));
 sg13g2_xnor2_1 _3703_ (.Y(_1132_),
    .A(\matt_venn_clock.pulse_min.count[2] ),
    .B(\matt_venn_clock.pulse_min.comp[2] ));
 sg13g2_xor2_1 _3704_ (.B(\matt_venn_clock.pulse_min.comp[0] ),
    .A(\matt_venn_clock.pulse_min.count[0] ),
    .X(_1133_));
 sg13g2_a221oi_1 _3705_ (.B2(\matt_venn_clock.pulse_min.count[1] ),
    .C1(_1133_),
    .B1(_1363_),
    .A1(_1359_),
    .Y(_1134_),
    .A2(\matt_venn_clock.pulse_min.comp[3] ));
 sg13g2_a22oi_1 _3706_ (.Y(_1135_),
    .B1(_1362_),
    .B2(\matt_venn_clock.pulse_min.count[3] ),
    .A2(\matt_venn_clock.pulse_min.comp[4] ),
    .A1(_1358_));
 sg13g2_nand4_1 _3707_ (.B(_1132_),
    .C(_1134_),
    .A(_1131_),
    .Y(_1136_),
    .D(_1135_));
 sg13g2_and3_1 _3708_ (.X(_1137_),
    .A(net2),
    .B(net301),
    .C(_1136_));
 sg13g2_nand2_1 _3709_ (.Y(_1138_),
    .A(net539),
    .B(net301));
 sg13g2_o21ai_1 _3710_ (.B1(_1138_),
    .Y(_1139_),
    .A1(net539),
    .A2(_1137_));
 sg13g2_nor2_1 _3711_ (.A(net358),
    .B(_1139_),
    .Y(_0174_));
 sg13g2_nand2_1 _3712_ (.Y(_1140_),
    .A(net454),
    .B(net296));
 sg13g2_nand2_2 _3713_ (.Y(_1141_),
    .A(net369),
    .B(_1137_));
 sg13g2_xnor2_1 _3714_ (.Y(_1142_),
    .A(net454),
    .B(\matt_venn_clock.pulse_min.count[0] ));
 sg13g2_o21ai_1 _3715_ (.B1(_1140_),
    .Y(_0175_),
    .A1(_1141_),
    .A2(_1142_));
 sg13g2_nand2_1 _3716_ (.Y(_1143_),
    .A(net395),
    .B(net296));
 sg13g2_nand3_1 _3717_ (.B(\matt_venn_clock.pulse_min.count[1] ),
    .C(\matt_venn_clock.pulse_min.count[0] ),
    .A(\matt_venn_clock.pulse_min.count[2] ),
    .Y(_1144_));
 sg13g2_a21o_1 _3718_ (.A2(\matt_venn_clock.pulse_min.count[0] ),
    .A1(net559),
    .B1(net395),
    .X(_1145_));
 sg13g2_nand2_1 _3719_ (.Y(_1146_),
    .A(_1144_),
    .B(net560));
 sg13g2_o21ai_1 _3720_ (.B1(_1143_),
    .Y(_0176_),
    .A1(_1141_),
    .A2(_1146_));
 sg13g2_nand2_1 _3721_ (.Y(_1147_),
    .A(net276),
    .B(net296));
 sg13g2_or2_1 _3722_ (.X(_1148_),
    .B(_1144_),
    .A(_1359_));
 sg13g2_xnor2_1 _3723_ (.Y(_1149_),
    .A(_1359_),
    .B(_1144_));
 sg13g2_o21ai_1 _3724_ (.B1(_1147_),
    .Y(_0177_),
    .A1(_1141_),
    .A2(_1149_));
 sg13g2_nand2_1 _3725_ (.Y(_1150_),
    .A(net256),
    .B(net295));
 sg13g2_xnor2_1 _3726_ (.Y(_1151_),
    .A(_0067_),
    .B(_1148_));
 sg13g2_o21ai_1 _3727_ (.B1(_1150_),
    .Y(_0178_),
    .A1(_1141_),
    .A2(_1151_));
 sg13g2_nor3_1 _3728_ (.A(\matt_venn_clock.pulse_sec.comp[4] ),
    .B(\matt_venn_clock.pulse_sec.comp[3] ),
    .C(\matt_venn_clock.pulse_sec.comp[2] ),
    .Y(_1152_));
 sg13g2_nor2_1 _3729_ (.A(net482),
    .B(\matt_venn_clock.pulse_sec.count[0] ),
    .Y(_1153_));
 sg13g2_nand4_1 _3730_ (.B(_1355_),
    .C(_0066_),
    .A(_1354_),
    .Y(_1154_),
    .D(_1153_));
 sg13g2_or2_1 _3731_ (.X(_1155_),
    .B(_1154_),
    .A(_1152_));
 sg13g2_or2_1 _3732_ (.X(_1156_),
    .B(_1155_),
    .A(net300));
 sg13g2_a21oi_1 _3733_ (.A1(net3),
    .A2(_1155_),
    .Y(_1157_),
    .B1(_0778_));
 sg13g2_o21ai_1 _3734_ (.B1(net443),
    .Y(_1158_),
    .A1(_1399_),
    .A2(_1156_));
 sg13g2_nand2_1 _3735_ (.Y(_1159_),
    .A(_1357_),
    .B(_1157_));
 sg13g2_nand3_1 _3736_ (.B(_1158_),
    .C(_1159_),
    .A(net369),
    .Y(_0179_));
 sg13g2_nand2_1 _3737_ (.Y(_1160_),
    .A(net373),
    .B(_1159_));
 sg13g2_a21oi_2 _3738_ (.B1(net357),
    .Y(_1161_),
    .A2(net302),
    .A1(_1399_));
 sg13g2_nand3_1 _3739_ (.B(_1357_),
    .C(_1157_),
    .A(_1356_),
    .Y(_1162_));
 sg13g2_nand3_1 _3740_ (.B(_1161_),
    .C(_1162_),
    .A(net374),
    .Y(_0180_));
 sg13g2_o21ai_1 _3741_ (.B1(_1161_),
    .Y(_1163_),
    .A1(net478),
    .A2(_1162_));
 sg13g2_a21o_1 _3742_ (.A2(_1162_),
    .A1(net478),
    .B1(_1163_),
    .X(_0181_));
 sg13g2_nor4_1 _3743_ (.A(net493),
    .B(net478),
    .C(net373),
    .D(net443),
    .Y(_1164_));
 sg13g2_nand2b_1 _3744_ (.Y(_1165_),
    .B(_1164_),
    .A_N(_1156_));
 sg13g2_o21ai_1 _3745_ (.B1(net493),
    .Y(_1166_),
    .A1(net478),
    .A2(_1162_));
 sg13g2_nand3_1 _3746_ (.B(_1165_),
    .C(_1166_),
    .A(_1161_),
    .Y(_0182_));
 sg13g2_and3_1 _3747_ (.X(_0183_),
    .A(net273),
    .B(_1161_),
    .C(_1165_));
 sg13g2_a22oi_1 _3748_ (.Y(_1167_),
    .B1(_1357_),
    .B2(\matt_venn_clock.pulse_sec.count[0] ),
    .A2(\matt_venn_clock.pulse_sec.comp[4] ),
    .A1(_1353_));
 sg13g2_nor2_1 _3749_ (.A(\matt_venn_clock.pulse_sec.count[0] ),
    .B(_1357_),
    .Y(_1168_));
 sg13g2_nor2_1 _3750_ (.A(_1354_),
    .B(\matt_venn_clock.pulse_sec.comp[3] ),
    .Y(_1169_));
 sg13g2_nor2_1 _3751_ (.A(\matt_venn_clock.pulse_sec.count[1] ),
    .B(_1356_),
    .Y(_1170_));
 sg13g2_nor2_1 _3752_ (.A(_1353_),
    .B(\matt_venn_clock.pulse_sec.comp[4] ),
    .Y(_1171_));
 sg13g2_a22oi_1 _3753_ (.Y(_1172_),
    .B1(_1356_),
    .B2(\matt_venn_clock.pulse_sec.count[1] ),
    .A2(\matt_venn_clock.pulse_sec.comp[3] ),
    .A1(_1354_));
 sg13g2_xnor2_1 _3754_ (.Y(_1173_),
    .A(\matt_venn_clock.pulse_sec.count[2] ),
    .B(\matt_venn_clock.pulse_sec.comp[2] ));
 sg13g2_nor4_1 _3755_ (.A(_1168_),
    .B(_1169_),
    .C(_1170_),
    .D(_1171_),
    .Y(_1174_));
 sg13g2_nand4_1 _3756_ (.B(_1172_),
    .C(_1173_),
    .A(_1167_),
    .Y(_1175_),
    .D(_1174_));
 sg13g2_and3_1 _3757_ (.X(_1176_),
    .A(net3),
    .B(net301),
    .C(_1175_));
 sg13g2_nand2_1 _3758_ (.Y(_1177_),
    .A(net516),
    .B(net301));
 sg13g2_o21ai_1 _3759_ (.B1(_1177_),
    .Y(_1178_),
    .A1(net516),
    .A2(_1176_));
 sg13g2_nor2_1 _3760_ (.A(net357),
    .B(_1178_),
    .Y(_0184_));
 sg13g2_nand2_1 _3761_ (.Y(_1179_),
    .A(net369),
    .B(_1176_));
 sg13g2_inv_1 _3762_ (.Y(_1180_),
    .A(_1179_));
 sg13g2_nand2_1 _3763_ (.Y(_1181_),
    .A(net482),
    .B(\matt_venn_clock.pulse_sec.count[0] ));
 sg13g2_a22oi_1 _3764_ (.Y(_1182_),
    .B1(_1180_),
    .B2(_1181_),
    .A2(net295),
    .A1(net482));
 sg13g2_nor2_1 _3765_ (.A(_1153_),
    .B(net483),
    .Y(_0185_));
 sg13g2_nand3_1 _3766_ (.B(\matt_venn_clock.pulse_sec.count[1] ),
    .C(\matt_venn_clock.pulse_sec.count[0] ),
    .A(net427),
    .Y(_1183_));
 sg13g2_a22oi_1 _3767_ (.Y(_1184_),
    .B1(_1180_),
    .B2(_1183_),
    .A2(net295),
    .A1(net427));
 sg13g2_a21oi_1 _3768_ (.A1(_1355_),
    .A2(_1181_),
    .Y(_0186_),
    .B1(_1184_));
 sg13g2_nand2_1 _3769_ (.Y(_1185_),
    .A(net248),
    .B(net295));
 sg13g2_or2_1 _3770_ (.X(_1186_),
    .B(_1183_),
    .A(_1354_));
 sg13g2_xnor2_1 _3771_ (.Y(_1187_),
    .A(_1354_),
    .B(_1183_));
 sg13g2_o21ai_1 _3772_ (.B1(_1185_),
    .Y(_0187_),
    .A1(_1179_),
    .A2(_1187_));
 sg13g2_nand2_1 _3773_ (.Y(_1188_),
    .A(net243),
    .B(net295));
 sg13g2_xnor2_1 _3774_ (.Y(_1189_),
    .A(_0066_),
    .B(_1186_));
 sg13g2_o21ai_1 _3775_ (.B1(_1188_),
    .Y(_0188_),
    .A1(_1179_),
    .A2(_1189_));
 sg13g2_nand3b_1 _3776_ (.B(\clock_sec_d[1] ),
    .C(\clock_sec_d[2] ),
    .Y(_1190_),
    .A_N(\clock_sec_d[0] ));
 sg13g2_and3_2 _3777_ (.X(_1191_),
    .A(net2),
    .B(net302),
    .C(_1119_));
 sg13g2_inv_1 _3778_ (.Y(_1192_),
    .A(_1191_));
 sg13g2_nand2_2 _3779_ (.Y(_1193_),
    .A(_1190_),
    .B(_1192_));
 sg13g2_o21ai_1 _3780_ (.B1(net365),
    .Y(_1194_),
    .A1(\clock_color_offset[0] ),
    .A2(_1193_));
 sg13g2_a21oi_1 _3781_ (.A1(_1352_),
    .A2(_1193_),
    .Y(_0189_),
    .B1(_1194_));
 sg13g2_a21oi_1 _3782_ (.A1(\clock_color_offset[0] ),
    .A2(_1193_),
    .Y(_1195_),
    .B1(net402));
 sg13g2_nand3_1 _3783_ (.B(\clock_color_offset[0] ),
    .C(_1193_),
    .A(net402),
    .Y(_1196_));
 sg13g2_nand2_1 _3784_ (.Y(_1197_),
    .A(net365),
    .B(_1196_));
 sg13g2_nor2_1 _3785_ (.A(net403),
    .B(_1197_),
    .Y(_0190_));
 sg13g2_o21ai_1 _3786_ (.B1(net365),
    .Y(_1198_),
    .A1(_1351_),
    .A2(_1196_));
 sg13g2_a21oi_1 _3787_ (.A1(_1351_),
    .A2(_1196_),
    .Y(_0191_),
    .B1(_1198_));
 sg13g2_nor2_1 _3788_ (.A(net431),
    .B(\clock_hrs_u[0] ),
    .Y(_1199_));
 sg13g2_nand3_1 _3789_ (.B(\clock_hrs_d[1] ),
    .C(_1199_),
    .A(\clock_hrs_u[2] ),
    .Y(_1200_));
 sg13g2_nor3_2 _3790_ (.A(\clock_hrs_u[3] ),
    .B(\clock_hrs_d[0] ),
    .C(_1200_),
    .Y(_1201_));
 sg13g2_nand2b_1 _3791_ (.Y(_1202_),
    .B(net366),
    .A_N(_1201_));
 sg13g2_nand2_1 _3792_ (.Y(_1203_),
    .A(\clock_hrs_u[3] ),
    .B(\clock_hrs_u[1] ));
 sg13g2_nor3_2 _3793_ (.A(\clock_hrs_u[2] ),
    .B(\clock_hrs_u[0] ),
    .C(_1203_),
    .Y(_1204_));
 sg13g2_nand2b_1 _3794_ (.Y(_1205_),
    .B(\clock_hrs_d[0] ),
    .A_N(_1204_));
 sg13g2_nand2_1 _3795_ (.Y(_1206_),
    .A(net230),
    .B(_1204_));
 sg13g2_a21oi_1 _3796_ (.A1(_1205_),
    .A2(net231),
    .Y(_0192_),
    .B1(_1202_));
 sg13g2_nand2_1 _3797_ (.Y(_1207_),
    .A(\clock_hrs_d[0] ),
    .B(_1204_));
 sg13g2_xor2_1 _3798_ (.B(_1207_),
    .A(net390),
    .X(_1208_));
 sg13g2_nor2_1 _3799_ (.A(_1202_),
    .B(net391),
    .Y(_0193_));
 sg13g2_nand3b_1 _3800_ (.B(\clock_min_d[1] ),
    .C(\clock_min_d[2] ),
    .Y(_1209_),
    .A_N(\clock_min_d[0] ));
 sg13g2_nor2_1 _3801_ (.A(_1201_),
    .B(_1204_),
    .Y(_1210_));
 sg13g2_and3_2 _3802_ (.X(_1211_),
    .A(net1),
    .B(_0780_),
    .C(_1082_));
 sg13g2_inv_1 _3803_ (.Y(_1212_),
    .A(_1211_));
 sg13g2_nand3_1 _3804_ (.B(_1210_),
    .C(_1212_),
    .A(_1209_),
    .Y(_1213_));
 sg13g2_nor4_1 _3805_ (.A(\clock_hrs_u[0] ),
    .B(_1201_),
    .C(_1204_),
    .D(_1211_),
    .Y(_1214_));
 sg13g2_a21oi_1 _3806_ (.A1(net375),
    .A2(_1211_),
    .Y(_1215_),
    .B1(_1214_));
 sg13g2_o21ai_1 _3807_ (.B1(net366),
    .Y(_1216_),
    .A1(_1213_),
    .A2(_1215_));
 sg13g2_a21oi_1 _3808_ (.A1(_1213_),
    .A2(net376),
    .Y(_0194_),
    .B1(_1216_));
 sg13g2_nand2_1 _3809_ (.Y(_1217_),
    .A(net431),
    .B(\clock_hrs_u[0] ));
 sg13g2_a21oi_1 _3810_ (.A1(_1204_),
    .A2(_1212_),
    .Y(_1218_),
    .B1(_1199_));
 sg13g2_nand2_1 _3811_ (.Y(_1219_),
    .A(_1217_),
    .B(_1218_));
 sg13g2_o21ai_1 _3812_ (.B1(net366),
    .Y(_1220_),
    .A1(net431),
    .A2(_1213_));
 sg13g2_a21oi_1 _3813_ (.A1(_1213_),
    .A2(_1219_),
    .Y(_0195_),
    .B1(_1220_));
 sg13g2_nor2_1 _3814_ (.A(_0042_),
    .B(_1217_),
    .Y(_1221_));
 sg13g2_xor2_1 _3815_ (.B(_1217_),
    .A(_0042_),
    .X(_1222_));
 sg13g2_o21ai_1 _3816_ (.B1(_1222_),
    .Y(_1223_),
    .A1(_1210_),
    .A2(_1211_));
 sg13g2_o21ai_1 _3817_ (.B1(net366),
    .Y(_1224_),
    .A1(net461),
    .A2(_1213_));
 sg13g2_a21oi_1 _3818_ (.A1(_1213_),
    .A2(_1223_),
    .Y(_0196_),
    .B1(_1224_));
 sg13g2_xnor2_1 _3819_ (.Y(_1225_),
    .A(_0039_),
    .B(_1221_));
 sg13g2_o21ai_1 _3820_ (.B1(_1225_),
    .Y(_1226_),
    .A1(_1210_),
    .A2(_1211_));
 sg13g2_nand2_1 _3821_ (.Y(_1227_),
    .A(_1213_),
    .B(_1226_));
 sg13g2_o21ai_1 _3822_ (.B1(_1227_),
    .Y(_1228_),
    .A1(net448),
    .A2(_1213_));
 sg13g2_nor2_1 _3823_ (.A(net359),
    .B(net449),
    .Y(_0197_));
 sg13g2_nand2_1 _3824_ (.Y(_1229_),
    .A(net238),
    .B(\clock_min_u[1] ));
 sg13g2_nor3_2 _3825_ (.A(net487),
    .B(\clock_min_u[0] ),
    .C(_1229_),
    .Y(_1230_));
 sg13g2_inv_1 _3826_ (.Y(_1231_),
    .A(_1230_));
 sg13g2_nor2_1 _3827_ (.A(net235),
    .B(_1231_),
    .Y(_1232_));
 sg13g2_nand2_1 _3828_ (.Y(_1233_),
    .A(net366),
    .B(_1209_));
 sg13g2_nor2_1 _3829_ (.A(\clock_min_d[0] ),
    .B(_1230_),
    .Y(_1234_));
 sg13g2_nor3_1 _3830_ (.A(_1232_),
    .B(_1233_),
    .C(_1234_),
    .Y(_0198_));
 sg13g2_nand3_1 _3831_ (.B(\clock_min_d[0] ),
    .C(_1230_),
    .A(net509),
    .Y(_1235_));
 sg13g2_a21oi_1 _3832_ (.A1(\clock_min_d[0] ),
    .A2(_1230_),
    .Y(_1236_),
    .B1(net509));
 sg13g2_nor2_1 _3833_ (.A(_1233_),
    .B(net510),
    .Y(_1237_));
 sg13g2_and2_1 _3834_ (.A(_1235_),
    .B(_1237_),
    .X(_0199_));
 sg13g2_xor2_1 _3835_ (.B(_1235_),
    .A(net409),
    .X(_1238_));
 sg13g2_nor2_1 _3836_ (.A(_1233_),
    .B(net410),
    .Y(_0200_));
 sg13g2_nor2_2 _3837_ (.A(_1193_),
    .B(_1230_),
    .Y(_1239_));
 sg13g2_nor3_1 _3838_ (.A(\clock_min_u[0] ),
    .B(_1191_),
    .C(_1230_),
    .Y(_1240_));
 sg13g2_a21o_1 _3839_ (.A2(_1191_),
    .A1(net397),
    .B1(_1240_),
    .X(_1241_));
 sg13g2_o21ai_1 _3840_ (.B1(net365),
    .Y(_1242_),
    .A1(_1239_),
    .A2(_1241_));
 sg13g2_a21oi_1 _3841_ (.A1(_1239_),
    .A2(_1241_),
    .Y(_0201_),
    .B1(_1242_));
 sg13g2_nand2_1 _3842_ (.Y(_1243_),
    .A(\clock_min_u[0] ),
    .B(_1193_));
 sg13g2_o21ai_1 _3843_ (.B1(net365),
    .Y(_1244_),
    .A1(_1191_),
    .A2(_1231_));
 sg13g2_nand2_1 _3844_ (.Y(_1245_),
    .A(\clock_min_u[1] ),
    .B(\clock_min_u[0] ));
 sg13g2_xor2_1 _3845_ (.B(_1243_),
    .A(net494),
    .X(_1246_));
 sg13g2_nor2_1 _3846_ (.A(_1244_),
    .B(net495),
    .Y(_0202_));
 sg13g2_nor2_1 _3847_ (.A(_0044_),
    .B(_1245_),
    .Y(_1247_));
 sg13g2_xnor2_1 _3848_ (.Y(_1248_),
    .A(_1404_),
    .B(_1245_));
 sg13g2_nor2_1 _3849_ (.A(_1239_),
    .B(_1248_),
    .Y(_1249_));
 sg13g2_nor3_1 _3850_ (.A(net487),
    .B(_1193_),
    .C(_1230_),
    .Y(_1250_));
 sg13g2_nor3_1 _3851_ (.A(_1244_),
    .B(_1249_),
    .C(_1250_),
    .Y(_0203_));
 sg13g2_xnor2_1 _3852_ (.Y(_1251_),
    .A(_0040_),
    .B(_1247_));
 sg13g2_nand2_1 _3853_ (.Y(_1252_),
    .A(_1193_),
    .B(_1251_));
 sg13g2_nand3_1 _3854_ (.B(net365),
    .C(_1239_),
    .A(net238),
    .Y(_1253_));
 sg13g2_o21ai_1 _3855_ (.B1(_1253_),
    .Y(_0204_),
    .A1(_1244_),
    .A2(_1252_));
 sg13g2_nand2_1 _3856_ (.Y(_1254_),
    .A(net250),
    .B(\clock_sec_u[1] ));
 sg13g2_nor3_2 _3857_ (.A(net258),
    .B(\clock_sec_u[0] ),
    .C(_1254_),
    .Y(_1255_));
 sg13g2_nor2b_1 _3858_ (.A(net271),
    .B_N(_1255_),
    .Y(_1256_));
 sg13g2_nand2_1 _3859_ (.Y(_1257_),
    .A(net366),
    .B(_1190_));
 sg13g2_nor2_1 _3860_ (.A(\clock_sec_d[0] ),
    .B(_1255_),
    .Y(_1258_));
 sg13g2_nor3_1 _3861_ (.A(_1256_),
    .B(_1257_),
    .C(_1258_),
    .Y(_0205_));
 sg13g2_nand3_1 _3862_ (.B(net525),
    .C(_1255_),
    .A(\clock_sec_d[1] ),
    .Y(_1259_));
 sg13g2_a21oi_1 _3863_ (.A1(net525),
    .A2(_1255_),
    .Y(_1260_),
    .B1(\clock_sec_d[1] ));
 sg13g2_nor2_1 _3864_ (.A(_1257_),
    .B(net526),
    .Y(_1261_));
 sg13g2_and2_1 _3865_ (.A(_1259_),
    .B(_1261_),
    .X(_0206_));
 sg13g2_xor2_1 _3866_ (.B(_1259_),
    .A(net392),
    .X(_1262_));
 sg13g2_nor2_1 _3867_ (.A(_1257_),
    .B(net393),
    .Y(_0207_));
 sg13g2_or3_1 _3868_ (.A(_1399_),
    .B(_0778_),
    .C(_1154_),
    .X(_1263_));
 sg13g2_and3_1 _3869_ (.X(_1264_),
    .A(\matt_venn_clock.sec_counter[0] ),
    .B(net240),
    .C(\matt_venn_clock.sec_counter[1] ));
 sg13g2_and2_1 _3870_ (.A(net252),
    .B(_1264_),
    .X(_1265_));
 sg13g2_and2_1 _3871_ (.A(net246),
    .B(_1265_),
    .X(_1266_));
 sg13g2_and2_1 _3872_ (.A(net264),
    .B(_1266_),
    .X(_1267_));
 sg13g2_and2_1 _3873_ (.A(net270),
    .B(_1267_),
    .X(_1268_));
 sg13g2_and2_1 _3874_ (.A(net275),
    .B(_1268_),
    .X(_1269_));
 sg13g2_nand3_1 _3875_ (.B(net506),
    .C(_1269_),
    .A(net561),
    .Y(_1270_));
 sg13g2_nor2_1 _3876_ (.A(_1389_),
    .B(_1270_),
    .Y(_1271_));
 sg13g2_and2_1 _3877_ (.A(\matt_venn_clock.sec_counter[11] ),
    .B(_1271_),
    .X(_1272_));
 sg13g2_and4_1 _3878_ (.A(\matt_venn_clock.sec_counter[12] ),
    .B(\matt_venn_clock.sec_counter[13] ),
    .C(\matt_venn_clock.sec_counter[14] ),
    .D(_1272_),
    .X(_1273_));
 sg13g2_nand4_1 _3879_ (.B(\matt_venn_clock.sec_counter[17] ),
    .C(\matt_venn_clock.sec_counter[15] ),
    .A(\matt_venn_clock.sec_counter[16] ),
    .Y(_1274_),
    .D(_1273_));
 sg13g2_nand2_1 _3880_ (.Y(_1275_),
    .A(\matt_venn_clock.sec_counter[18] ),
    .B(net384));
 sg13g2_nor2_2 _3881_ (.A(_1274_),
    .B(_1275_),
    .Y(_1276_));
 sg13g2_and3_1 _3882_ (.X(_1277_),
    .A(\matt_venn_clock.sec_counter[12] ),
    .B(\matt_venn_clock.sec_counter[13] ),
    .C(_1272_));
 sg13g2_and4_1 _3883_ (.A(\matt_venn_clock.sec_counter[14] ),
    .B(\matt_venn_clock.sec_counter[16] ),
    .C(net470),
    .D(_1277_),
    .X(_1278_));
 sg13g2_nand2_1 _3884_ (.Y(_1279_),
    .A(net476),
    .B(_1278_));
 sg13g2_and3_1 _3885_ (.X(_1280_),
    .A(\matt_venn_clock.sec_counter[20] ),
    .B(net260),
    .C(_1276_));
 sg13g2_and2_1 _3886_ (.A(\matt_venn_clock.sec_counter[22] ),
    .B(_1280_),
    .X(_1281_));
 sg13g2_nand2_1 _3887_ (.Y(_1282_),
    .A(\matt_venn_clock.sec_counter[23] ),
    .B(_1281_));
 sg13g2_xor2_1 _3888_ (.B(_1281_),
    .A(net515),
    .X(_1283_));
 sg13g2_a21oi_1 _3889_ (.A1(net470),
    .A2(_1273_),
    .Y(_1284_),
    .B1(net522));
 sg13g2_or2_1 _3890_ (.X(_1285_),
    .B(_1284_),
    .A(_1278_));
 sg13g2_xnor2_1 _3891_ (.Y(_1286_),
    .A(net470),
    .B(_1273_));
 sg13g2_xor2_1 _3892_ (.B(_1277_),
    .A(net504),
    .X(_1287_));
 sg13g2_nor2b_1 _3893_ (.A(net412),
    .B_N(_1272_),
    .Y(_1288_));
 sg13g2_xor2_1 _3894_ (.B(_1272_),
    .A(net412),
    .X(_1289_));
 sg13g2_xnor2_1 _3895_ (.Y(_1290_),
    .A(net472),
    .B(_1271_));
 sg13g2_xnor2_1 _3896_ (.Y(_1291_),
    .A(_1389_),
    .B(_1270_));
 sg13g2_a21o_1 _3897_ (.A2(_1269_),
    .A1(\matt_venn_clock.sec_counter[8] ),
    .B1(net506),
    .X(_1292_));
 sg13g2_nand2_1 _3898_ (.Y(_1293_),
    .A(_1270_),
    .B(net507));
 sg13g2_xor2_1 _3899_ (.B(_1269_),
    .A(net537),
    .X(_1294_));
 sg13g2_nor2_1 _3900_ (.A(\matt_venn_clock.sec_counter[6] ),
    .B(\matt_venn_clock.sec_counter[7] ),
    .Y(_1295_));
 sg13g2_nand2_1 _3901_ (.Y(_1296_),
    .A(\matt_venn_clock.sec_counter[19] ),
    .B(\matt_venn_clock.sec_counter[24] ));
 sg13g2_and3_1 _3902_ (.X(_1297_),
    .A(\matt_venn_clock.sec_counter[13] ),
    .B(\matt_venn_clock.sec_counter[20] ),
    .C(\matt_venn_clock.sec_counter[21] ));
 sg13g2_nand4_1 _3903_ (.B(_1267_),
    .C(_1295_),
    .A(\matt_venn_clock.sec_counter[22] ),
    .Y(_1298_),
    .D(_1297_));
 sg13g2_nor4_2 _3904_ (.A(\matt_venn_clock.sec_counter[17] ),
    .B(_0054_),
    .C(_1296_),
    .Y(_1299_),
    .D(_1298_));
 sg13g2_nand3_1 _3905_ (.B(_1293_),
    .C(_1299_),
    .A(_1291_),
    .Y(_1300_));
 sg13g2_nor4_2 _3906_ (.A(_1289_),
    .B(_1290_),
    .C(_1294_),
    .Y(_1301_),
    .D(_1300_));
 sg13g2_nand3_1 _3907_ (.B(_1287_),
    .C(_1301_),
    .A(_1286_),
    .Y(_1302_));
 sg13g2_nor3_2 _3908_ (.A(_1283_),
    .B(_1285_),
    .C(_1302_),
    .Y(_1303_));
 sg13g2_xnor2_1 _3909_ (.Y(_1304_),
    .A(\clock_sec_u[0] ),
    .B(_1303_));
 sg13g2_nor3_2 _3910_ (.A(_1399_),
    .B(_0781_),
    .C(_1154_),
    .Y(_1305_));
 sg13g2_o21ai_1 _3911_ (.B1(net365),
    .Y(_1306_),
    .A1(net404),
    .A2(_1263_));
 sg13g2_a21oi_1 _3912_ (.A1(_1263_),
    .A2(_1304_),
    .Y(_0208_),
    .B1(_1306_));
 sg13g2_nor2_1 _3913_ (.A(_1303_),
    .B(_1305_),
    .Y(_1307_));
 sg13g2_nor3_1 _3914_ (.A(_1255_),
    .B(_1303_),
    .C(_1305_),
    .Y(_1308_));
 sg13g2_nand2_1 _3915_ (.Y(_1309_),
    .A(net479),
    .B(_1308_));
 sg13g2_nand2_1 _3916_ (.Y(_1310_),
    .A(\clock_sec_u[1] ),
    .B(\clock_sec_u[0] ));
 sg13g2_or2_1 _3917_ (.X(_1311_),
    .B(\clock_sec_u[0] ),
    .A(\clock_sec_u[1] ));
 sg13g2_nand3b_1 _3918_ (.B(_1310_),
    .C(_1311_),
    .Y(_1312_),
    .A_N(_1307_));
 sg13g2_a21oi_1 _3919_ (.A1(_1309_),
    .A2(_1312_),
    .Y(_0209_),
    .B1(net359));
 sg13g2_nor2_1 _3920_ (.A(_0046_),
    .B(_1310_),
    .Y(_1313_));
 sg13g2_xor2_1 _3921_ (.B(_1310_),
    .A(_0046_),
    .X(_1314_));
 sg13g2_o21ai_1 _3922_ (.B1(net365),
    .Y(_1315_),
    .A1(_1307_),
    .A2(_1314_));
 sg13g2_a21oi_1 _3923_ (.A1(_1349_),
    .A2(_1307_),
    .Y(_0210_),
    .B1(_1315_));
 sg13g2_nand2_1 _3924_ (.Y(_1316_),
    .A(net250),
    .B(_1308_));
 sg13g2_xnor2_1 _3925_ (.Y(_1317_),
    .A(_0041_),
    .B(_1313_));
 sg13g2_o21ai_1 _3926_ (.B1(_1317_),
    .Y(_1318_),
    .A1(_1303_),
    .A2(_1305_));
 sg13g2_a21oi_1 _3927_ (.A1(_1316_),
    .A2(_1318_),
    .Y(_0211_),
    .B1(net359));
 sg13g2_nor4_1 _3928_ (.A(\matt_venn_vga.x_block_q[5] ),
    .B(\matt_venn_vga.y_block_q[4] ),
    .C(\matt_venn_vga.y_block_q[3] ),
    .D(net414),
    .Y(_1319_));
 sg13g2_nor3_1 _3929_ (.A(\matt_venn_vga.font_0.dout[3] ),
    .B(\matt_venn_vga.col_index_q[0] ),
    .C(\matt_venn_vga.col_index_q[1] ),
    .Y(_1320_));
 sg13g2_o21ai_1 _3930_ (.B1(\matt_venn_vga.y_block_q[2] ),
    .Y(_1321_),
    .A1(\matt_venn_vga.y_block_q[1] ),
    .A2(\matt_venn_vga.y_block_q[0] ));
 sg13g2_o21ai_1 _3931_ (.B1(\matt_venn_vga.col_index_q[0] ),
    .Y(_1322_),
    .A1(_1406_),
    .A2(\matt_venn_vga.col_index_q[1] ));
 sg13g2_nand2_1 _3932_ (.Y(_1323_),
    .A(_1321_),
    .B(_1322_));
 sg13g2_o21ai_1 _3933_ (.B1(net415),
    .Y(_1324_),
    .A1(\matt_venn_vga.font_0.dout[1] ),
    .A2(_1407_));
 sg13g2_nor3_2 _3934_ (.A(_1320_),
    .B(_1323_),
    .C(net416),
    .Y(_0212_));
 sg13g2_nand2b_1 _3935_ (.Y(_1325_),
    .B(net363),
    .A_N(_1303_));
 sg13g2_inv_1 _3936_ (.Y(_1326_),
    .A(net282));
 sg13g2_and2_1 _3937_ (.A(net224),
    .B(_1326_),
    .X(_0213_));
 sg13g2_xnor2_1 _3938_ (.Y(_1327_),
    .A(\matt_venn_clock.sec_counter[0] ),
    .B(net371));
 sg13g2_nor2_1 _3939_ (.A(net280),
    .B(net372),
    .Y(_0214_));
 sg13g2_a21oi_1 _3940_ (.A1(\matt_venn_clock.sec_counter[0] ),
    .A2(\matt_venn_clock.sec_counter[1] ),
    .Y(_1328_),
    .B1(net240));
 sg13g2_nor3_1 _3941_ (.A(_1264_),
    .B(net280),
    .C(net241),
    .Y(_0215_));
 sg13g2_nor2_1 _3942_ (.A(net252),
    .B(_1264_),
    .Y(_1329_));
 sg13g2_nor3_1 _3943_ (.A(_1265_),
    .B(net280),
    .C(net253),
    .Y(_0216_));
 sg13g2_nor2_1 _3944_ (.A(net246),
    .B(_1265_),
    .Y(_1330_));
 sg13g2_nor3_1 _3945_ (.A(_1266_),
    .B(net280),
    .C(net247),
    .Y(_0217_));
 sg13g2_nor2_1 _3946_ (.A(net264),
    .B(_1266_),
    .Y(_1331_));
 sg13g2_nor3_1 _3947_ (.A(_1267_),
    .B(net280),
    .C(_1331_),
    .Y(_0218_));
 sg13g2_nor2_1 _3948_ (.A(net270),
    .B(_1267_),
    .Y(_1332_));
 sg13g2_nor3_1 _3949_ (.A(_1268_),
    .B(net280),
    .C(_1332_),
    .Y(_0219_));
 sg13g2_nor2_1 _3950_ (.A(net275),
    .B(_1268_),
    .Y(_1333_));
 sg13g2_nor3_1 _3951_ (.A(_1269_),
    .B(net280),
    .C(_1333_),
    .Y(_0220_));
 sg13g2_and2_1 _3952_ (.A(_1294_),
    .B(_1326_),
    .X(_0221_));
 sg13g2_nor2_1 _3953_ (.A(_1293_),
    .B(net282),
    .Y(_0222_));
 sg13g2_nor2_1 _3954_ (.A(net499),
    .B(net282),
    .Y(_0223_));
 sg13g2_nor2_1 _3955_ (.A(net473),
    .B(net280),
    .Y(_0224_));
 sg13g2_nor2_1 _3956_ (.A(_1289_),
    .B(net281),
    .Y(_0225_));
 sg13g2_xnor2_1 _3957_ (.Y(_1334_),
    .A(\matt_venn_clock.sec_counter[13] ),
    .B(_1288_));
 sg13g2_nor2_1 _3958_ (.A(net281),
    .B(net413),
    .Y(_0226_));
 sg13g2_and2_1 _3959_ (.A(net505),
    .B(_1326_),
    .X(_0227_));
 sg13g2_nor2_1 _3960_ (.A(net471),
    .B(net281),
    .Y(_0228_));
 sg13g2_nor2_1 _3961_ (.A(_1285_),
    .B(net281),
    .Y(_0229_));
 sg13g2_o21ai_1 _3962_ (.B1(net362),
    .Y(_1335_),
    .A1(net476),
    .A2(_1278_));
 sg13g2_nor2b_1 _3963_ (.A(net477),
    .B_N(_1279_),
    .Y(_0230_));
 sg13g2_and2_1 _3964_ (.A(net378),
    .B(_1274_),
    .X(_1336_));
 sg13g2_nor2_1 _3965_ (.A(net378),
    .B(_1279_),
    .Y(_1337_));
 sg13g2_nor3_1 _3966_ (.A(net282),
    .B(net379),
    .C(_1337_),
    .Y(_0231_));
 sg13g2_xnor2_1 _3967_ (.Y(_1338_),
    .A(net384),
    .B(_1337_));
 sg13g2_nor2_1 _3968_ (.A(net281),
    .B(net385),
    .Y(_0232_));
 sg13g2_xnor2_1 _3969_ (.Y(_1339_),
    .A(net423),
    .B(_1276_));
 sg13g2_nor2_1 _3970_ (.A(net281),
    .B(net424),
    .Y(_0233_));
 sg13g2_a21oi_1 _3971_ (.A1(\matt_venn_clock.sec_counter[20] ),
    .A2(_1276_),
    .Y(_1340_),
    .B1(net260));
 sg13g2_nor3_1 _3972_ (.A(_1280_),
    .B(net281),
    .C(net261),
    .Y(_0234_));
 sg13g2_xnor2_1 _3973_ (.Y(_1341_),
    .A(net386),
    .B(_1280_));
 sg13g2_nor2_1 _3974_ (.A(net281),
    .B(net387),
    .Y(_0235_));
 sg13g2_and2_1 _3975_ (.A(net363),
    .B(_1283_),
    .X(_0236_));
 sg13g2_xor2_1 _3976_ (.B(_1282_),
    .A(net420),
    .X(_1342_));
 sg13g2_nor2_1 _3977_ (.A(net282),
    .B(net421),
    .Y(_0237_));
 sg13g2_and2_1 _3978_ (.A(net366),
    .B(_0503_),
    .X(_0238_));
 sg13g2_and2_1 _3979_ (.A(net363),
    .B(_0580_),
    .X(_0239_));
 sg13g2_and2_1 _3980_ (.A(net363),
    .B(_0579_),
    .X(_0240_));
 sg13g2_nor3_1 _3981_ (.A(net360),
    .B(_1441_),
    .C(_1606_),
    .Y(_0241_));
 sg13g2_and2_1 _3982_ (.A(net363),
    .B(_0577_),
    .X(_0242_));
 sg13g2_and2_1 _3983_ (.A(net363),
    .B(_0591_),
    .X(_0243_));
 sg13g2_and2_1 _3984_ (.A(net363),
    .B(_0601_),
    .X(_0244_));
 sg13g2_nor4_1 _3985_ (.A(\matt_venn_vga_shadow.x_block_q[5] ),
    .B(\matt_venn_vga_shadow.y_block_q[4] ),
    .C(\matt_venn_vga_shadow.y_block_q[3] ),
    .D(\matt_venn_vga_shadow.y_block_q[5] ),
    .Y(_1343_));
 sg13g2_nor3_1 _3986_ (.A(\matt_venn_vga_shadow.font_0.dout[3] ),
    .B(\matt_venn_vga_shadow.col_index_q[0] ),
    .C(\matt_venn_vga_shadow.col_index_q[1] ),
    .Y(_1344_));
 sg13g2_o21ai_1 _3987_ (.B1(net466),
    .Y(_1345_),
    .A1(\matt_venn_vga_shadow.y_block_q[1] ),
    .A2(\matt_venn_vga_shadow.y_block_q[0] ));
 sg13g2_o21ai_1 _3988_ (.B1(\matt_venn_vga_shadow.col_index_q[0] ),
    .Y(_1346_),
    .A1(_1408_),
    .A2(\matt_venn_vga_shadow.col_index_q[1] ));
 sg13g2_nand2_1 _3989_ (.Y(_1347_),
    .A(net467),
    .B(_1346_));
 sg13g2_o21ai_1 _3990_ (.B1(_1343_),
    .Y(_1348_),
    .A1(\matt_venn_vga_shadow.font_0.dout[1] ),
    .A2(_1409_));
 sg13g2_nor3_2 _3991_ (.A(_1344_),
    .B(net468),
    .C(_1348_),
    .Y(_0245_));
 sg13g2_or2_1 _3992_ (.X(_0247_),
    .B(_0503_),
    .A(net316));
 sg13g2_nor2_1 _3993_ (.A(net360),
    .B(_0520_),
    .Y(_0248_));
 sg13g2_and2_1 _3994_ (.A(net362),
    .B(_0649_),
    .X(_0249_));
 sg13g2_and2_1 _3995_ (.A(net362),
    .B(_0647_),
    .X(_0250_));
 sg13g2_and2_1 _3996_ (.A(net362),
    .B(_0645_),
    .X(_0251_));
 sg13g2_and2_1 _3997_ (.A(net362),
    .B(_0643_),
    .X(_0252_));
 sg13g2_nor2_1 _3998_ (.A(net360),
    .B(_0660_),
    .Y(_0253_));
 sg13g2_and2_1 _3999_ (.A(net362),
    .B(_0671_),
    .X(_0254_));
 sg13g2_dfrbp_1 _4000_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net15),
    .D(_0079_),
    .Q_N(_1966_),
    .Q(\matt_venn_vga.color[0] ));
 sg13g2_dfrbp_1 _4001_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net16),
    .D(_0080_),
    .Q_N(_1967_),
    .Q(\matt_venn_vga.color[1] ));
 sg13g2_dfrbp_1 _4002_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net17),
    .D(_0000_),
    .Q_N(_1968_),
    .Q(\matt_venn_vga.digit_0.digit_index[0] ));
 sg13g2_dfrbp_1 _4003_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net18),
    .D(_0001_),
    .Q_N(_1969_),
    .Q(\matt_venn_vga.digit_0.digit_index[1] ));
 sg13g2_dfrbp_1 _4004_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net19),
    .D(_0002_),
    .Q_N(_1970_),
    .Q(\matt_venn_vga.digit_0.digit_index[2] ));
 sg13g2_dfrbp_1 _4005_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net20),
    .D(_0003_),
    .Q_N(_1971_),
    .Q(\matt_venn_vga.digit_0.digit_index[3] ));
 sg13g2_dfrbp_1 _4006_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net21),
    .D(_0004_),
    .Q_N(_1972_),
    .Q(\matt_venn_vga.digit_0.digit_index[4] ));
 sg13g2_dfrbp_1 _4007_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net22),
    .D(_0005_),
    .Q_N(_1973_),
    .Q(\matt_venn_vga.digit_0.digit_index[5] ));
 sg13g2_dfrbp_1 _4008_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net23),
    .D(_0011_),
    .Q_N(_1974_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[0] ));
 sg13g2_dfrbp_1 _4009_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net24),
    .D(_0012_),
    .Q_N(_1975_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[1] ));
 sg13g2_dfrbp_1 _4010_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net25),
    .D(_0013_),
    .Q_N(_1976_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[2] ));
 sg13g2_dfrbp_1 _4011_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net26),
    .D(_0014_),
    .Q_N(_1977_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[3] ));
 sg13g2_dfrbp_1 _4012_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net27),
    .D(_0015_),
    .Q_N(_1978_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[4] ));
 sg13g2_dfrbp_1 _4013_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net28),
    .D(_0016_),
    .Q_N(_1979_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[5] ));
 sg13g2_dfrbp_1 _4014_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net29),
    .D(_0017_),
    .Q_N(_1980_),
    .Q(\matt_venn_vga_shadow.color[4] ));
 sg13g2_dfrbp_1 _4015_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net30),
    .D(_0018_),
    .Q_N(_1981_),
    .Q(\matt_venn_vga_shadow.color[5] ));
 sg13g2_dfrbp_1 _4016_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net31),
    .D(_0008_),
    .Q_N(_1982_),
    .Q(\matt_venn_vga.font_0.dout[1] ));
 sg13g2_dfrbp_1 _4017_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net75),
    .D(_0009_),
    .Q_N(_1983_),
    .Q(\matt_venn_vga.font_0.dout[2] ));
 sg13g2_dfrbp_1 _4018_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net123),
    .D(_0010_),
    .Q_N(_1965_),
    .Q(\matt_venn_vga.font_0.dout[3] ));
 sg13g2_dfrbp_1 _4019_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net122),
    .D(net269),
    .Q_N(_0049_),
    .Q(\ydelta[0] ));
 sg13g2_dfrbp_1 _4020_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net120),
    .D(_0082_),
    .Q_N(_1964_),
    .Q(\ydelta[1] ));
 sg13g2_dfrbp_1 _4021_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net118),
    .D(_0083_),
    .Q_N(_1963_),
    .Q(\ydelta[2] ));
 sg13g2_dfrbp_1 _4022_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net117),
    .D(_0084_),
    .Q_N(_1962_),
    .Q(\ydelta[3] ));
 sg13g2_dfrbp_1 _4023_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net115),
    .D(_0085_),
    .Q_N(_1961_),
    .Q(\ydelta[4] ));
 sg13g2_dfrbp_1 _4024_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net114),
    .D(_0086_),
    .Q_N(_1960_),
    .Q(\ydelta[5] ));
 sg13g2_dfrbp_1 _4025_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net112),
    .D(net442),
    .Q_N(_1959_),
    .Q(\ydelta[6] ));
 sg13g2_dfrbp_1 _4026_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net111),
    .D(net408),
    .Q_N(_0058_),
    .Q(\ydelta[7] ));
 sg13g2_dfrbp_1 _4027_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net109),
    .D(_0089_),
    .Q_N(_0078_),
    .Q(\pxm[0] ));
 sg13g2_dfrbp_1 _4028_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net108),
    .D(_0090_),
    .Q_N(_1958_),
    .Q(\pxm[1] ));
 sg13g2_dfrbp_1 _4029_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net106),
    .D(_0091_),
    .Q_N(_0050_),
    .Q(\px[0] ));
 sg13g2_dfrbp_1 _4030_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net105),
    .D(_0092_),
    .Q_N(_1957_),
    .Q(\px[1] ));
 sg13g2_dfrbp_1 _4031_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net103),
    .D(_0093_),
    .Q_N(_1956_),
    .Q(\px[2] ));
 sg13g2_dfrbp_1 _4032_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net101),
    .D(_0094_),
    .Q_N(_1955_),
    .Q(\px[3] ));
 sg13g2_dfrbp_1 _4033_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net99),
    .D(_0095_),
    .Q_N(_1954_),
    .Q(\px[4] ));
 sg13g2_dfrbp_1 _4034_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net95),
    .D(_0096_),
    .Q_N(_1953_),
    .Q(\px[5] ));
 sg13g2_dfrbp_1 _4035_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net93),
    .D(_0097_),
    .Q_N(_1952_),
    .Q(\px[6] ));
 sg13g2_dfrbp_1 _4036_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net91),
    .D(_0098_),
    .Q_N(_0028_),
    .Q(\px[7] ));
 sg13g2_dfrbp_1 _4037_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net89),
    .D(_0099_),
    .Q_N(_1951_),
    .Q(\px[8] ));
 sg13g2_dfrbp_1 _4038_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net87),
    .D(_0100_),
    .Q_N(_1950_),
    .Q(\px[9] ));
 sg13g2_dfrbp_1 _4039_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net85),
    .D(net502),
    .Q_N(_1949_),
    .Q(\py[0] ));
 sg13g2_dfrbp_1 _4040_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net83),
    .D(_0102_),
    .Q_N(_0063_),
    .Q(\py[1] ));
 sg13g2_dfrbp_1 _4041_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net81),
    .D(_0103_),
    .Q_N(_0062_),
    .Q(\py[2] ));
 sg13g2_dfrbp_1 _4042_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net79),
    .D(_0104_),
    .Q_N(_0027_),
    .Q(\py[3] ));
 sg13g2_dfrbp_1 _4043_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net74),
    .D(_0105_),
    .Q_N(_0061_),
    .Q(\py[4] ));
 sg13g2_dfrbp_1 _4044_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net72),
    .D(_0106_),
    .Q_N(_0060_),
    .Q(\py[5] ));
 sg13g2_dfrbp_1 _4045_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net70),
    .D(_0107_),
    .Q_N(_0059_),
    .Q(\py[6] ));
 sg13g2_dfrbp_1 _4046_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net68),
    .D(_0108_),
    .Q_N(_0064_),
    .Q(\py[7] ));
 sg13g2_dfrbp_1 _4047_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net66),
    .D(_0109_),
    .Q_N(_0024_),
    .Q(\py[8] ));
 sg13g2_dfrbp_1 _4048_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net64),
    .D(_0110_),
    .Q_N(_0022_),
    .Q(\py[9] ));
 sg13g2_dfrbp_1 _4049_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net62),
    .D(_0111_),
    .Q_N(_1948_),
    .Q(\pym[10] ));
 sg13g2_dfrbp_1 _4050_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net60),
    .D(_0112_),
    .Q_N(_1947_),
    .Q(\pym[11] ));
 sg13g2_dfrbp_1 _4051_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net58),
    .D(_0113_),
    .Q_N(_0077_),
    .Q(\t[0] ));
 sg13g2_dfrbp_1 _4052_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net57),
    .D(net465),
    .Q_N(_1946_),
    .Q(\t[1] ));
 sg13g2_dfrbp_1 _4053_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net55),
    .D(net457),
    .Q_N(_1945_),
    .Q(\t[2] ));
 sg13g2_dfrbp_1 _4054_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net54),
    .D(net279),
    .Q_N(_1944_),
    .Q(\t[3] ));
 sg13g2_dfrbp_1 _4055_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net52),
    .D(_0117_),
    .Q_N(_1943_),
    .Q(\product_comp[0] ));
 sg13g2_dfrbp_1 _4056_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net51),
    .D(_0118_),
    .Q_N(_1942_),
    .Q(\product_comp[1] ));
 sg13g2_dfrbp_1 _4057_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net49),
    .D(_0119_),
    .Q_N(_1941_),
    .Q(\product_comp[2] ));
 sg13g2_dfrbp_1 _4058_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net48),
    .D(_0120_),
    .Q_N(_1940_),
    .Q(\product_comp[3] ));
 sg13g2_dfrbp_1 _4059_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net46),
    .D(net486),
    .Q_N(_0037_),
    .Q(\product_comp[4] ));
 sg13g2_dfrbp_1 _4060_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net45),
    .D(_0122_),
    .Q_N(_0036_),
    .Q(\product_comp[5] ));
 sg13g2_dfrbp_1 _4061_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net43),
    .D(net440),
    .Q_N(_0035_),
    .Q(\product_comp[6] ));
 sg13g2_dfrbp_1 _4062_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net41),
    .D(_0124_),
    .Q_N(_1939_),
    .Q(\product_comp[7] ));
 sg13g2_dfrbp_1 _4063_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net39),
    .D(_0125_),
    .Q_N(_0034_),
    .Q(\product_comp[8] ));
 sg13g2_dfrbp_1 _4064_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net37),
    .D(_0126_),
    .Q_N(_0033_),
    .Q(\product_comp[9] ));
 sg13g2_dfrbp_1 _4065_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net35),
    .D(_0127_),
    .Q_N(_0065_),
    .Q(\product_comp[10] ));
 sg13g2_dfrbp_1 _4066_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net76),
    .D(_0128_),
    .Q_N(_1984_),
    .Q(dx));
 sg13g2_dfrbp_1 _4067_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net77),
    .D(_0019_),
    .Q_N(_1985_),
    .Q(\matt_venn_vga_shadow.font_0.dout[1] ));
 sg13g2_dfrbp_1 _4068_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net96),
    .D(_0020_),
    .Q_N(_1986_),
    .Q(\matt_venn_vga_shadow.font_0.dout[2] ));
 sg13g2_dfrbp_1 _4069_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net33),
    .D(_0021_),
    .Q_N(_1938_),
    .Q(\matt_venn_vga_shadow.font_0.dout[3] ));
 sg13g2_dfrbp_1 _4070_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net14),
    .D(_0129_),
    .Q_N(_1937_),
    .Q(\matt_venn_vga.color[2] ));
 sg13g2_dfrbp_1 _4071_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net13),
    .D(_0130_),
    .Q_N(_1936_),
    .Q(\matt_venn_vga_shadow.color[0] ));
 sg13g2_dfrbp_1 _4072_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net214),
    .D(_0131_),
    .Q_N(_1935_),
    .Q(\matt_venn_vga_shadow.color[1] ));
 sg13g2_dfrbp_1 _4073_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net213),
    .D(_0132_),
    .Q_N(_1934_),
    .Q(\matt_venn_vga_shadow.color[3] ));
 sg13g2_dfrbp_1 _4074_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net212),
    .D(_0133_),
    .Q_N(_0070_),
    .Q(\vga_sync.hsync ));
 sg13g2_dfrbp_1 _4075_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net211),
    .D(_0134_),
    .Q_N(_1933_),
    .Q(\matt_venn_vga.y_px[0] ));
 sg13g2_dfrbp_1 _4076_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net209),
    .D(_0135_),
    .Q_N(_0031_),
    .Q(\matt_venn_vga.y_px[1] ));
 sg13g2_dfrbp_1 _4077_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net207),
    .D(_0136_),
    .Q_N(_0030_),
    .Q(\matt_venn_vga.y_px[2] ));
 sg13g2_dfrbp_1 _4078_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net205),
    .D(_0137_),
    .Q_N(_0032_),
    .Q(\matt_venn_vga.y_px[3] ));
 sg13g2_dfrbp_1 _4079_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net203),
    .D(_0138_),
    .Q_N(_0026_),
    .Q(\matt_venn_vga.y_px[4] ));
 sg13g2_dfrbp_1 _4080_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net199),
    .D(net530),
    .Q_N(_0069_),
    .Q(\matt_venn_vga.y_px[5] ));
 sg13g2_dfrbp_1 _4081_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net197),
    .D(_0140_),
    .Q_N(_0029_),
    .Q(\matt_venn_vga.y_px[6] ));
 sg13g2_dfrbp_1 _4082_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net195),
    .D(_0141_),
    .Q_N(_0025_),
    .Q(\matt_venn_vga.y_px[7] ));
 sg13g2_dfrbp_1 _4083_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net193),
    .D(_0142_),
    .Q_N(_0023_),
    .Q(\matt_venn_vga.y_px[8] ));
 sg13g2_dfrbp_1 _4084_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net191),
    .D(_0143_),
    .Q_N(_0057_),
    .Q(\matt_venn_vga.y_px[9] ));
 sg13g2_dfrbp_1 _4085_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net189),
    .D(_0144_),
    .Q_N(_1932_),
    .Q(\vga_sync.vsync ));
 sg13g2_dfrbp_1 _4086_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net188),
    .D(_0145_),
    .Q_N(_1931_),
    .Q(\matt_venn_vga_shadow.col_index[0] ));
 sg13g2_dfrbp_1 _4087_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net97),
    .D(_0146_),
    .Q_N(_1987_),
    .Q(\matt_venn_vga_shadow.col_index[1] ));
 sg13g2_dfrbp_1 _4088_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net184),
    .D(_0006_),
    .Q_N(_1988_),
    .Q(\matt_venn_vga.color[4] ));
 sg13g2_dfrbp_1 _4089_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net187),
    .D(_0007_),
    .Q_N(_1930_),
    .Q(\matt_venn_vga.color[5] ));
 sg13g2_dfrbp_1 _4090_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net186),
    .D(_0147_),
    .Q_N(_1929_),
    .Q(\matt_venn_vga.color[3] ));
 sg13g2_dfrbp_1 _4091_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net183),
    .D(_0148_),
    .Q_N(_1928_),
    .Q(\matt_venn_vga_shadow.color[2] ));
 sg13g2_dfrbp_1 _4092_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net182),
    .D(_0149_),
    .Q_N(_0076_),
    .Q(\h[0] ));
 sg13g2_dfrbp_1 _4093_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net181),
    .D(_0150_),
    .Q_N(_1927_),
    .Q(\h[1] ));
 sg13g2_dfrbp_1 _4094_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net180),
    .D(_0151_),
    .Q_N(_1926_),
    .Q(\h[2] ));
 sg13g2_dfrbp_1 _4095_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net179),
    .D(_0152_),
    .Q_N(_1925_),
    .Q(\h[3] ));
 sg13g2_dfrbp_1 _4096_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net178),
    .D(_0153_),
    .Q_N(_1924_),
    .Q(\h[4] ));
 sg13g2_dfrbp_1 _4097_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net177),
    .D(_0154_),
    .Q_N(_1923_),
    .Q(\h[5] ));
 sg13g2_dfrbp_1 _4098_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net176),
    .D(_0155_),
    .Q_N(\matt_venn_vga.digit_0.char[0] ),
    .Q(\matt_venn_vga.x_px[6] ));
 sg13g2_dfrbp_1 _4099_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net175),
    .D(_0156_),
    .Q_N(_1922_),
    .Q(\matt_venn_vga.x_px[7] ));
 sg13g2_dfrbp_1 _4100_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net174),
    .D(_0157_),
    .Q_N(_0055_),
    .Q(\matt_venn_vga.x_px[8] ));
 sg13g2_dfrbp_1 _4101_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net173),
    .D(_0158_),
    .Q_N(_1921_),
    .Q(\matt_venn_vga.x_px[9] ));
 sg13g2_dfrbp_1 _4102_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net172),
    .D(_0159_),
    .Q_N(_1920_),
    .Q(\matt_venn_clock.pulse_hrs.comp[0] ));
 sg13g2_dfrbp_1 _4103_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net170),
    .D(_0160_),
    .Q_N(_1919_),
    .Q(\matt_venn_clock.pulse_hrs.comp[1] ));
 sg13g2_dfrbp_1 _4104_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net168),
    .D(net452),
    .Q_N(_1918_),
    .Q(\matt_venn_clock.pulse_hrs.comp[2] ));
 sg13g2_dfrbp_1 _4105_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net166),
    .D(net433),
    .Q_N(_1917_),
    .Q(\matt_venn_clock.pulse_hrs.comp[3] ));
 sg13g2_dfrbp_1 _4106_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net164),
    .D(_0163_),
    .Q_N(_1916_),
    .Q(\matt_venn_clock.pulse_hrs.comp[4] ));
 sg13g2_dfrbp_1 _4107_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net162),
    .D(_0164_),
    .Q_N(_1915_),
    .Q(\matt_venn_clock.pulse_hrs.count[0] ));
 sg13g2_dfrbp_1 _4108_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net160),
    .D(net497),
    .Q_N(_1914_),
    .Q(\matt_venn_clock.pulse_hrs.count[1] ));
 sg13g2_dfrbp_1 _4109_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net158),
    .D(net401),
    .Q_N(_1913_),
    .Q(\matt_venn_clock.pulse_hrs.count[2] ));
 sg13g2_dfrbp_1 _4110_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net156),
    .D(net445),
    .Q_N(_1912_),
    .Q(\matt_venn_clock.pulse_hrs.count[3] ));
 sg13g2_dfrbp_1 _4111_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net154),
    .D(net266),
    .Q_N(_0068_),
    .Q(\matt_venn_clock.pulse_hrs.count[4] ));
 sg13g2_dfrbp_1 _4112_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0169_),
    .Q_N(_1911_),
    .Q(\matt_venn_clock.pulse_min.comp[0] ));
 sg13g2_dfrbp_1 _4113_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net150),
    .D(_0170_),
    .Q_N(_1910_),
    .Q(\matt_venn_clock.pulse_min.comp[1] ));
 sg13g2_dfrbp_1 _4114_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net148),
    .D(_0171_),
    .Q_N(_1909_),
    .Q(\matt_venn_clock.pulse_min.comp[2] ));
 sg13g2_dfrbp_1 _4115_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net146),
    .D(net460),
    .Q_N(_1908_),
    .Q(\matt_venn_clock.pulse_min.comp[3] ));
 sg13g2_dfrbp_1 _4116_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net144),
    .D(_0173_),
    .Q_N(_1907_),
    .Q(\matt_venn_clock.pulse_min.comp[4] ));
 sg13g2_dfrbp_1 _4117_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net142),
    .D(_0174_),
    .Q_N(_1906_),
    .Q(\matt_venn_clock.pulse_min.count[0] ));
 sg13g2_dfrbp_1 _4118_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net140),
    .D(net455),
    .Q_N(_1905_),
    .Q(\matt_venn_clock.pulse_min.count[1] ));
 sg13g2_dfrbp_1 _4119_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net138),
    .D(_0176_),
    .Q_N(_1904_),
    .Q(\matt_venn_clock.pulse_min.count[2] ));
 sg13g2_dfrbp_1 _4120_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net136),
    .D(net277),
    .Q_N(_1903_),
    .Q(\matt_venn_clock.pulse_min.count[3] ));
 sg13g2_dfrbp_1 _4121_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net134),
    .D(net257),
    .Q_N(_0067_),
    .Q(\matt_venn_clock.pulse_min.count[4] ));
 sg13g2_dfrbp_1 _4122_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net132),
    .D(_0179_),
    .Q_N(_1902_),
    .Q(\matt_venn_clock.pulse_sec.comp[0] ));
 sg13g2_dfrbp_1 _4123_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net130),
    .D(_0180_),
    .Q_N(_1901_),
    .Q(\matt_venn_clock.pulse_sec.comp[1] ));
 sg13g2_dfrbp_1 _4124_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net128),
    .D(_0181_),
    .Q_N(_1900_),
    .Q(\matt_venn_clock.pulse_sec.comp[2] ));
 sg13g2_dfrbp_1 _4125_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net126),
    .D(_0182_),
    .Q_N(_1899_),
    .Q(\matt_venn_clock.pulse_sec.comp[3] ));
 sg13g2_dfrbp_1 _4126_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net124),
    .D(net274),
    .Q_N(_1898_),
    .Q(\matt_venn_clock.pulse_sec.comp[4] ));
 sg13g2_dfrbp_1 _4127_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net119),
    .D(_0184_),
    .Q_N(_1897_),
    .Q(\matt_venn_clock.pulse_sec.count[0] ));
 sg13g2_dfrbp_1 _4128_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net116),
    .D(net484),
    .Q_N(_1896_),
    .Q(\matt_venn_clock.pulse_sec.count[1] ));
 sg13g2_dfrbp_1 _4129_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net113),
    .D(net428),
    .Q_N(_1895_),
    .Q(\matt_venn_clock.pulse_sec.count[2] ));
 sg13g2_dfrbp_1 _4130_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net110),
    .D(net249),
    .Q_N(_1894_),
    .Q(\matt_venn_clock.pulse_sec.count[3] ));
 sg13g2_dfrbp_1 _4131_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net107),
    .D(net244),
    .Q_N(_0066_),
    .Q(\matt_venn_clock.pulse_sec.count[4] ));
 sg13g2_dfrbp_1 _4132_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net104),
    .D(net229),
    .Q_N(_0075_),
    .Q(\clock_color_offset[0] ));
 sg13g2_dfrbp_1 _4133_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net100),
    .D(_0190_),
    .Q_N(_0056_),
    .Q(\clock_color_offset[1] ));
 sg13g2_dfrbp_1 _4134_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net94),
    .D(net426),
    .Q_N(_1893_),
    .Q(\clock_color_offset[2] ));
 sg13g2_dfrbp_1 _4135_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net90),
    .D(net232),
    .Q_N(_0074_),
    .Q(\clock_hrs_d[0] ));
 sg13g2_dfrbp_1 _4136_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net86),
    .D(_0193_),
    .Q_N(_0047_),
    .Q(\clock_hrs_d[1] ));
 sg13g2_dfrbp_1 _4137_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net82),
    .D(_0194_),
    .Q_N(_0052_),
    .Q(\clock_hrs_u[0] ));
 sg13g2_dfrbp_1 _4138_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net78),
    .D(_0195_),
    .Q_N(_0048_),
    .Q(\clock_hrs_u[1] ));
 sg13g2_dfrbp_1 _4139_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net71),
    .D(net462),
    .Q_N(_0042_),
    .Q(\clock_hrs_u[2] ));
 sg13g2_dfrbp_1 _4140_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net67),
    .D(_0197_),
    .Q_N(_0039_),
    .Q(\clock_hrs_u[3] ));
 sg13g2_dfrbp_1 _4141_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net63),
    .D(net236),
    .Q_N(_0073_),
    .Q(\clock_min_d[0] ));
 sg13g2_dfrbp_1 _4142_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net59),
    .D(net511),
    .Q_N(_1892_),
    .Q(\clock_min_d[1] ));
 sg13g2_dfrbp_1 _4143_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net56),
    .D(net411),
    .Q_N(_0043_),
    .Q(\clock_min_d[2] ));
 sg13g2_dfrbp_1 _4144_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net53),
    .D(net398),
    .Q_N(_0051_),
    .Q(\clock_min_u[0] ));
 sg13g2_dfrbp_1 _4145_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net50),
    .D(_0202_),
    .Q_N(_1891_),
    .Q(\clock_min_u[1] ));
 sg13g2_dfrbp_1 _4146_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net47),
    .D(net488),
    .Q_N(_0044_),
    .Q(\clock_min_u[2] ));
 sg13g2_dfrbp_1 _4147_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net44),
    .D(net239),
    .Q_N(_0040_),
    .Q(\clock_min_u[3] ));
 sg13g2_dfrbp_1 _4148_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net40),
    .D(net272),
    .Q_N(_0072_),
    .Q(\clock_sec_d[0] ));
 sg13g2_dfrbp_1 _4149_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net36),
    .D(net527),
    .Q_N(_1890_),
    .Q(\clock_sec_d[1] ));
 sg13g2_dfrbp_1 _4150_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net32),
    .D(net394),
    .Q_N(_0045_),
    .Q(\clock_sec_d[2] ));
 sg13g2_dfrbp_1 _4151_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net208),
    .D(net405),
    .Q_N(_0038_),
    .Q(\clock_sec_u[0] ));
 sg13g2_dfrbp_1 _4152_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net204),
    .D(net480),
    .Q_N(_1889_),
    .Q(\clock_sec_u[1] ));
 sg13g2_dfrbp_1 _4153_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net198),
    .D(net259),
    .Q_N(_0046_),
    .Q(\clock_sec_u[2] ));
 sg13g2_dfrbp_1 _4154_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net194),
    .D(net251),
    .Q_N(_0041_),
    .Q(\clock_sec_u[3] ));
 sg13g2_dfrbp_1 _4155_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net190),
    .D(net417),
    .Q_N(_1888_),
    .Q(\matt_venn_vga.draw ));
 sg13g2_dfrbp_1 _4156_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net171),
    .D(_0213_),
    .Q_N(_0071_),
    .Q(\matt_venn_clock.sec_counter[0] ));
 sg13g2_dfrbp_1 _4157_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net169),
    .D(_0214_),
    .Q_N(_1887_),
    .Q(\matt_venn_clock.sec_counter[1] ));
 sg13g2_dfrbp_1 _4158_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net167),
    .D(net242),
    .Q_N(_1886_),
    .Q(\matt_venn_clock.sec_counter[2] ));
 sg13g2_dfrbp_1 _4159_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net165),
    .D(_0216_),
    .Q_N(_1885_),
    .Q(\matt_venn_clock.sec_counter[3] ));
 sg13g2_dfrbp_1 _4160_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net163),
    .D(_0217_),
    .Q_N(_1884_),
    .Q(\matt_venn_clock.sec_counter[4] ));
 sg13g2_dfrbp_1 _4161_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net161),
    .D(_0218_),
    .Q_N(_1883_),
    .Q(\matt_venn_clock.sec_counter[5] ));
 sg13g2_dfrbp_1 _4162_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net159),
    .D(_0219_),
    .Q_N(_1882_),
    .Q(\matt_venn_clock.sec_counter[6] ));
 sg13g2_dfrbp_1 _4163_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net157),
    .D(_0220_),
    .Q_N(_1881_),
    .Q(\matt_venn_clock.sec_counter[7] ));
 sg13g2_dfrbp_1 _4164_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net155),
    .D(_0221_),
    .Q_N(_1880_),
    .Q(\matt_venn_clock.sec_counter[8] ));
 sg13g2_dfrbp_1 _4165_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net153),
    .D(_0222_),
    .Q_N(_1879_),
    .Q(\matt_venn_clock.sec_counter[9] ));
 sg13g2_dfrbp_1 _4166_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net151),
    .D(_0223_),
    .Q_N(_1878_),
    .Q(\matt_venn_clock.sec_counter[10] ));
 sg13g2_dfrbp_1 _4167_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net149),
    .D(_0224_),
    .Q_N(_1877_),
    .Q(\matt_venn_clock.sec_counter[11] ));
 sg13g2_dfrbp_1 _4168_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net147),
    .D(_0225_),
    .Q_N(_0053_),
    .Q(\matt_venn_clock.sec_counter[12] ));
 sg13g2_dfrbp_1 _4169_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net145),
    .D(_0226_),
    .Q_N(_1876_),
    .Q(\matt_venn_clock.sec_counter[13] ));
 sg13g2_dfrbp_1 _4170_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net143),
    .D(_0227_),
    .Q_N(_1875_),
    .Q(\matt_venn_clock.sec_counter[14] ));
 sg13g2_dfrbp_1 _4171_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net141),
    .D(_0228_),
    .Q_N(_1874_),
    .Q(\matt_venn_clock.sec_counter[15] ));
 sg13g2_dfrbp_1 _4172_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net139),
    .D(_0229_),
    .Q_N(_1873_),
    .Q(\matt_venn_clock.sec_counter[16] ));
 sg13g2_dfrbp_1 _4173_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net137),
    .D(_0230_),
    .Q_N(_1872_),
    .Q(\matt_venn_clock.sec_counter[17] ));
 sg13g2_dfrbp_1 _4174_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net135),
    .D(net380),
    .Q_N(_0054_),
    .Q(\matt_venn_clock.sec_counter[18] ));
 sg13g2_dfrbp_1 _4175_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net133),
    .D(_0232_),
    .Q_N(_1871_),
    .Q(\matt_venn_clock.sec_counter[19] ));
 sg13g2_dfrbp_1 _4176_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net131),
    .D(_0233_),
    .Q_N(_1870_),
    .Q(\matt_venn_clock.sec_counter[20] ));
 sg13g2_dfrbp_1 _4177_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net129),
    .D(net262),
    .Q_N(_1869_),
    .Q(\matt_venn_clock.sec_counter[21] ));
 sg13g2_dfrbp_1 _4178_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net127),
    .D(_0235_),
    .Q_N(_1868_),
    .Q(\matt_venn_clock.sec_counter[22] ));
 sg13g2_dfrbp_1 _4179_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net125),
    .D(_0236_),
    .Q_N(_1867_),
    .Q(\matt_venn_clock.sec_counter[23] ));
 sg13g2_dfrbp_1 _4180_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net185),
    .D(_0237_),
    .Q_N(_1989_),
    .Q(\matt_venn_clock.sec_counter[24] ));
 sg13g2_dfrbp_1 _4181_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net201),
    .D(net222),
    .Q_N(_1990_),
    .Q(\matt_venn_vga.col_index_q[0] ));
 sg13g2_dfrbp_1 _4182_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net121),
    .D(net220),
    .Q_N(_1866_),
    .Q(\matt_venn_vga.col_index_q[1] ));
 sg13g2_dfrbp_1 _4183_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net102),
    .D(_0238_),
    .Q_N(_1865_),
    .Q(\matt_venn_vga.x_block_q[5] ));
 sg13g2_dfrbp_1 _4184_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net98),
    .D(_0239_),
    .Q_N(_1864_),
    .Q(\matt_venn_vga.y_block_q[0] ));
 sg13g2_dfrbp_1 _4185_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net92),
    .D(_0240_),
    .Q_N(_1863_),
    .Q(\matt_venn_vga.y_block_q[1] ));
 sg13g2_dfrbp_1 _4186_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net88),
    .D(_0241_),
    .Q_N(_1862_),
    .Q(\matt_venn_vga.y_block_q[2] ));
 sg13g2_dfrbp_1 _4187_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net84),
    .D(_0242_),
    .Q_N(_1861_),
    .Q(\matt_venn_vga.y_block_q[3] ));
 sg13g2_dfrbp_1 _4188_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net80),
    .D(_0243_),
    .Q_N(_1860_),
    .Q(\matt_venn_vga.y_block_q[4] ));
 sg13g2_dfrbp_1 _4189_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net73),
    .D(_0244_),
    .Q_N(_1859_),
    .Q(\matt_venn_vga.y_block_q[5] ));
 sg13g2_dfrbp_1 _4190_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net69),
    .D(net469),
    .Q_N(_1858_),
    .Q(\matt_venn_vga_shadow.draw ));
 sg13g2_dfrbp_1 _4191_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net65),
    .D(_0246_),
    .Q_N(_1857_),
    .Q(\matt_venn_vga.col_index[0] ));
 sg13g2_dfrbp_1 _4192_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net202),
    .D(_0247_),
    .Q_N(_1991_),
    .Q(\matt_venn_vga.col_index[1] ));
 sg13g2_dfrbp_1 _4193_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net192),
    .D(net221),
    .Q_N(_1992_),
    .Q(\matt_venn_vga_shadow.col_index_q[0] ));
 sg13g2_dfrbp_1 _4194_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net61),
    .D(net223),
    .Q_N(_1856_),
    .Q(\matt_venn_vga_shadow.col_index_q[1] ));
 sg13g2_dfrbp_1 _4195_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net42),
    .D(_0248_),
    .Q_N(_1855_),
    .Q(\matt_venn_vga_shadow.x_block_q[5] ));
 sg13g2_dfrbp_1 _4196_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net38),
    .D(_0249_),
    .Q_N(_1854_),
    .Q(\matt_venn_vga_shadow.y_block_q[0] ));
 sg13g2_dfrbp_1 _4197_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net34),
    .D(_0250_),
    .Q_N(_1853_),
    .Q(\matt_venn_vga_shadow.y_block_q[1] ));
 sg13g2_dfrbp_1 _4198_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net210),
    .D(_0251_),
    .Q_N(_1852_),
    .Q(\matt_venn_vga_shadow.y_block_q[2] ));
 sg13g2_dfrbp_1 _4199_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net206),
    .D(_0252_),
    .Q_N(_1851_),
    .Q(\matt_venn_vga_shadow.y_block_q[3] ));
 sg13g2_dfrbp_1 _4200_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net200),
    .D(_0253_),
    .Q_N(_1850_),
    .Q(\matt_venn_vga_shadow.y_block_q[4] ));
 sg13g2_dfrbp_1 _4201_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net196),
    .D(_0254_),
    .Q_N(_1849_),
    .Q(\matt_venn_vga_shadow.y_block_q[5] ));
 sg13g2_tiehi _4070__14 (.L_HI(net14));
 sg13g2_tiehi _4000__15 (.L_HI(net15));
 sg13g2_tiehi _4001__16 (.L_HI(net16));
 sg13g2_tiehi _4002__17 (.L_HI(net17));
 sg13g2_tiehi _4003__18 (.L_HI(net18));
 sg13g2_tiehi _4004__19 (.L_HI(net19));
 sg13g2_tiehi _4005__20 (.L_HI(net20));
 sg13g2_tiehi _4006__21 (.L_HI(net21));
 sg13g2_tiehi _4007__22 (.L_HI(net22));
 sg13g2_tiehi _4008__23 (.L_HI(net23));
 sg13g2_tiehi _4009__24 (.L_HI(net24));
 sg13g2_tiehi _4010__25 (.L_HI(net25));
 sg13g2_tiehi _4011__26 (.L_HI(net26));
 sg13g2_tiehi _4012__27 (.L_HI(net27));
 sg13g2_tiehi _4013__28 (.L_HI(net28));
 sg13g2_tiehi _4014__29 (.L_HI(net29));
 sg13g2_tiehi _4015__30 (.L_HI(net30));
 sg13g2_tiehi _4016__31 (.L_HI(net31));
 sg13g2_tiehi _4150__32 (.L_HI(net32));
 sg13g2_tiehi _4069__33 (.L_HI(net33));
 sg13g2_tiehi _4197__34 (.L_HI(net34));
 sg13g2_tiehi _4065__35 (.L_HI(net35));
 sg13g2_tiehi _4149__36 (.L_HI(net36));
 sg13g2_tiehi _4064__37 (.L_HI(net37));
 sg13g2_tiehi _4196__38 (.L_HI(net38));
 sg13g2_tiehi _4063__39 (.L_HI(net39));
 sg13g2_tiehi _4148__40 (.L_HI(net40));
 sg13g2_tiehi _4062__41 (.L_HI(net41));
 sg13g2_tiehi _4195__42 (.L_HI(net42));
 sg13g2_tiehi _4061__43 (.L_HI(net43));
 sg13g2_tiehi _4147__44 (.L_HI(net44));
 sg13g2_tiehi _4060__45 (.L_HI(net45));
 sg13g2_tiehi _4059__46 (.L_HI(net46));
 sg13g2_tiehi _4146__47 (.L_HI(net47));
 sg13g2_tiehi _4058__48 (.L_HI(net48));
 sg13g2_tiehi _4057__49 (.L_HI(net49));
 sg13g2_tiehi _4145__50 (.L_HI(net50));
 sg13g2_tiehi _4056__51 (.L_HI(net51));
 sg13g2_tiehi _4055__52 (.L_HI(net52));
 sg13g2_tiehi _4144__53 (.L_HI(net53));
 sg13g2_tiehi _4054__54 (.L_HI(net54));
 sg13g2_tiehi _4053__55 (.L_HI(net55));
 sg13g2_tiehi _4143__56 (.L_HI(net56));
 sg13g2_tiehi _4052__57 (.L_HI(net57));
 sg13g2_tiehi _4051__58 (.L_HI(net58));
 sg13g2_tiehi _4142__59 (.L_HI(net59));
 sg13g2_tiehi _4050__60 (.L_HI(net60));
 sg13g2_tiehi _4194__61 (.L_HI(net61));
 sg13g2_tiehi _4049__62 (.L_HI(net62));
 sg13g2_tiehi _4141__63 (.L_HI(net63));
 sg13g2_tiehi _4048__64 (.L_HI(net64));
 sg13g2_tiehi _4191__65 (.L_HI(net65));
 sg13g2_tiehi _4047__66 (.L_HI(net66));
 sg13g2_tiehi _4140__67 (.L_HI(net67));
 sg13g2_tiehi _4046__68 (.L_HI(net68));
 sg13g2_tiehi _4190__69 (.L_HI(net69));
 sg13g2_tiehi _4045__70 (.L_HI(net70));
 sg13g2_tiehi _4139__71 (.L_HI(net71));
 sg13g2_tiehi _4044__72 (.L_HI(net72));
 sg13g2_tiehi _4189__73 (.L_HI(net73));
 sg13g2_tiehi _4043__74 (.L_HI(net74));
 sg13g2_tiehi _4017__75 (.L_HI(net75));
 sg13g2_tiehi _4066__76 (.L_HI(net76));
 sg13g2_tiehi _4067__77 (.L_HI(net77));
 sg13g2_tiehi _4138__78 (.L_HI(net78));
 sg13g2_tiehi _4042__79 (.L_HI(net79));
 sg13g2_tiehi _4188__80 (.L_HI(net80));
 sg13g2_tiehi _4041__81 (.L_HI(net81));
 sg13g2_tiehi _4137__82 (.L_HI(net82));
 sg13g2_tiehi _4040__83 (.L_HI(net83));
 sg13g2_tiehi _4187__84 (.L_HI(net84));
 sg13g2_tiehi _4039__85 (.L_HI(net85));
 sg13g2_tiehi _4136__86 (.L_HI(net86));
 sg13g2_tiehi _4038__87 (.L_HI(net87));
 sg13g2_tiehi _4186__88 (.L_HI(net88));
 sg13g2_tiehi _4037__89 (.L_HI(net89));
 sg13g2_tiehi _4135__90 (.L_HI(net90));
 sg13g2_tiehi _4036__91 (.L_HI(net91));
 sg13g2_tiehi _4185__92 (.L_HI(net92));
 sg13g2_tiehi _4035__93 (.L_HI(net93));
 sg13g2_tiehi _4134__94 (.L_HI(net94));
 sg13g2_tiehi _4034__95 (.L_HI(net95));
 sg13g2_tiehi _4068__96 (.L_HI(net96));
 sg13g2_tiehi _4087__97 (.L_HI(net97));
 sg13g2_tiehi _4184__98 (.L_HI(net98));
 sg13g2_tiehi _4033__99 (.L_HI(net99));
 sg13g2_tiehi _4133__100 (.L_HI(net100));
 sg13g2_tiehi _4032__101 (.L_HI(net101));
 sg13g2_tiehi _4183__102 (.L_HI(net102));
 sg13g2_tiehi _4031__103 (.L_HI(net103));
 sg13g2_tiehi _4132__104 (.L_HI(net104));
 sg13g2_tiehi _4030__105 (.L_HI(net105));
 sg13g2_tiehi _4029__106 (.L_HI(net106));
 sg13g2_tiehi _4131__107 (.L_HI(net107));
 sg13g2_tiehi _4028__108 (.L_HI(net108));
 sg13g2_tiehi _4027__109 (.L_HI(net109));
 sg13g2_tiehi _4130__110 (.L_HI(net110));
 sg13g2_tiehi _4026__111 (.L_HI(net111));
 sg13g2_tiehi _4025__112 (.L_HI(net112));
 sg13g2_tiehi _4129__113 (.L_HI(net113));
 sg13g2_tiehi _4024__114 (.L_HI(net114));
 sg13g2_tiehi _4023__115 (.L_HI(net115));
 sg13g2_tiehi _4128__116 (.L_HI(net116));
 sg13g2_tiehi _4022__117 (.L_HI(net117));
 sg13g2_tiehi _4021__118 (.L_HI(net118));
 sg13g2_tiehi _4127__119 (.L_HI(net119));
 sg13g2_tiehi _4020__120 (.L_HI(net120));
 sg13g2_tiehi _4182__121 (.L_HI(net121));
 sg13g2_tiehi _4019__122 (.L_HI(net122));
 sg13g2_tiehi _4018__123 (.L_HI(net123));
 sg13g2_tiehi _4126__124 (.L_HI(net124));
 sg13g2_tiehi _4179__125 (.L_HI(net125));
 sg13g2_tiehi _4125__126 (.L_HI(net126));
 sg13g2_tiehi _4178__127 (.L_HI(net127));
 sg13g2_tiehi _4124__128 (.L_HI(net128));
 sg13g2_tiehi _4177__129 (.L_HI(net129));
 sg13g2_tiehi _4123__130 (.L_HI(net130));
 sg13g2_tiehi _4176__131 (.L_HI(net131));
 sg13g2_tiehi _4122__132 (.L_HI(net132));
 sg13g2_tiehi _4175__133 (.L_HI(net133));
 sg13g2_tiehi _4121__134 (.L_HI(net134));
 sg13g2_tiehi _4174__135 (.L_HI(net135));
 sg13g2_tiehi _4120__136 (.L_HI(net136));
 sg13g2_tiehi _4173__137 (.L_HI(net137));
 sg13g2_tiehi _4119__138 (.L_HI(net138));
 sg13g2_tiehi _4172__139 (.L_HI(net139));
 sg13g2_tiehi _4118__140 (.L_HI(net140));
 sg13g2_tiehi _4171__141 (.L_HI(net141));
 sg13g2_tiehi _4117__142 (.L_HI(net142));
 sg13g2_tiehi _4170__143 (.L_HI(net143));
 sg13g2_tiehi _4116__144 (.L_HI(net144));
 sg13g2_tiehi _4169__145 (.L_HI(net145));
 sg13g2_tiehi _4115__146 (.L_HI(net146));
 sg13g2_tiehi _4168__147 (.L_HI(net147));
 sg13g2_tiehi _4114__148 (.L_HI(net148));
 sg13g2_tiehi _4167__149 (.L_HI(net149));
 sg13g2_tiehi _4113__150 (.L_HI(net150));
 sg13g2_tiehi _4166__151 (.L_HI(net151));
 sg13g2_tiehi _4112__152 (.L_HI(net152));
 sg13g2_tiehi _4165__153 (.L_HI(net153));
 sg13g2_tiehi _4111__154 (.L_HI(net154));
 sg13g2_tiehi _4164__155 (.L_HI(net155));
 sg13g2_tiehi _4110__156 (.L_HI(net156));
 sg13g2_tiehi _4163__157 (.L_HI(net157));
 sg13g2_tiehi _4109__158 (.L_HI(net158));
 sg13g2_tiehi _4162__159 (.L_HI(net159));
 sg13g2_tiehi _4108__160 (.L_HI(net160));
 sg13g2_tiehi _4161__161 (.L_HI(net161));
 sg13g2_tiehi _4107__162 (.L_HI(net162));
 sg13g2_tiehi _4160__163 (.L_HI(net163));
 sg13g2_tiehi _4106__164 (.L_HI(net164));
 sg13g2_tiehi _4159__165 (.L_HI(net165));
 sg13g2_tiehi _4105__166 (.L_HI(net166));
 sg13g2_tiehi _4158__167 (.L_HI(net167));
 sg13g2_tiehi _4104__168 (.L_HI(net168));
 sg13g2_tiehi _4157__169 (.L_HI(net169));
 sg13g2_tiehi _4103__170 (.L_HI(net170));
 sg13g2_tiehi _4156__171 (.L_HI(net171));
 sg13g2_tiehi _4102__172 (.L_HI(net172));
 sg13g2_tiehi _4101__173 (.L_HI(net173));
 sg13g2_tiehi _4100__174 (.L_HI(net174));
 sg13g2_tiehi _4099__175 (.L_HI(net175));
 sg13g2_tiehi _4098__176 (.L_HI(net176));
 sg13g2_tiehi _4097__177 (.L_HI(net177));
 sg13g2_tiehi _4096__178 (.L_HI(net178));
 sg13g2_tiehi _4095__179 (.L_HI(net179));
 sg13g2_tiehi _4094__180 (.L_HI(net180));
 sg13g2_tiehi _4093__181 (.L_HI(net181));
 sg13g2_tiehi _4092__182 (.L_HI(net182));
 sg13g2_tiehi _4091__183 (.L_HI(net183));
 sg13g2_tiehi _4088__184 (.L_HI(net184));
 sg13g2_tiehi _4180__185 (.L_HI(net185));
 sg13g2_tiehi _4090__186 (.L_HI(net186));
 sg13g2_tiehi _4089__187 (.L_HI(net187));
 sg13g2_tiehi _4086__188 (.L_HI(net188));
 sg13g2_tiehi _4085__189 (.L_HI(net189));
 sg13g2_tiehi _4155__190 (.L_HI(net190));
 sg13g2_tiehi _4084__191 (.L_HI(net191));
 sg13g2_tiehi _4193__192 (.L_HI(net192));
 sg13g2_tiehi _4083__193 (.L_HI(net193));
 sg13g2_tiehi _4154__194 (.L_HI(net194));
 sg13g2_tiehi _4082__195 (.L_HI(net195));
 sg13g2_tiehi _4201__196 (.L_HI(net196));
 sg13g2_tiehi _4081__197 (.L_HI(net197));
 sg13g2_tiehi _4153__198 (.L_HI(net198));
 sg13g2_tiehi _4080__199 (.L_HI(net199));
 sg13g2_tiehi _4200__200 (.L_HI(net200));
 sg13g2_tiehi _4181__201 (.L_HI(net201));
 sg13g2_tiehi _4192__202 (.L_HI(net202));
 sg13g2_tiehi _4079__203 (.L_HI(net203));
 sg13g2_tiehi _4152__204 (.L_HI(net204));
 sg13g2_tiehi _4078__205 (.L_HI(net205));
 sg13g2_tiehi _4199__206 (.L_HI(net206));
 sg13g2_tiehi _4077__207 (.L_HI(net207));
 sg13g2_tiehi _4151__208 (.L_HI(net208));
 sg13g2_tiehi _4076__209 (.L_HI(net209));
 sg13g2_tiehi _4198__210 (.L_HI(net210));
 sg13g2_tiehi _4075__211 (.L_HI(net211));
 sg13g2_tiehi _4074__212 (.L_HI(net212));
 sg13g2_tiehi _4073__213 (.L_HI(net213));
 sg13g2_tiehi _4072__214 (.L_HI(net214));
 sg13g2_tiehi tt_um_algofoogle_fun_vga_clock_215 (.L_HI(net215));
 sg13g2_tiehi tt_um_algofoogle_fun_vga_clock_216 (.L_HI(net216));
 sg13g2_tiehi tt_um_algofoogle_fun_vga_clock_217 (.L_HI(net217));
 sg13g2_tiehi tt_um_algofoogle_fun_vga_clock_218 (.L_HI(net218));
 sg13g2_tiehi tt_um_algofoogle_fun_vga_clock_219 (.L_HI(net219));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_algofoogle_fun_vga_clock_8 (.L_LO(net8));
 sg13g2_tielo tt_um_algofoogle_fun_vga_clock_9 (.L_LO(net9));
 sg13g2_tielo tt_um_algofoogle_fun_vga_clock_10 (.L_LO(net10));
 sg13g2_tielo tt_um_algofoogle_fun_vga_clock_11 (.L_LO(net11));
 sg13g2_tielo tt_um_algofoogle_fun_vga_clock_12 (.L_LO(net12));
 sg13g2_tiehi _4071__13 (.L_HI(net13));
 sg13g2_buf_2 _4415_ (.A(hmax),
    .X(uio_out[0]));
 sg13g2_buf_2 _4416_ (.A(\vga_sync.o_vmax ),
    .X(uio_out[1]));
 sg13g2_buf_2 _4417_ (.A(hblank),
    .X(uio_out[2]));
 sg13g2_buf_2 _4418_ (.A(vblank),
    .X(uio_out[3]));
 sg13g2_buf_2 _4419_ (.A(\matt_venn_vga.activevideo ),
    .X(uio_out[4]));
 sg13g2_buf_2 fanout280 (.A(net282),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_1325_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_0985_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(net285),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_0829_),
    .X(net285));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_0821_));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_0598_),
    .X(net288));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(_0828_));
 sg13g2_buf_2 fanout290 (.A(net292),
    .X(net290));
 sg13g2_buf_1 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_1 fanout292 (.A(net293),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_0824_));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_1 fanout296 (.A(net297),
    .X(net296));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(_0824_));
 sg13g2_buf_2 fanout298 (.A(_0676_),
    .X(net298));
 sg13g2_buf_1 fanout299 (.A(_0676_),
    .X(net299));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(_0781_));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(net302));
 sg13g2_buf_2 fanout302 (.A(_0777_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_0505_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_1600_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_1546_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_0503_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_1556_),
    .X(net307));
 sg13g2_buf_4 fanout308 (.X(net308),
    .A(_1549_));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net311));
 sg13g2_buf_2 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(\matt_venn_vga.x_px[9] ),
    .X(net311));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(\matt_venn_vga.x_px[7] ));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(net314));
 sg13g2_buf_2 fanout314 (.A(net315),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(\matt_venn_vga.x_px[6] ),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(\h[5] ));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(net382));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(net536));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(\h[2] ));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(\h[1] ));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(\h[0] ));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(net524));
 sg13g2_buf_1 fanout324 (.A(\matt_venn_vga.y_px[9] ),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net326),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net544),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(\matt_venn_vga.y_px[7] ),
    .X(net328));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(\matt_venn_vga.y_px[6] ));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(net529));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(\matt_venn_vga.y_px[5] ));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(net512));
 sg13g2_buf_2 fanout333 (.A(\matt_venn_vga.y_px[4] ),
    .X(net333));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net535));
 sg13g2_buf_1 fanout335 (.A(\matt_venn_vga.y_px[3] ),
    .X(net335));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(net538));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(\matt_venn_vga.y_px[2] ));
 sg13g2_buf_2 fanout338 (.A(net339),
    .X(net338));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(\matt_venn_vga.y_px[1] ));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(net341));
 sg13g2_buf_2 fanout341 (.A(\matt_venn_vga.y_px[0] ),
    .X(net341));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(net343));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(dx));
 sg13g2_buf_2 fanout344 (.A(net553),
    .X(net344));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(net540));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(net554));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(net348));
 sg13g2_buf_2 fanout348 (.A(\py[0] ),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(net547),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(\px[7] ),
    .X(net350));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(\px[6] ));
 sg13g2_buf_2 fanout352 (.A(\px[5] ),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(\px[1] ),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(\px[0] ),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(\ydelta[7] ));
 sg13g2_buf_1 fanout356 (.A(\ydelta[7] ),
    .X(net356));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net359));
 sg13g2_buf_2 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(net360));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(_1398_));
 sg13g2_buf_2 fanout361 (.A(net4),
    .X(net361));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net364));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(net370));
 sg13g2_buf_2 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(net370));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(net369));
 sg13g2_buf_1 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(net370));
 sg13g2_buf_2 fanout370 (.A(rst_n),
    .X(net370));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[7]));
 sg13g2_tielo tt_um_algofoogle_fun_vga_clock_7 (.L_LO(net7));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_26_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_27_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_31_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_13_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_15_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_18_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_20_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\matt_venn_vga.col_index[1] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold2 (.A(\matt_venn_vga_shadow.col_index[0] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold3 (.A(\matt_venn_vga.col_index[0] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold4 (.A(\matt_venn_vga_shadow.col_index[1] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0071_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0076_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0077_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0967_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0075_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0189_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0074_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold12 (.A(_1206_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0192_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0078_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0846_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0073_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0198_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold18 (.A(\px[7] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold19 (.A(\clock_min_u[3] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0204_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold21 (.A(\matt_venn_clock.sec_counter[2] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold22 (.A(_1328_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0215_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold24 (.A(\matt_venn_clock.pulse_sec.count[4] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0188_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold26 (.A(\pxm[1] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold27 (.A(\matt_venn_clock.sec_counter[4] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold28 (.A(_1330_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold29 (.A(\matt_venn_clock.pulse_sec.count[3] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0187_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold31 (.A(\clock_sec_u[3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0211_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold33 (.A(\matt_venn_clock.sec_counter[3] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold34 (.A(_1329_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold35 (.A(\matt_venn_clock.pulse_hrs.comp[4] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold36 (.A(\matt_venn_clock.pulse_min.comp[4] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold37 (.A(\matt_venn_clock.pulse_min.count[4] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0178_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold39 (.A(\clock_sec_u[2] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0210_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold41 (.A(\matt_venn_clock.sec_counter[21] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold42 (.A(_1340_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0234_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold44 (.A(\px[6] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold45 (.A(\matt_venn_clock.sec_counter[5] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold46 (.A(\matt_venn_clock.pulse_hrs.count[4] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0168_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold48 (.A(\px[5] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0049_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0081_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold51 (.A(\matt_venn_clock.sec_counter[6] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0072_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0205_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold54 (.A(\matt_venn_clock.pulse_sec.comp[4] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0183_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold56 (.A(\matt_venn_clock.sec_counter[7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold57 (.A(\matt_venn_clock.pulse_min.count[3] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0177_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold59 (.A(\t[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0116_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold61 (.A(\matt_venn_clock.sec_counter[1] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1327_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold63 (.A(\matt_venn_clock.pulse_sec.comp[1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold64 (.A(_1160_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0052_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold66 (.A(_1215_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold67 (.A(\pym[11] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0054_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold69 (.A(_1336_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0231_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ydelta[3] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold72 (.A(\h[4] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold73 (.A(\vga_sync.vsync ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold74 (.A(\matt_venn_clock.sec_counter[19] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold75 (.A(_1338_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold76 (.A(\matt_venn_clock.sec_counter[22] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1341_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold78 (.A(\product_comp[10] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold79 (.A(_1016_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold80 (.A(\clock_hrs_d[1] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold81 (.A(_1208_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold82 (.A(\clock_sec_d[2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold83 (.A(_1262_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0207_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold85 (.A(\matt_venn_clock.pulse_min.count[2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pym[10] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0051_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0201_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold89 (.A(\matt_venn_clock.pulse_hrs.count[2] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold90 (.A(_1109_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0166_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold92 (.A(\clock_color_offset[1] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold93 (.A(_1195_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0038_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0208_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold96 (.A(\vga_sync.hsync ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0058_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0088_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold99 (.A(\clock_min_d[2] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold100 (.A(_1238_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0200_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0053_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold103 (.A(_1334_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold104 (.A(\matt_venn_vga.y_block_q[5] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold105 (.A(_1319_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold106 (.A(_1324_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0212_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold108 (.A(\matt_venn_clock.pulse_min.comp[1] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold109 (.A(_1125_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold110 (.A(\matt_venn_clock.sec_counter[24] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold111 (.A(_1342_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold112 (.A(\px[3] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold113 (.A(\matt_venn_clock.sec_counter[20] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold114 (.A(_1339_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold115 (.A(\clock_color_offset[2] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0191_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold117 (.A(\matt_venn_clock.pulse_sec.count[2] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0186_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0036_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold120 (.A(_1001_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold121 (.A(\clock_hrs_u[1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold122 (.A(\matt_venn_clock.pulse_hrs.comp[3] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0162_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold124 (.A(\matt_venn_clock.pulse_min.comp[2] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0033_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold126 (.A(_1013_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0034_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold128 (.A(_1010_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0035_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0123_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold131 (.A(\ydelta[6] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0087_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold133 (.A(\matt_venn_clock.pulse_sec.comp[0] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold134 (.A(\matt_venn_clock.pulse_hrs.count[3] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0167_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ydelta[5] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold137 (.A(\py[7] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold138 (.A(\clock_hrs_u[3] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold139 (.A(_1228_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold140 (.A(\matt_venn_clock.pulse_hrs.comp[2] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold141 (.A(_1092_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0161_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold143 (.A(\py[6] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold144 (.A(\matt_venn_clock.pulse_min.count[1] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0175_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold146 (.A(\t[2] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0115_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold148 (.A(\matt_venn_clock.pulse_min.comp[0] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold149 (.A(\matt_venn_clock.pulse_min.comp[3] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0172_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold151 (.A(\clock_hrs_u[2] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0196_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold153 (.A(\t[0] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0968_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0114_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold156 (.A(\matt_venn_vga_shadow.y_block_q[2] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold157 (.A(_1345_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold158 (.A(_1347_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0245_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold160 (.A(\matt_venn_clock.sec_counter[15] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold161 (.A(_1286_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold162 (.A(\matt_venn_clock.sec_counter[11] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold163 (.A(_1290_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold164 (.A(\matt_venn_clock.pulse_hrs.comp[1] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ydelta[4] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold166 (.A(\matt_venn_clock.sec_counter[17] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold167 (.A(_1335_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold168 (.A(\matt_venn_clock.pulse_sec.comp[2] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold169 (.A(\clock_sec_u[1] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0209_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold171 (.A(\ydelta[1] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold172 (.A(\matt_venn_clock.pulse_sec.count[1] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold173 (.A(_1182_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0185_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0037_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0121_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold177 (.A(\clock_min_u[2] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0203_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold179 (.A(\product_comp[0] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold180 (.A(\px[9] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold181 (.A(\px[4] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold182 (.A(\matt_venn_clock.pulse_hrs.comp[0] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold183 (.A(\matt_venn_clock.pulse_sec.comp[3] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold184 (.A(\clock_min_u[1] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold185 (.A(_1246_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold186 (.A(\matt_venn_clock.pulse_hrs.count[1] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0165_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold188 (.A(\matt_venn_clock.sec_counter[10] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1291_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ydelta[0] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0909_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0101_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold193 (.A(\py[5] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold194 (.A(\matt_venn_clock.sec_counter[14] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold195 (.A(_1287_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold196 (.A(\matt_venn_clock.sec_counter[9] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold197 (.A(_1292_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold198 (.A(\clock_hrs_d[0] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold199 (.A(\clock_min_d[1] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold200 (.A(_1236_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0199_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold202 (.A(\matt_venn_vga.y_px[4] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold203 (.A(\py[9] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold204 (.A(\product_comp[1] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold205 (.A(\matt_venn_clock.sec_counter[23] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold206 (.A(\matt_venn_clock.pulse_sec.count[0] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0025_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold208 (.A(\matt_venn_vga.digit_0.char[0] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold209 (.A(_1074_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold210 (.A(_1075_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold211 (.A(\px[2] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold212 (.A(\matt_venn_clock.sec_counter[16] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold213 (.A(\product_comp[2] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold214 (.A(\matt_venn_vga.y_px[9] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold215 (.A(\clock_sec_d[0] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold216 (.A(_1260_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0206_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold218 (.A(\py[8] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold219 (.A(\matt_venn_vga.y_px[5] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0139_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold221 (.A(\ydelta[2] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold222 (.A(\h[1] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold223 (.A(_1411_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold224 (.A(_1066_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold225 (.A(\matt_venn_vga.y_px[3] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold226 (.A(\h[3] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold227 (.A(\matt_venn_clock.sec_counter[8] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold228 (.A(\matt_venn_vga.y_px[2] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold229 (.A(\matt_venn_clock.pulse_min.count[0] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold230 (.A(\py[3] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold231 (.A(\py[2] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold232 (.A(\matt_venn_clock.pulse_hrs.count[0] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0047_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold234 (.A(\matt_venn_vga.y_px[8] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold235 (.A(\h[0] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold236 (.A(_1071_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold237 (.A(\px[8] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold238 (.A(\py[4] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold239 (.A(\product_comp[3] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold240 (.A(\matt_venn_vga.x_px[8] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold241 (.A(_1077_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0029_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold243 (.A(\product_comp[7] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold244 (.A(\py[1] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold245 (.A(\matt_venn_vga.y_px[7] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0056_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold247 (.A(\pxm[0] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold248 (.A(\matt_venn_vga.x_px[7] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold249 (.A(\matt_venn_clock.pulse_min.count[1] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold250 (.A(_1145_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold251 (.A(\matt_venn_clock.sec_counter[8] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold252 (.A(\clock_color_offset[1] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold253 (.A(\clock_color_offset[1] ),
    .X(net563));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(rst_n));
 sg13g2_antennanp ANTENNA_4 (.A(rst_n));
 sg13g2_antennanp ANTENNA_5 (.A(rst_n));
 sg13g2_antennanp ANTENNA_6 (.A(rst_n));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_4 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_decap_4 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_237 ();
 sg13g2_decap_8 FILLER_6_248 ();
 sg13g2_decap_4 FILLER_6_255 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_219 ();
 sg13g2_decap_4 FILLER_7_259 ();
 sg13g2_fill_2 FILLER_7_263 ();
 sg13g2_decap_4 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_decap_4 FILLER_7_283 ();
 sg13g2_fill_1 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_fill_2 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_163 ();
 sg13g2_decap_4 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_174 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_214 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_fill_1 FILLER_8_222 ();
 sg13g2_fill_1 FILLER_8_231 ();
 sg13g2_fill_2 FILLER_8_269 ();
 sg13g2_fill_2 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_310 ();
 sg13g2_decap_8 FILLER_8_317 ();
 sg13g2_decap_8 FILLER_8_324 ();
 sg13g2_decap_8 FILLER_8_331 ();
 sg13g2_decap_8 FILLER_8_338 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_221 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_fill_2 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_238 ();
 sg13g2_decap_4 FILLER_9_244 ();
 sg13g2_fill_1 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_4 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_4 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_204 ();
 sg13g2_fill_2 FILLER_10_251 ();
 sg13g2_fill_2 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_275 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_fill_2 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_208 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_fill_2 FILLER_11_237 ();
 sg13g2_decap_4 FILLER_11_244 ();
 sg13g2_fill_1 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_262 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_fill_2 FILLER_11_273 ();
 sg13g2_decap_4 FILLER_11_290 ();
 sg13g2_fill_2 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_fill_2 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_195 ();
 sg13g2_decap_8 FILLER_12_202 ();
 sg13g2_decap_8 FILLER_12_209 ();
 sg13g2_decap_4 FILLER_12_216 ();
 sg13g2_fill_2 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_311 ();
 sg13g2_decap_8 FILLER_12_318 ();
 sg13g2_decap_8 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_decap_8 FILLER_13_184 ();
 sg13g2_decap_8 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_220 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_decap_4 FILLER_13_263 ();
 sg13g2_decap_4 FILLER_13_272 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_decap_4 FILLER_13_282 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_decap_4 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_181 ();
 sg13g2_decap_8 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_fill_2 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_fill_2 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_4 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_4 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_decap_4 FILLER_15_194 ();
 sg13g2_decap_4 FILLER_15_229 ();
 sg13g2_fill_2 FILLER_15_233 ();
 sg13g2_decap_4 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_113 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_41 ();
 sg13g2_decap_8 FILLER_17_48 ();
 sg13g2_decap_8 FILLER_17_55 ();
 sg13g2_decap_8 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_69 ();
 sg13g2_decap_4 FILLER_17_76 ();
 sg13g2_fill_1 FILLER_17_118 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_decap_4 FILLER_17_213 ();
 sg13g2_fill_2 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_4 FILLER_17_241 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_292 ();
 sg13g2_decap_4 FILLER_17_299 ();
 sg13g2_fill_2 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_fill_2 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_2 FILLER_18_40 ();
 sg13g2_fill_2 FILLER_18_51 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_decap_8 FILLER_18_64 ();
 sg13g2_decap_8 FILLER_18_71 ();
 sg13g2_decap_8 FILLER_18_78 ();
 sg13g2_decap_4 FILLER_18_85 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_128 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_decap_8 FILLER_18_177 ();
 sg13g2_decap_4 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_198 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_4 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_4 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_18 ();
 sg13g2_fill_2 FILLER_19_45 ();
 sg13g2_fill_2 FILLER_19_61 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_73 ();
 sg13g2_decap_8 FILLER_19_80 ();
 sg13g2_decap_8 FILLER_19_87 ();
 sg13g2_decap_8 FILLER_19_94 ();
 sg13g2_decap_8 FILLER_19_101 ();
 sg13g2_decap_8 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_115 ();
 sg13g2_decap_8 FILLER_19_122 ();
 sg13g2_decap_8 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_decap_8 FILLER_19_150 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_decap_8 FILLER_19_164 ();
 sg13g2_decap_4 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_220 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_4 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_4 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_decap_4 FILLER_20_132 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_decap_4 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_decap_4 FILLER_20_177 ();
 sg13g2_fill_1 FILLER_20_207 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_357 ();
 sg13g2_fill_2 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_16 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_decap_8 FILLER_21_72 ();
 sg13g2_decap_8 FILLER_21_79 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_167 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_fill_2 FILLER_21_348 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_decap_4 FILLER_21_366 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_51 ();
 sg13g2_decap_8 FILLER_22_58 ();
 sg13g2_decap_8 FILLER_22_65 ();
 sg13g2_decap_8 FILLER_22_72 ();
 sg13g2_decap_4 FILLER_22_79 ();
 sg13g2_fill_2 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_147 ();
 sg13g2_fill_2 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_188 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_241 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_8 FILLER_22_293 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_fill_2 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_fill_1 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_66 ();
 sg13g2_decap_8 FILLER_23_73 ();
 sg13g2_decap_4 FILLER_23_80 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_fill_2 FILLER_23_197 ();
 sg13g2_decap_4 FILLER_23_222 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_250 ();
 sg13g2_decap_8 FILLER_23_257 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_288 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_4 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_351 ();
 sg13g2_decap_4 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_4 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_decap_4 FILLER_24_83 ();
 sg13g2_decap_4 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_111 ();
 sg13g2_decap_8 FILLER_24_118 ();
 sg13g2_decap_4 FILLER_24_125 ();
 sg13g2_fill_2 FILLER_24_129 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_decap_4 FILLER_24_153 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_decap_4 FILLER_24_173 ();
 sg13g2_decap_4 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_4 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_decap_4 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_decap_4 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_4 FILLER_24_329 ();
 sg13g2_decap_4 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_34 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_103 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_4 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_145 ();
 sg13g2_decap_8 FILLER_25_152 ();
 sg13g2_decap_4 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_fill_2 FILLER_25_243 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_decap_4 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_decap_4 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_64 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_118 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_decap_4 FILLER_26_132 ();
 sg13g2_decap_4 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_decap_4 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_287 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_decap_4 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_16 ();
 sg13g2_fill_1 FILLER_27_18 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_54 ();
 sg13g2_fill_1 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_66 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_decap_8 FILLER_27_79 ();
 sg13g2_decap_4 FILLER_27_86 ();
 sg13g2_decap_4 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_decap_8 FILLER_27_162 ();
 sg13g2_decap_4 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_2 FILLER_27_178 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_256 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_4 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_fill_2 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_fill_2 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_4 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_fill_2 FILLER_27_379 ();
 sg13g2_fill_1 FILLER_27_381 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_58 ();
 sg13g2_decap_4 FILLER_28_65 ();
 sg13g2_fill_1 FILLER_28_69 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_decap_4 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_187 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_65 ();
 sg13g2_decap_8 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_decap_8 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_103 ();
 sg13g2_decap_8 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_decap_4 FILLER_29_129 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_decap_4 FILLER_29_192 ();
 sg13g2_decap_4 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_fill_2 FILLER_29_393 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_109 ();
 sg13g2_decap_4 FILLER_30_119 ();
 sg13g2_fill_2 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_139 ();
 sg13g2_decap_4 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_decap_4 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_204 ();
 sg13g2_fill_1 FILLER_30_206 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_4 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_decap_4 FILLER_30_380 ();
 sg13g2_fill_1 FILLER_31_40 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_decap_4 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_241 ();
 sg13g2_decap_8 FILLER_31_250 ();
 sg13g2_decap_4 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_decap_4 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_decap_8 FILLER_32_44 ();
 sg13g2_decap_4 FILLER_32_51 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_decap_8 FILLER_32_97 ();
 sg13g2_decap_8 FILLER_32_104 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_150 ();
 sg13g2_decap_4 FILLER_32_157 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_208 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_289 ();
 sg13g2_decap_8 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_385 ();
 sg13g2_decap_4 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_23 ();
 sg13g2_fill_2 FILLER_33_29 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_39 ();
 sg13g2_decap_8 FILLER_33_54 ();
 sg13g2_decap_4 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_79 ();
 sg13g2_fill_2 FILLER_33_106 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_4 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_decap_8 FILLER_33_248 ();
 sg13g2_decap_4 FILLER_33_255 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_362 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_13 ();
 sg13g2_decap_4 FILLER_34_20 ();
 sg13g2_fill_2 FILLER_34_24 ();
 sg13g2_fill_2 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_89 ();
 sg13g2_fill_2 FILLER_34_95 ();
 sg13g2_decap_8 FILLER_34_127 ();
 sg13g2_decap_8 FILLER_34_134 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_decap_4 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_decap_4 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_decap_4 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_decap_4 FILLER_35_113 ();
 sg13g2_fill_2 FILLER_35_117 ();
 sg13g2_decap_8 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_decap_4 FILLER_35_195 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_decap_4 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_fill_2 FILLER_35_350 ();
 sg13g2_decap_4 FILLER_35_393 ();
 sg13g2_decap_4 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_74 ();
 sg13g2_decap_4 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_211 ();
 sg13g2_decap_4 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_307 ();
 sg13g2_decap_8 FILLER_36_314 ();
 sg13g2_decap_8 FILLER_36_321 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_fill_2 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_4 FILLER_37_39 ();
 sg13g2_fill_1 FILLER_37_43 ();
 sg13g2_decap_8 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_74 ();
 sg13g2_decap_4 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_85 ();
 sg13g2_decap_8 FILLER_37_90 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_decap_8 FILLER_37_104 ();
 sg13g2_fill_2 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_121 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_decap_8 FILLER_37_134 ();
 sg13g2_fill_2 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_143 ();
 sg13g2_decap_8 FILLER_37_153 ();
 sg13g2_fill_2 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_162 ();
 sg13g2_decap_8 FILLER_37_176 ();
 sg13g2_decap_8 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_219 ();
 sg13g2_decap_8 FILLER_37_226 ();
 sg13g2_decap_8 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_decap_4 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_330 ();
 sg13g2_decap_4 FILLER_37_362 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_fill_2 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_5 ();
 sg13g2_decap_4 FILLER_38_12 ();
 sg13g2_fill_2 FILLER_38_16 ();
 sg13g2_fill_1 FILLER_38_23 ();
 sg13g2_decap_4 FILLER_38_38 ();
 sg13g2_decap_4 FILLER_38_58 ();
 sg13g2_fill_2 FILLER_38_62 ();
 sg13g2_decap_4 FILLER_38_90 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_decap_8 FILLER_38_111 ();
 sg13g2_decap_4 FILLER_38_118 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_decap_4 FILLER_38_127 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_decap_8 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_decap_8 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_158 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_235 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_decap_4 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_19 ();
 sg13g2_decap_4 FILLER_39_37 ();
 sg13g2_decap_8 FILLER_39_62 ();
 sg13g2_fill_2 FILLER_39_69 ();
 sg13g2_fill_1 FILLER_39_71 ();
 sg13g2_decap_4 FILLER_39_80 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_fill_2 FILLER_39_111 ();
 sg13g2_fill_1 FILLER_39_113 ();
 sg13g2_decap_4 FILLER_39_140 ();
 sg13g2_fill_2 FILLER_39_160 ();
 sg13g2_fill_2 FILLER_39_167 ();
 sg13g2_fill_1 FILLER_39_169 ();
 sg13g2_fill_2 FILLER_39_182 ();
 sg13g2_fill_1 FILLER_39_198 ();
 sg13g2_decap_4 FILLER_39_204 ();
 sg13g2_fill_2 FILLER_39_229 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_fill_1 FILLER_39_242 ();
 sg13g2_fill_2 FILLER_39_255 ();
 sg13g2_fill_2 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_281 ();
 sg13g2_fill_1 FILLER_39_283 ();
 sg13g2_fill_2 FILLER_39_292 ();
 sg13g2_decap_8 FILLER_39_328 ();
 sg13g2_decap_8 FILLER_39_335 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_decap_4 FILLER_39_360 ();
 sg13g2_fill_1 FILLER_39_364 ();
 sg13g2_fill_2 FILLER_39_371 ();
 sg13g2_fill_2 FILLER_39_389 ();
 sg13g2_fill_1 FILLER_39_391 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_fill_1 FILLER_40_35 ();
 sg13g2_fill_2 FILLER_40_139 ();
 sg13g2_fill_1 FILLER_40_189 ();
 sg13g2_fill_2 FILLER_40_197 ();
 sg13g2_fill_1 FILLER_40_199 ();
 sg13g2_decap_8 FILLER_40_209 ();
 sg13g2_fill_2 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_218 ();
 sg13g2_decap_8 FILLER_40_230 ();
 sg13g2_decap_8 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_fill_1 FILLER_40_282 ();
 sg13g2_decap_8 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_decap_8 FILLER_40_309 ();
 sg13g2_decap_4 FILLER_40_316 ();
 sg13g2_fill_1 FILLER_40_320 ();
 sg13g2_decap_4 FILLER_40_346 ();
 sg13g2_fill_2 FILLER_40_350 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_fill_2 FILLER_40_375 ();
 sg13g2_fill_2 FILLER_40_385 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_59 ();
 sg13g2_decap_8 FILLER_41_66 ();
 sg13g2_decap_8 FILLER_41_73 ();
 sg13g2_decap_8 FILLER_41_80 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_fill_1 FILLER_41_89 ();
 sg13g2_decap_4 FILLER_41_100 ();
 sg13g2_fill_2 FILLER_41_114 ();
 sg13g2_fill_1 FILLER_41_116 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_fill_1 FILLER_41_151 ();
 sg13g2_fill_1 FILLER_41_160 ();
 sg13g2_decap_4 FILLER_41_179 ();
 sg13g2_fill_2 FILLER_41_183 ();
 sg13g2_decap_4 FILLER_41_193 ();
 sg13g2_fill_1 FILLER_41_205 ();
 sg13g2_decap_8 FILLER_41_219 ();
 sg13g2_fill_2 FILLER_41_226 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_fill_2 FILLER_41_237 ();
 sg13g2_decap_8 FILLER_41_244 ();
 sg13g2_decap_4 FILLER_41_251 ();
 sg13g2_fill_2 FILLER_41_255 ();
 sg13g2_decap_8 FILLER_41_261 ();
 sg13g2_decap_8 FILLER_41_268 ();
 sg13g2_fill_2 FILLER_41_275 ();
 sg13g2_fill_1 FILLER_41_277 ();
 sg13g2_fill_2 FILLER_41_291 ();
 sg13g2_fill_1 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_299 ();
 sg13g2_decap_8 FILLER_41_319 ();
 sg13g2_decap_8 FILLER_41_326 ();
 sg13g2_decap_4 FILLER_41_333 ();
 sg13g2_fill_2 FILLER_41_337 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_4 FILLER_41_357 ();
 sg13g2_fill_2 FILLER_41_361 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_381 ();
 sg13g2_fill_2 FILLER_42_55 ();
 sg13g2_fill_1 FILLER_42_57 ();
 sg13g2_decap_4 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_75 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_4 FILLER_42_119 ();
 sg13g2_fill_1 FILLER_42_123 ();
 sg13g2_decap_4 FILLER_42_136 ();
 sg13g2_fill_1 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_163 ();
 sg13g2_decap_8 FILLER_42_170 ();
 sg13g2_decap_8 FILLER_42_177 ();
 sg13g2_decap_8 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_191 ();
 sg13g2_fill_2 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_205 ();
 sg13g2_fill_1 FILLER_42_207 ();
 sg13g2_fill_2 FILLER_42_213 ();
 sg13g2_decap_8 FILLER_42_220 ();
 sg13g2_decap_8 FILLER_42_257 ();
 sg13g2_decap_4 FILLER_42_264 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_decap_4 FILLER_42_284 ();
 sg13g2_fill_2 FILLER_42_288 ();
 sg13g2_decap_8 FILLER_42_316 ();
 sg13g2_decap_4 FILLER_42_323 ();
 sg13g2_fill_2 FILLER_42_327 ();
 sg13g2_fill_2 FILLER_42_352 ();
 sg13g2_fill_1 FILLER_42_354 ();
 sg13g2_fill_1 FILLER_42_365 ();
 sg13g2_decap_8 FILLER_42_381 ();
 sg13g2_decap_8 FILLER_42_388 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_16 ();
 sg13g2_fill_2 FILLER_43_93 ();
 sg13g2_fill_1 FILLER_43_95 ();
 sg13g2_decap_8 FILLER_43_109 ();
 sg13g2_decap_8 FILLER_43_116 ();
 sg13g2_decap_8 FILLER_43_123 ();
 sg13g2_decap_8 FILLER_43_130 ();
 sg13g2_decap_8 FILLER_43_137 ();
 sg13g2_decap_8 FILLER_43_144 ();
 sg13g2_decap_8 FILLER_43_151 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_fill_2 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_215 ();
 sg13g2_fill_2 FILLER_43_241 ();
 sg13g2_decap_8 FILLER_43_254 ();
 sg13g2_decap_8 FILLER_43_261 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_fill_2 FILLER_43_294 ();
 sg13g2_fill_1 FILLER_43_316 ();
 sg13g2_decap_4 FILLER_43_333 ();
 sg13g2_fill_1 FILLER_43_337 ();
 sg13g2_fill_2 FILLER_43_347 ();
 sg13g2_fill_2 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_365 ();
 sg13g2_decap_8 FILLER_43_372 ();
 sg13g2_fill_2 FILLER_43_379 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_4 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_4 FILLER_44_70 ();
 sg13g2_fill_1 FILLER_44_74 ();
 sg13g2_decap_4 FILLER_44_83 ();
 sg13g2_fill_1 FILLER_44_87 ();
 sg13g2_decap_8 FILLER_44_113 ();
 sg13g2_decap_8 FILLER_44_120 ();
 sg13g2_decap_8 FILLER_44_127 ();
 sg13g2_fill_2 FILLER_44_134 ();
 sg13g2_fill_1 FILLER_44_136 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_fill_1 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_fill_2 FILLER_44_240 ();
 sg13g2_fill_2 FILLER_44_250 ();
 sg13g2_fill_1 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_decap_4 FILLER_44_332 ();
 sg13g2_fill_2 FILLER_44_336 ();
 sg13g2_fill_2 FILLER_44_346 ();
 sg13g2_fill_2 FILLER_44_356 ();
 sg13g2_fill_1 FILLER_44_358 ();
 sg13g2_fill_2 FILLER_44_372 ();
 sg13g2_fill_2 FILLER_44_395 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_15 ();
 sg13g2_decap_8 FILLER_45_61 ();
 sg13g2_decap_8 FILLER_45_68 ();
 sg13g2_decap_8 FILLER_45_75 ();
 sg13g2_decap_4 FILLER_45_82 ();
 sg13g2_fill_2 FILLER_45_104 ();
 sg13g2_fill_1 FILLER_45_195 ();
 sg13g2_fill_1 FILLER_45_205 ();
 sg13g2_decap_4 FILLER_45_211 ();
 sg13g2_decap_8 FILLER_45_219 ();
 sg13g2_decap_8 FILLER_45_226 ();
 sg13g2_decap_8 FILLER_45_233 ();
 sg13g2_fill_2 FILLER_45_240 ();
 sg13g2_decap_4 FILLER_45_258 ();
 sg13g2_fill_1 FILLER_45_262 ();
 sg13g2_decap_8 FILLER_45_276 ();
 sg13g2_decap_4 FILLER_45_283 ();
 sg13g2_fill_2 FILLER_45_287 ();
 sg13g2_fill_2 FILLER_45_314 ();
 sg13g2_decap_8 FILLER_45_324 ();
 sg13g2_decap_8 FILLER_45_331 ();
 sg13g2_decap_8 FILLER_45_338 ();
 sg13g2_decap_8 FILLER_45_345 ();
 sg13g2_decap_8 FILLER_45_352 ();
 sg13g2_decap_8 FILLER_45_359 ();
 sg13g2_decap_8 FILLER_45_366 ();
 sg13g2_decap_8 FILLER_45_373 ();
 sg13g2_decap_8 FILLER_45_380 ();
 sg13g2_fill_2 FILLER_45_387 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_39 ();
 sg13g2_decap_8 FILLER_46_53 ();
 sg13g2_decap_8 FILLER_46_60 ();
 sg13g2_fill_1 FILLER_46_67 ();
 sg13g2_fill_1 FILLER_46_89 ();
 sg13g2_fill_2 FILLER_46_94 ();
 sg13g2_fill_1 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_102 ();
 sg13g2_fill_2 FILLER_46_110 ();
 sg13g2_fill_1 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_139 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_decap_8 FILLER_46_177 ();
 sg13g2_decap_8 FILLER_46_184 ();
 sg13g2_decap_4 FILLER_46_191 ();
 sg13g2_fill_2 FILLER_46_195 ();
 sg13g2_fill_1 FILLER_46_254 ();
 sg13g2_fill_1 FILLER_46_286 ();
 sg13g2_fill_2 FILLER_46_296 ();
 sg13g2_decap_8 FILLER_46_304 ();
 sg13g2_decap_8 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_318 ();
 sg13g2_fill_2 FILLER_46_325 ();
 sg13g2_fill_1 FILLER_46_327 ();
 sg13g2_fill_2 FILLER_46_336 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_decap_4 FILLER_46_376 ();
 sg13g2_fill_2 FILLER_46_380 ();
 sg13g2_decap_8 FILLER_47_110 ();
 sg13g2_decap_8 FILLER_47_117 ();
 sg13g2_fill_2 FILLER_47_124 ();
 sg13g2_decap_4 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_143 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_164 ();
 sg13g2_decap_8 FILLER_47_169 ();
 sg13g2_decap_8 FILLER_47_176 ();
 sg13g2_decap_4 FILLER_47_183 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_decap_8 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_265 ();
 sg13g2_decap_8 FILLER_47_270 ();
 sg13g2_fill_2 FILLER_47_277 ();
 sg13g2_fill_1 FILLER_47_279 ();
 sg13g2_decap_8 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_291 ();
 sg13g2_decap_8 FILLER_47_296 ();
 sg13g2_decap_4 FILLER_47_303 ();
 sg13g2_fill_2 FILLER_47_307 ();
 sg13g2_decap_8 FILLER_47_333 ();
 sg13g2_decap_4 FILLER_47_340 ();
 sg13g2_fill_1 FILLER_47_344 ();
 sg13g2_fill_2 FILLER_47_349 ();
 sg13g2_fill_1 FILLER_47_351 ();
 sg13g2_fill_2 FILLER_47_356 ();
 sg13g2_fill_1 FILLER_47_358 ();
 sg13g2_decap_4 FILLER_47_378 ();
 sg13g2_fill_2 FILLER_47_382 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_15 ();
 sg13g2_decap_8 FILLER_48_22 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_fill_1 FILLER_48_39 ();
 sg13g2_decap_8 FILLER_48_52 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_fill_1 FILLER_48_70 ();
 sg13g2_fill_1 FILLER_48_78 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_4 FILLER_48_133 ();
 sg13g2_fill_1 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_167 ();
 sg13g2_fill_1 FILLER_48_174 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_fill_1 FILLER_48_245 ();
 sg13g2_fill_2 FILLER_48_251 ();
 sg13g2_fill_1 FILLER_48_253 ();
 sg13g2_fill_1 FILLER_48_271 ();
 sg13g2_fill_2 FILLER_48_280 ();
 sg13g2_fill_2 FILLER_48_299 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_fill_2 FILLER_48_350 ();
 sg13g2_fill_1 FILLER_48_352 ();
 sg13g2_fill_1 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_fill_2 FILLER_48_392 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_decap_4 FILLER_48_403 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_1 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_fill_1 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_143 ();
 sg13g2_decap_4 FILLER_49_150 ();
 sg13g2_fill_1 FILLER_49_154 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_fill_1 FILLER_49_197 ();
 sg13g2_decap_8 FILLER_49_208 ();
 sg13g2_decap_8 FILLER_49_215 ();
 sg13g2_decap_8 FILLER_49_222 ();
 sg13g2_decap_8 FILLER_49_229 ();
 sg13g2_decap_4 FILLER_49_236 ();
 sg13g2_fill_1 FILLER_49_240 ();
 sg13g2_fill_2 FILLER_49_246 ();
 sg13g2_fill_1 FILLER_49_248 ();
 sg13g2_fill_1 FILLER_49_265 ();
 sg13g2_fill_1 FILLER_49_292 ();
 sg13g2_decap_8 FILLER_49_344 ();
 sg13g2_decap_4 FILLER_49_351 ();
 sg13g2_fill_1 FILLER_49_360 ();
 sg13g2_decap_8 FILLER_49_383 ();
 sg13g2_decap_4 FILLER_49_390 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_35 ();
 sg13g2_fill_1 FILLER_50_37 ();
 sg13g2_fill_1 FILLER_50_47 ();
 sg13g2_decap_4 FILLER_50_74 ();
 sg13g2_fill_1 FILLER_50_78 ();
 sg13g2_fill_2 FILLER_50_108 ();
 sg13g2_fill_1 FILLER_50_140 ();
 sg13g2_decap_4 FILLER_50_147 ();
 sg13g2_fill_2 FILLER_50_151 ();
 sg13g2_decap_8 FILLER_50_169 ();
 sg13g2_decap_8 FILLER_50_176 ();
 sg13g2_decap_4 FILLER_50_183 ();
 sg13g2_decap_8 FILLER_50_192 ();
 sg13g2_decap_8 FILLER_50_199 ();
 sg13g2_decap_4 FILLER_50_206 ();
 sg13g2_fill_1 FILLER_50_210 ();
 sg13g2_decap_4 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_237 ();
 sg13g2_decap_4 FILLER_50_256 ();
 sg13g2_fill_1 FILLER_50_265 ();
 sg13g2_fill_2 FILLER_50_274 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_decap_8 FILLER_50_341 ();
 sg13g2_decap_4 FILLER_50_348 ();
 sg13g2_fill_1 FILLER_50_352 ();
 sg13g2_decap_8 FILLER_50_357 ();
 sg13g2_decap_4 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_377 ();
 sg13g2_decap_4 FILLER_50_384 ();
 sg13g2_fill_2 FILLER_50_388 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_18 ();
 sg13g2_fill_2 FILLER_51_27 ();
 sg13g2_decap_4 FILLER_51_55 ();
 sg13g2_decap_4 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_74 ();
 sg13g2_decap_4 FILLER_51_81 ();
 sg13g2_fill_1 FILLER_51_85 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_107 ();
 sg13g2_decap_4 FILLER_51_114 ();
 sg13g2_fill_2 FILLER_51_125 ();
 sg13g2_fill_2 FILLER_51_131 ();
 sg13g2_fill_2 FILLER_51_179 ();
 sg13g2_fill_1 FILLER_51_198 ();
 sg13g2_decap_8 FILLER_51_204 ();
 sg13g2_decap_8 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_218 ();
 sg13g2_decap_8 FILLER_51_225 ();
 sg13g2_decap_8 FILLER_51_232 ();
 sg13g2_decap_8 FILLER_51_239 ();
 sg13g2_decap_8 FILLER_51_246 ();
 sg13g2_decap_8 FILLER_51_253 ();
 sg13g2_decap_8 FILLER_51_260 ();
 sg13g2_decap_8 FILLER_51_267 ();
 sg13g2_fill_1 FILLER_51_274 ();
 sg13g2_decap_8 FILLER_51_279 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_decap_8 FILLER_51_291 ();
 sg13g2_fill_1 FILLER_51_298 ();
 sg13g2_decap_8 FILLER_51_304 ();
 sg13g2_decap_8 FILLER_51_311 ();
 sg13g2_decap_4 FILLER_51_318 ();
 sg13g2_decap_8 FILLER_51_327 ();
 sg13g2_fill_2 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_decap_4 FILLER_51_385 ();
 sg13g2_fill_2 FILLER_51_394 ();
 sg13g2_fill_1 FILLER_51_396 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_81 ();
 sg13g2_decap_8 FILLER_52_88 ();
 sg13g2_decap_8 FILLER_52_95 ();
 sg13g2_decap_8 FILLER_52_102 ();
 sg13g2_decap_4 FILLER_52_109 ();
 sg13g2_decap_8 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_235 ();
 sg13g2_fill_1 FILLER_52_237 ();
 sg13g2_decap_8 FILLER_52_251 ();
 sg13g2_decap_8 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_265 ();
 sg13g2_decap_8 FILLER_52_271 ();
 sg13g2_decap_4 FILLER_52_278 ();
 sg13g2_fill_2 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_326 ();
 sg13g2_fill_2 FILLER_52_353 ();
 sg13g2_fill_1 FILLER_52_355 ();
 sg13g2_fill_2 FILLER_52_365 ();
 sg13g2_fill_2 FILLER_52_387 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_fill_2 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_37 ();
 sg13g2_decap_4 FILLER_53_50 ();
 sg13g2_fill_1 FILLER_53_54 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_89 ();
 sg13g2_decap_8 FILLER_53_96 ();
 sg13g2_fill_1 FILLER_53_103 ();
 sg13g2_fill_2 FILLER_53_135 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_fill_1 FILLER_53_150 ();
 sg13g2_fill_1 FILLER_53_168 ();
 sg13g2_fill_1 FILLER_53_177 ();
 sg13g2_decap_8 FILLER_53_202 ();
 sg13g2_decap_4 FILLER_53_209 ();
 sg13g2_fill_1 FILLER_53_213 ();
 sg13g2_fill_2 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_224 ();
 sg13g2_decap_4 FILLER_53_279 ();
 sg13g2_decap_4 FILLER_53_288 ();
 sg13g2_fill_1 FILLER_53_328 ();
 sg13g2_fill_2 FILLER_53_333 ();
 sg13g2_fill_1 FILLER_53_335 ();
 sg13g2_decap_4 FILLER_53_383 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_4 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_25 ();
 sg13g2_fill_2 FILLER_54_57 ();
 sg13g2_fill_1 FILLER_54_59 ();
 sg13g2_fill_2 FILLER_54_65 ();
 sg13g2_fill_1 FILLER_54_67 ();
 sg13g2_decap_8 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_fill_1 FILLER_54_91 ();
 sg13g2_fill_1 FILLER_54_118 ();
 sg13g2_decap_8 FILLER_54_127 ();
 sg13g2_decap_8 FILLER_54_134 ();
 sg13g2_fill_1 FILLER_54_141 ();
 sg13g2_fill_2 FILLER_54_148 ();
 sg13g2_fill_1 FILLER_54_150 ();
 sg13g2_fill_1 FILLER_54_156 ();
 sg13g2_decap_4 FILLER_54_176 ();
 sg13g2_decap_8 FILLER_54_195 ();
 sg13g2_decap_4 FILLER_54_202 ();
 sg13g2_decap_8 FILLER_54_209 ();
 sg13g2_decap_4 FILLER_54_216 ();
 sg13g2_fill_2 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_226 ();
 sg13g2_fill_2 FILLER_54_233 ();
 sg13g2_fill_1 FILLER_54_235 ();
 sg13g2_fill_2 FILLER_54_257 ();
 sg13g2_fill_2 FILLER_54_337 ();
 sg13g2_fill_2 FILLER_54_361 ();
 sg13g2_fill_2 FILLER_54_376 ();
 sg13g2_decap_4 FILLER_54_383 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_11 ();
 sg13g2_decap_8 FILLER_55_69 ();
 sg13g2_fill_1 FILLER_55_76 ();
 sg13g2_decap_8 FILLER_55_80 ();
 sg13g2_decap_8 FILLER_55_87 ();
 sg13g2_decap_8 FILLER_55_94 ();
 sg13g2_decap_4 FILLER_55_101 ();
 sg13g2_fill_1 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_115 ();
 sg13g2_decap_8 FILLER_55_122 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_fill_1 FILLER_55_131 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_186 ();
 sg13g2_decap_8 FILLER_55_193 ();
 sg13g2_decap_8 FILLER_55_235 ();
 sg13g2_decap_8 FILLER_55_242 ();
 sg13g2_decap_8 FILLER_55_249 ();
 sg13g2_fill_2 FILLER_55_256 ();
 sg13g2_fill_1 FILLER_55_258 ();
 sg13g2_decap_8 FILLER_55_276 ();
 sg13g2_fill_2 FILLER_55_283 ();
 sg13g2_fill_1 FILLER_55_285 ();
 sg13g2_decap_8 FILLER_55_290 ();
 sg13g2_decap_8 FILLER_55_297 ();
 sg13g2_fill_2 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_306 ();
 sg13g2_decap_4 FILLER_55_311 ();
 sg13g2_fill_2 FILLER_55_315 ();
 sg13g2_decap_8 FILLER_55_326 ();
 sg13g2_decap_4 FILLER_55_333 ();
 sg13g2_fill_1 FILLER_55_345 ();
 sg13g2_decap_8 FILLER_55_362 ();
 sg13g2_decap_8 FILLER_55_369 ();
 sg13g2_decap_8 FILLER_55_376 ();
 sg13g2_fill_1 FILLER_55_383 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_11 ();
 sg13g2_fill_2 FILLER_56_41 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_fill_1 FILLER_56_62 ();
 sg13g2_decap_8 FILLER_56_80 ();
 sg13g2_decap_8 FILLER_56_93 ();
 sg13g2_fill_1 FILLER_56_100 ();
 sg13g2_fill_1 FILLER_56_106 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_decap_4 FILLER_56_133 ();
 sg13g2_fill_1 FILLER_56_137 ();
 sg13g2_decap_8 FILLER_56_164 ();
 sg13g2_fill_1 FILLER_56_180 ();
 sg13g2_decap_8 FILLER_56_192 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_201 ();
 sg13g2_decap_8 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_242 ();
 sg13g2_decap_8 FILLER_56_249 ();
 sg13g2_decap_8 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_263 ();
 sg13g2_fill_1 FILLER_56_265 ();
 sg13g2_decap_8 FILLER_56_271 ();
 sg13g2_decap_4 FILLER_56_278 ();
 sg13g2_fill_2 FILLER_56_282 ();
 sg13g2_fill_2 FILLER_56_313 ();
 sg13g2_fill_2 FILLER_56_341 ();
 sg13g2_decap_4 FILLER_56_360 ();
 sg13g2_fill_1 FILLER_56_364 ();
 sg13g2_decap_4 FILLER_56_391 ();
 sg13g2_decap_4 FILLER_56_405 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_22 ();
 sg13g2_fill_1 FILLER_57_24 ();
 sg13g2_fill_1 FILLER_57_104 ();
 sg13g2_fill_1 FILLER_57_111 ();
 sg13g2_fill_2 FILLER_57_120 ();
 sg13g2_fill_2 FILLER_57_136 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_159 ();
 sg13g2_fill_2 FILLER_57_177 ();
 sg13g2_fill_1 FILLER_57_206 ();
 sg13g2_fill_1 FILLER_57_245 ();
 sg13g2_fill_2 FILLER_57_254 ();
 sg13g2_fill_1 FILLER_57_256 ();
 sg13g2_decap_4 FILLER_57_277 ();
 sg13g2_fill_2 FILLER_57_307 ();
 sg13g2_fill_1 FILLER_57_309 ();
 sg13g2_decap_4 FILLER_57_322 ();
 sg13g2_fill_2 FILLER_57_330 ();
 sg13g2_fill_1 FILLER_57_332 ();
 sg13g2_decap_8 FILLER_57_356 ();
 sg13g2_fill_2 FILLER_57_373 ();
 sg13g2_fill_1 FILLER_57_396 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_fill_1 FILLER_58_35 ();
 sg13g2_fill_2 FILLER_58_41 ();
 sg13g2_fill_1 FILLER_58_43 ();
 sg13g2_decap_4 FILLER_58_74 ();
 sg13g2_decap_8 FILLER_58_92 ();
 sg13g2_decap_4 FILLER_58_99 ();
 sg13g2_fill_2 FILLER_58_103 ();
 sg13g2_fill_1 FILLER_58_108 ();
 sg13g2_fill_2 FILLER_58_129 ();
 sg13g2_fill_2 FILLER_58_148 ();
 sg13g2_fill_2 FILLER_58_154 ();
 sg13g2_decap_4 FILLER_58_167 ();
 sg13g2_fill_2 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_204 ();
 sg13g2_fill_1 FILLER_58_206 ();
 sg13g2_decap_4 FILLER_58_212 ();
 sg13g2_decap_4 FILLER_58_231 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_fill_2 FILLER_58_283 ();
 sg13g2_fill_1 FILLER_58_285 ();
 sg13g2_decap_4 FILLER_58_316 ();
 sg13g2_fill_2 FILLER_58_320 ();
 sg13g2_decap_8 FILLER_58_327 ();
 sg13g2_decap_4 FILLER_58_334 ();
 sg13g2_decap_4 FILLER_58_351 ();
 sg13g2_fill_2 FILLER_58_359 ();
 sg13g2_fill_2 FILLER_58_366 ();
 sg13g2_decap_4 FILLER_58_386 ();
 sg13g2_fill_1 FILLER_58_390 ();
 sg13g2_fill_1 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_fill_2 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_32 ();
 sg13g2_fill_2 FILLER_59_56 ();
 sg13g2_fill_1 FILLER_59_83 ();
 sg13g2_decap_8 FILLER_59_88 ();
 sg13g2_decap_4 FILLER_59_95 ();
 sg13g2_fill_1 FILLER_59_99 ();
 sg13g2_fill_2 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_fill_2 FILLER_59_119 ();
 sg13g2_fill_1 FILLER_59_121 ();
 sg13g2_decap_8 FILLER_59_138 ();
 sg13g2_decap_4 FILLER_59_145 ();
 sg13g2_fill_1 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_decap_8 FILLER_59_169 ();
 sg13g2_decap_4 FILLER_59_176 ();
 sg13g2_fill_2 FILLER_59_180 ();
 sg13g2_fill_1 FILLER_59_203 ();
 sg13g2_fill_1 FILLER_59_233 ();
 sg13g2_decap_8 FILLER_59_249 ();
 sg13g2_fill_2 FILLER_59_256 ();
 sg13g2_fill_1 FILLER_59_258 ();
 sg13g2_fill_2 FILLER_59_262 ();
 sg13g2_fill_1 FILLER_59_264 ();
 sg13g2_fill_2 FILLER_59_281 ();
 sg13g2_fill_1 FILLER_59_283 ();
 sg13g2_fill_1 FILLER_59_288 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_4 FILLER_59_308 ();
 sg13g2_fill_1 FILLER_59_312 ();
 sg13g2_fill_2 FILLER_59_325 ();
 sg13g2_fill_1 FILLER_59_350 ();
 sg13g2_fill_2 FILLER_59_376 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_48 ();
 sg13g2_fill_1 FILLER_60_50 ();
 sg13g2_decap_4 FILLER_60_71 ();
 sg13g2_decap_8 FILLER_60_85 ();
 sg13g2_decap_4 FILLER_60_92 ();
 sg13g2_fill_1 FILLER_60_148 ();
 sg13g2_fill_2 FILLER_60_174 ();
 sg13g2_decap_8 FILLER_60_180 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_decap_4 FILLER_60_194 ();
 sg13g2_fill_2 FILLER_60_198 ();
 sg13g2_decap_8 FILLER_60_204 ();
 sg13g2_decap_4 FILLER_60_211 ();
 sg13g2_fill_1 FILLER_60_215 ();
 sg13g2_decap_8 FILLER_60_240 ();
 sg13g2_decap_4 FILLER_60_247 ();
 sg13g2_decap_8 FILLER_60_256 ();
 sg13g2_fill_2 FILLER_60_263 ();
 sg13g2_decap_4 FILLER_60_309 ();
 sg13g2_fill_1 FILLER_60_313 ();
 sg13g2_fill_2 FILLER_60_323 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_fill_1 FILLER_60_359 ();
 sg13g2_fill_2 FILLER_60_371 ();
 sg13g2_fill_1 FILLER_60_373 ();
 sg13g2_fill_1 FILLER_60_391 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_14 ();
 sg13g2_fill_1 FILLER_61_56 ();
 sg13g2_fill_1 FILLER_61_66 ();
 sg13g2_decap_4 FILLER_61_83 ();
 sg13g2_decap_4 FILLER_61_117 ();
 sg13g2_fill_2 FILLER_61_121 ();
 sg13g2_fill_2 FILLER_61_132 ();
 sg13g2_fill_1 FILLER_61_134 ();
 sg13g2_fill_2 FILLER_61_180 ();
 sg13g2_decap_8 FILLER_61_204 ();
 sg13g2_fill_2 FILLER_61_211 ();
 sg13g2_fill_1 FILLER_61_213 ();
 sg13g2_decap_4 FILLER_61_228 ();
 sg13g2_fill_2 FILLER_61_232 ();
 sg13g2_fill_2 FILLER_61_287 ();
 sg13g2_fill_1 FILLER_61_303 ();
 sg13g2_decap_4 FILLER_61_335 ();
 sg13g2_fill_2 FILLER_61_339 ();
 sg13g2_decap_4 FILLER_61_351 ();
 sg13g2_fill_1 FILLER_61_355 ();
 sg13g2_fill_1 FILLER_61_364 ();
 sg13g2_fill_2 FILLER_61_369 ();
 sg13g2_fill_2 FILLER_61_381 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_4 FILLER_62_28 ();
 sg13g2_fill_2 FILLER_62_32 ();
 sg13g2_decap_4 FILLER_62_69 ();
 sg13g2_fill_1 FILLER_62_73 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_137 ();
 sg13g2_fill_1 FILLER_62_144 ();
 sg13g2_decap_4 FILLER_62_149 ();
 sg13g2_decap_4 FILLER_62_158 ();
 sg13g2_decap_8 FILLER_62_211 ();
 sg13g2_fill_2 FILLER_62_218 ();
 sg13g2_fill_1 FILLER_62_220 ();
 sg13g2_fill_1 FILLER_62_226 ();
 sg13g2_decap_8 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_253 ();
 sg13g2_decap_8 FILLER_62_258 ();
 sg13g2_decap_4 FILLER_62_265 ();
 sg13g2_decap_4 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_323 ();
 sg13g2_decap_4 FILLER_62_330 ();
 sg13g2_fill_2 FILLER_62_334 ();
 sg13g2_decap_4 FILLER_62_355 ();
 sg13g2_fill_1 FILLER_62_397 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_35 ();
 sg13g2_fill_2 FILLER_63_50 ();
 sg13g2_decap_4 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_95 ();
 sg13g2_decap_8 FILLER_63_102 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_decap_8 FILLER_63_116 ();
 sg13g2_fill_2 FILLER_63_123 ();
 sg13g2_fill_1 FILLER_63_125 ();
 sg13g2_decap_4 FILLER_63_134 ();
 sg13g2_fill_1 FILLER_63_190 ();
 sg13g2_decap_8 FILLER_63_195 ();
 sg13g2_decap_8 FILLER_63_202 ();
 sg13g2_fill_2 FILLER_63_209 ();
 sg13g2_fill_1 FILLER_63_211 ();
 sg13g2_fill_1 FILLER_63_231 ();
 sg13g2_fill_1 FILLER_63_251 ();
 sg13g2_fill_1 FILLER_63_260 ();
 sg13g2_fill_1 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_330 ();
 sg13g2_decap_4 FILLER_63_337 ();
 sg13g2_fill_1 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_350 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_14 ();
 sg13g2_decap_4 FILLER_64_55 ();
 sg13g2_fill_2 FILLER_64_59 ();
 sg13g2_decap_4 FILLER_64_64 ();
 sg13g2_fill_1 FILLER_64_81 ();
 sg13g2_fill_1 FILLER_64_92 ();
 sg13g2_decap_8 FILLER_64_108 ();
 sg13g2_fill_2 FILLER_64_115 ();
 sg13g2_decap_4 FILLER_64_126 ();
 sg13g2_fill_2 FILLER_64_130 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_4 FILLER_64_147 ();
 sg13g2_fill_2 FILLER_64_151 ();
 sg13g2_decap_8 FILLER_64_157 ();
 sg13g2_decap_4 FILLER_64_164 ();
 sg13g2_fill_1 FILLER_64_168 ();
 sg13g2_fill_1 FILLER_64_174 ();
 sg13g2_decap_8 FILLER_64_179 ();
 sg13g2_decap_8 FILLER_64_186 ();
 sg13g2_decap_8 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_200 ();
 sg13g2_fill_1 FILLER_64_206 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_fill_1 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_352 ();
 sg13g2_fill_1 FILLER_64_359 ();
 sg13g2_fill_2 FILLER_64_386 ();
 sg13g2_fill_1 FILLER_64_388 ();
 sg13g2_decap_8 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_62 ();
 sg13g2_decap_8 FILLER_65_69 ();
 sg13g2_decap_8 FILLER_65_134 ();
 sg13g2_decap_4 FILLER_65_193 ();
 sg13g2_fill_1 FILLER_65_197 ();
 sg13g2_fill_2 FILLER_65_215 ();
 sg13g2_fill_2 FILLER_65_237 ();
 sg13g2_fill_2 FILLER_65_245 ();
 sg13g2_fill_2 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_260 ();
 sg13g2_decap_4 FILLER_65_266 ();
 sg13g2_fill_2 FILLER_65_270 ();
 sg13g2_decap_8 FILLER_65_276 ();
 sg13g2_decap_4 FILLER_65_283 ();
 sg13g2_fill_2 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_302 ();
 sg13g2_fill_2 FILLER_65_322 ();
 sg13g2_fill_1 FILLER_65_324 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_decap_4 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_339 ();
 sg13g2_fill_2 FILLER_65_380 ();
 sg13g2_fill_1 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_4 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_25 ();
 sg13g2_fill_2 FILLER_66_79 ();
 sg13g2_fill_1 FILLER_66_81 ();
 sg13g2_fill_2 FILLER_66_125 ();
 sg13g2_fill_1 FILLER_66_127 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_fill_2 FILLER_66_175 ();
 sg13g2_fill_1 FILLER_66_177 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_fill_2 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_decap_8 FILLER_66_247 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_decap_8 FILLER_66_261 ();
 sg13g2_decap_8 FILLER_66_276 ();
 sg13g2_fill_1 FILLER_66_283 ();
 sg13g2_fill_2 FILLER_66_297 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_327 ();
 sg13g2_fill_1 FILLER_66_349 ();
 sg13g2_decap_8 FILLER_66_363 ();
 sg13g2_decap_8 FILLER_66_370 ();
 sg13g2_decap_4 FILLER_66_377 ();
 sg13g2_decap_4 FILLER_66_389 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_23 ();
 sg13g2_fill_2 FILLER_67_79 ();
 sg13g2_decap_4 FILLER_67_102 ();
 sg13g2_decap_8 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_128 ();
 sg13g2_fill_2 FILLER_67_145 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_157 ();
 sg13g2_decap_8 FILLER_67_164 ();
 sg13g2_decap_4 FILLER_67_171 ();
 sg13g2_fill_2 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_4 FILLER_67_238 ();
 sg13g2_decap_4 FILLER_67_250 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_fill_2 FILLER_67_286 ();
 sg13g2_decap_8 FILLER_67_362 ();
 sg13g2_decap_4 FILLER_67_369 ();
 sg13g2_decap_4 FILLER_67_390 ();
 sg13g2_fill_1 FILLER_67_394 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_fill_1 FILLER_68_44 ();
 sg13g2_fill_2 FILLER_68_50 ();
 sg13g2_fill_1 FILLER_68_52 ();
 sg13g2_decap_4 FILLER_68_72 ();
 sg13g2_decap_8 FILLER_68_81 ();
 sg13g2_fill_2 FILLER_68_88 ();
 sg13g2_fill_1 FILLER_68_90 ();
 sg13g2_fill_1 FILLER_68_96 ();
 sg13g2_decap_8 FILLER_68_107 ();
 sg13g2_decap_8 FILLER_68_114 ();
 sg13g2_decap_8 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_141 ();
 sg13g2_fill_1 FILLER_68_143 ();
 sg13g2_decap_8 FILLER_68_152 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_8 FILLER_68_166 ();
 sg13g2_decap_8 FILLER_68_173 ();
 sg13g2_fill_1 FILLER_68_180 ();
 sg13g2_decap_8 FILLER_68_207 ();
 sg13g2_decap_8 FILLER_68_214 ();
 sg13g2_decap_8 FILLER_68_221 ();
 sg13g2_decap_4 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_241 ();
 sg13g2_fill_1 FILLER_68_243 ();
 sg13g2_fill_2 FILLER_68_251 ();
 sg13g2_fill_1 FILLER_68_253 ();
 sg13g2_fill_2 FILLER_68_273 ();
 sg13g2_fill_1 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_358 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_fill_1 FILLER_68_373 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_4 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_39 ();
 sg13g2_decap_8 FILLER_69_58 ();
 sg13g2_fill_2 FILLER_69_65 ();
 sg13g2_decap_8 FILLER_69_79 ();
 sg13g2_decap_8 FILLER_69_86 ();
 sg13g2_decap_8 FILLER_69_93 ();
 sg13g2_decap_8 FILLER_69_100 ();
 sg13g2_fill_2 FILLER_69_107 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_fill_1 FILLER_69_137 ();
 sg13g2_fill_2 FILLER_69_143 ();
 sg13g2_fill_2 FILLER_69_158 ();
 sg13g2_fill_1 FILLER_69_160 ();
 sg13g2_fill_1 FILLER_69_182 ();
 sg13g2_fill_2 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_193 ();
 sg13g2_decap_8 FILLER_69_220 ();
 sg13g2_fill_1 FILLER_69_227 ();
 sg13g2_fill_2 FILLER_69_280 ();
 sg13g2_fill_2 FILLER_69_321 ();
 sg13g2_fill_1 FILLER_69_382 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_21 ();
 sg13g2_fill_1 FILLER_70_25 ();
 sg13g2_fill_2 FILLER_70_62 ();
 sg13g2_decap_8 FILLER_70_88 ();
 sg13g2_decap_4 FILLER_70_95 ();
 sg13g2_fill_1 FILLER_70_99 ();
 sg13g2_fill_1 FILLER_70_130 ();
 sg13g2_fill_1 FILLER_70_140 ();
 sg13g2_fill_2 FILLER_70_150 ();
 sg13g2_fill_2 FILLER_70_168 ();
 sg13g2_fill_2 FILLER_70_180 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_fill_1 FILLER_70_301 ();
 sg13g2_fill_1 FILLER_70_315 ();
 sg13g2_decap_4 FILLER_70_349 ();
 sg13g2_fill_2 FILLER_70_383 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_4 FILLER_71_28 ();
 sg13g2_fill_2 FILLER_71_32 ();
 sg13g2_fill_2 FILLER_71_64 ();
 sg13g2_fill_2 FILLER_71_92 ();
 sg13g2_fill_1 FILLER_71_94 ();
 sg13g2_fill_2 FILLER_71_109 ();
 sg13g2_fill_2 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_183 ();
 sg13g2_decap_8 FILLER_71_218 ();
 sg13g2_decap_8 FILLER_71_225 ();
 sg13g2_decap_8 FILLER_71_232 ();
 sg13g2_decap_4 FILLER_71_239 ();
 sg13g2_decap_8 FILLER_71_250 ();
 sg13g2_decap_8 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_264 ();
 sg13g2_fill_2 FILLER_71_277 ();
 sg13g2_decap_8 FILLER_71_283 ();
 sg13g2_decap_4 FILLER_71_298 ();
 sg13g2_fill_2 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_308 ();
 sg13g2_fill_2 FILLER_71_316 ();
 sg13g2_fill_2 FILLER_71_325 ();
 sg13g2_fill_2 FILLER_71_332 ();
 sg13g2_decap_8 FILLER_71_338 ();
 sg13g2_decap_8 FILLER_71_345 ();
 sg13g2_decap_8 FILLER_71_352 ();
 sg13g2_fill_1 FILLER_71_359 ();
 sg13g2_fill_1 FILLER_71_364 ();
 sg13g2_fill_2 FILLER_71_375 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_fill_2 FILLER_71_397 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_35 ();
 sg13g2_fill_1 FILLER_72_59 ();
 sg13g2_fill_1 FILLER_72_125 ();
 sg13g2_fill_2 FILLER_72_130 ();
 sg13g2_decap_4 FILLER_72_174 ();
 sg13g2_decap_4 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_212 ();
 sg13g2_decap_8 FILLER_72_219 ();
 sg13g2_decap_8 FILLER_72_226 ();
 sg13g2_decap_4 FILLER_72_233 ();
 sg13g2_decap_8 FILLER_72_277 ();
 sg13g2_fill_2 FILLER_72_284 ();
 sg13g2_decap_8 FILLER_72_292 ();
 sg13g2_fill_2 FILLER_72_299 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_decap_4 FILLER_72_333 ();
 sg13g2_fill_1 FILLER_72_337 ();
 sg13g2_decap_8 FILLER_72_342 ();
 sg13g2_decap_8 FILLER_72_355 ();
 sg13g2_decap_8 FILLER_72_362 ();
 sg13g2_fill_2 FILLER_72_369 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_66 ();
 sg13g2_fill_1 FILLER_73_103 ();
 sg13g2_fill_2 FILLER_73_117 ();
 sg13g2_fill_2 FILLER_73_128 ();
 sg13g2_fill_1 FILLER_73_130 ();
 sg13g2_fill_1 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_173 ();
 sg13g2_decap_8 FILLER_73_180 ();
 sg13g2_decap_8 FILLER_73_187 ();
 sg13g2_fill_2 FILLER_73_194 ();
 sg13g2_fill_1 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_205 ();
 sg13g2_decap_8 FILLER_73_212 ();
 sg13g2_decap_8 FILLER_73_219 ();
 sg13g2_decap_4 FILLER_73_226 ();
 sg13g2_fill_1 FILLER_73_274 ();
 sg13g2_fill_2 FILLER_73_314 ();
 sg13g2_fill_2 FILLER_73_330 ();
 sg13g2_fill_2 FILLER_73_363 ();
 sg13g2_fill_2 FILLER_73_386 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_4 FILLER_74_49 ();
 sg13g2_fill_1 FILLER_74_53 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_84 ();
 sg13g2_fill_2 FILLER_74_129 ();
 sg13g2_fill_1 FILLER_74_152 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_4 FILLER_74_203 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_235 ();
 sg13g2_fill_1 FILLER_74_242 ();
 sg13g2_fill_2 FILLER_74_257 ();
 sg13g2_decap_4 FILLER_74_293 ();
 sg13g2_fill_2 FILLER_74_297 ();
 sg13g2_fill_2 FILLER_74_318 ();
 sg13g2_fill_2 FILLER_74_334 ();
 sg13g2_fill_2 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_4 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_82 ();
 sg13g2_decap_8 FILLER_75_131 ();
 sg13g2_fill_2 FILLER_75_138 ();
 sg13g2_decap_8 FILLER_75_143 ();
 sg13g2_decap_4 FILLER_75_154 ();
 sg13g2_fill_1 FILLER_75_158 ();
 sg13g2_decap_8 FILLER_75_163 ();
 sg13g2_decap_4 FILLER_75_170 ();
 sg13g2_decap_8 FILLER_75_181 ();
 sg13g2_decap_8 FILLER_75_188 ();
 sg13g2_decap_8 FILLER_75_195 ();
 sg13g2_fill_2 FILLER_75_202 ();
 sg13g2_decap_8 FILLER_75_258 ();
 sg13g2_fill_2 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_4 FILLER_75_287 ();
 sg13g2_fill_2 FILLER_75_295 ();
 sg13g2_fill_1 FILLER_75_297 ();
 sg13g2_fill_2 FILLER_75_303 ();
 sg13g2_decap_8 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_fill_1 FILLER_75_342 ();
 sg13g2_decap_4 FILLER_75_347 ();
 sg13g2_fill_1 FILLER_75_351 ();
 sg13g2_decap_4 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_360 ();
 sg13g2_fill_1 FILLER_75_369 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_4 FILLER_76_35 ();
 sg13g2_fill_2 FILLER_76_81 ();
 sg13g2_fill_2 FILLER_76_129 ();
 sg13g2_fill_2 FILLER_76_145 ();
 sg13g2_fill_2 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_195 ();
 sg13g2_decap_8 FILLER_76_202 ();
 sg13g2_decap_4 FILLER_76_209 ();
 sg13g2_fill_1 FILLER_76_213 ();
 sg13g2_fill_1 FILLER_76_260 ();
 sg13g2_fill_2 FILLER_76_269 ();
 sg13g2_fill_1 FILLER_76_271 ();
 sg13g2_decap_8 FILLER_76_281 ();
 sg13g2_decap_4 FILLER_76_288 ();
 sg13g2_fill_2 FILLER_76_292 ();
 sg13g2_fill_1 FILLER_76_307 ();
 sg13g2_decap_8 FILLER_76_328 ();
 sg13g2_decap_4 FILLER_76_335 ();
 sg13g2_fill_2 FILLER_76_339 ();
 sg13g2_fill_2 FILLER_76_362 ();
 sg13g2_fill_1 FILLER_76_375 ();
 sg13g2_fill_1 FILLER_76_383 ();
 sg13g2_fill_2 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_4 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_46 ();
 sg13g2_fill_1 FILLER_77_83 ();
 sg13g2_fill_1 FILLER_77_98 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_fill_2 FILLER_77_217 ();
 sg13g2_fill_1 FILLER_77_219 ();
 sg13g2_fill_1 FILLER_77_224 ();
 sg13g2_fill_2 FILLER_77_258 ();
 sg13g2_fill_2 FILLER_77_302 ();
 sg13g2_fill_1 FILLER_77_304 ();
 sg13g2_fill_1 FILLER_77_314 ();
 sg13g2_decap_4 FILLER_77_344 ();
 sg13g2_fill_2 FILLER_77_348 ();
 sg13g2_decap_4 FILLER_77_360 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_fill_1 FILLER_78_49 ();
 sg13g2_decap_4 FILLER_78_127 ();
 sg13g2_decap_4 FILLER_78_205 ();
 sg13g2_fill_1 FILLER_78_209 ();
 sg13g2_fill_2 FILLER_78_263 ();
 sg13g2_fill_1 FILLER_78_265 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_4 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_53 ();
 sg13g2_fill_2 FILLER_79_63 ();
 sg13g2_fill_1 FILLER_79_65 ();
 sg13g2_fill_2 FILLER_79_110 ();
 sg13g2_decap_8 FILLER_79_142 ();
 sg13g2_decap_8 FILLER_79_149 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_fill_1 FILLER_79_189 ();
 sg13g2_decap_4 FILLER_79_198 ();
 sg13g2_fill_1 FILLER_79_242 ();
 sg13g2_fill_2 FILLER_79_248 ();
 sg13g2_fill_1 FILLER_79_250 ();
 sg13g2_fill_1 FILLER_79_312 ();
 sg13g2_fill_2 FILLER_79_344 ();
 sg13g2_fill_1 FILLER_79_346 ();
 sg13g2_fill_1 FILLER_79_382 ();
 sg13g2_fill_1 FILLER_79_392 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_fill_2 FILLER_80_49 ();
 sg13g2_fill_1 FILLER_80_84 ();
 sg13g2_fill_1 FILLER_80_103 ();
 sg13g2_fill_2 FILLER_80_116 ();
 sg13g2_fill_1 FILLER_80_118 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_8 FILLER_80_140 ();
 sg13g2_decap_8 FILLER_80_147 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_4 FILLER_80_161 ();
 sg13g2_fill_2 FILLER_80_165 ();
 sg13g2_decap_8 FILLER_80_171 ();
 sg13g2_decap_8 FILLER_80_178 ();
 sg13g2_decap_8 FILLER_80_185 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_217 ();
 sg13g2_decap_4 FILLER_80_237 ();
 sg13g2_decap_4 FILLER_80_245 ();
 sg13g2_fill_1 FILLER_80_249 ();
 sg13g2_decap_4 FILLER_80_260 ();
 sg13g2_fill_1 FILLER_80_264 ();
 sg13g2_decap_4 FILLER_80_270 ();
 sg13g2_decap_4 FILLER_80_278 ();
 sg13g2_fill_2 FILLER_80_282 ();
 sg13g2_decap_8 FILLER_80_288 ();
 sg13g2_decap_8 FILLER_80_295 ();
 sg13g2_fill_1 FILLER_80_302 ();
 sg13g2_fill_2 FILLER_80_341 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_356 ();
 sg13g2_fill_2 FILLER_80_372 ();
 sg13g2_fill_1 FILLER_80_374 ();
 sg13g2_fill_2 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net215;
 assign uio_oe[1] = net216;
 assign uio_oe[2] = net217;
 assign uio_oe[3] = net218;
 assign uio_oe[4] = net219;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[5] = net10;
 assign uio_out[6] = net11;
 assign uio_out[7] = net12;
endmodule
