module tt_um_a1k0n_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire audio;
 wire hsync;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire \vgademo.a_cos[0] ;
 wire \vgademo.a_cos[10] ;
 wire \vgademo.a_cos[11] ;
 wire \vgademo.a_cos[12] ;
 wire \vgademo.a_cos[13] ;
 wire \vgademo.a_cos[14] ;
 wire \vgademo.a_cos[1] ;
 wire \vgademo.a_cos[2] ;
 wire \vgademo.a_cos[3] ;
 wire \vgademo.a_cos[4] ;
 wire \vgademo.a_cos[5] ;
 wire \vgademo.a_cos[6] ;
 wire \vgademo.a_cos[7] ;
 wire \vgademo.a_cos[8] ;
 wire \vgademo.a_cos[9] ;
 wire \vgademo.a_scrolly[10] ;
 wire \vgademo.a_scrolly[11] ;
 wire \vgademo.a_scrolly[12] ;
 wire \vgademo.a_scrolly[13] ;
 wire \vgademo.a_scrolly[3] ;
 wire \vgademo.a_scrolly[4] ;
 wire \vgademo.a_scrolly[5] ;
 wire \vgademo.a_scrolly[6] ;
 wire \vgademo.a_scrolly[7] ;
 wire \vgademo.a_scrolly[8] ;
 wire \vgademo.a_scrolly[9] ;
 wire \vgademo.a_sin[0] ;
 wire \vgademo.a_sin[10] ;
 wire \vgademo.a_sin[11] ;
 wire \vgademo.a_sin[12] ;
 wire \vgademo.a_sin[13] ;
 wire \vgademo.a_sin[14] ;
 wire \vgademo.a_sin[1] ;
 wire \vgademo.a_sin[2] ;
 wire \vgademo.a_sin[3] ;
 wire \vgademo.a_sin[4] ;
 wire \vgademo.a_sin[5] ;
 wire \vgademo.a_sin[6] ;
 wire \vgademo.a_sin[7] ;
 wire \vgademo.a_sin[8] ;
 wire \vgademo.a_sin[9] ;
 wire \vgademo.audio_beat_out[0] ;
 wire \vgademo.audio_beat_out[1] ;
 wire \vgademo.audio_beat_out[2] ;
 wire \vgademo.audio_beat_out[3] ;
 wire \vgademo.audio_beat_out[4] ;
 wire \vgademo.audio_kick_frames[0] ;
 wire \vgademo.audio_kick_frames[1] ;
 wire \vgademo.audio_kick_frames[2] ;
 wire \vgademo.audio_snare_frames[0] ;
 wire \vgademo.audio_snare_frames[1] ;
 wire \vgademo.audio_snare_frames[2] ;
 wire \vgademo.audio_snare_frames[3] ;
 wire \vgademo.audio_songpos[0] ;
 wire \vgademo.audio_songpos[1] ;
 wire \vgademo.audio_songpos[2] ;
 wire \vgademo.audio_songpos[3] ;
 wire \vgademo.audio_songpos[4] ;
 wire \vgademo.audio_songpos[5] ;
 wire \vgademo.audio_songpos[6] ;
 wire \vgademo.audio_songpos[7] ;
 wire \vgademo.b_cos[0] ;
 wire \vgademo.b_cos[10] ;
 wire \vgademo.b_cos[11] ;
 wire \vgademo.b_cos[1] ;
 wire \vgademo.b_cos[2] ;
 wire \vgademo.b_cos[3] ;
 wire \vgademo.b_cos[4] ;
 wire \vgademo.b_cos[5] ;
 wire \vgademo.b_cos[6] ;
 wire \vgademo.b_cos[7] ;
 wire \vgademo.b_cos[8] ;
 wire \vgademo.b_cos[9] ;
 wire \vgademo.b_sin[0] ;
 wire \vgademo.b_sin[10] ;
 wire \vgademo.b_sin[11] ;
 wire \vgademo.b_sin[1] ;
 wire \vgademo.b_sin[2] ;
 wire \vgademo.b_sin[3] ;
 wire \vgademo.b_sin[4] ;
 wire \vgademo.b_sin[5] ;
 wire \vgademo.b_sin[6] ;
 wire \vgademo.b_sin[7] ;
 wire \vgademo.b_sin[8] ;
 wire \vgademo.b_sin[9] ;
 wire \vgademo.bayer_j[0] ;
 wire \vgademo.bayer_j[1] ;
 wire \vgademo.h_count[0] ;
 wire \vgademo.h_count[10] ;
 wire \vgademo.h_count[1] ;
 wire \vgademo.h_count[2] ;
 wire \vgademo.h_count[3] ;
 wire \vgademo.h_count[4] ;
 wire \vgademo.h_count[5] ;
 wire \vgademo.h_count[6] ;
 wire \vgademo.h_count[7] ;
 wire \vgademo.h_count[8] ;
 wire \vgademo.h_count[9] ;
 wire \vgademo.linelfsr[0] ;
 wire \vgademo.linelfsr[10] ;
 wire \vgademo.linelfsr[11] ;
 wire \vgademo.linelfsr[12] ;
 wire \vgademo.linelfsr[1] ;
 wire \vgademo.linelfsr[2] ;
 wire \vgademo.linelfsr[3] ;
 wire \vgademo.linelfsr[4] ;
 wire \vgademo.linelfsr[5] ;
 wire \vgademo.linelfsr[6] ;
 wire \vgademo.linelfsr[7] ;
 wire \vgademo.linelfsr[8] ;
 wire \vgademo.linelfsr[9] ;
 wire \vgademo.plane_du[0] ;
 wire \vgademo.plane_du[10] ;
 wire \vgademo.plane_du[1] ;
 wire \vgademo.plane_du[2] ;
 wire \vgademo.plane_du[3] ;
 wire \vgademo.plane_du[4] ;
 wire \vgademo.plane_du[5] ;
 wire \vgademo.plane_du[6] ;
 wire \vgademo.plane_du[7] ;
 wire \vgademo.plane_du[8] ;
 wire \vgademo.plane_du[9] ;
 wire \vgademo.plane_dx[0] ;
 wire \vgademo.plane_dx[1] ;
 wire \vgademo.plane_dx[2] ;
 wire \vgademo.plane_dx[3] ;
 wire \vgademo.plane_dx_div.d[16] ;
 wire \vgademo.plane_dx_div.d[17] ;
 wire \vgademo.plane_dx_div.d[18] ;
 wire \vgademo.plane_dx_div.d[19] ;
 wire \vgademo.plane_dx_div.d[20] ;
 wire \vgademo.plane_dx_div.d[21] ;
 wire \vgademo.plane_dx_div.d[22] ;
 wire \vgademo.plane_dx_div.d[23] ;
 wire \vgademo.plane_dx_div.d[24] ;
 wire \vgademo.plane_dx_div.i[0] ;
 wire \vgademo.plane_dx_div.i[1] ;
 wire \vgademo.plane_dx_div.i[2] ;
 wire \vgademo.plane_dx_div.i[3] ;
 wire \vgademo.plane_dx_div.q[3] ;
 wire \vgademo.plane_dx_div.q[4] ;
 wire \vgademo.plane_dx_div.q[5] ;
 wire \vgademo.plane_dx_div.q[6] ;
 wire \vgademo.plane_dx_div.q[7] ;
 wire \vgademo.plane_dx_div.q[8] ;
 wire \vgademo.plane_dx_div.q[9] ;
 wire \vgademo.plane_dx_div.r[16] ;
 wire \vgademo.plane_dx_div.r[17] ;
 wire \vgademo.plane_dx_div.r[18] ;
 wire \vgademo.plane_dx_div.r[19] ;
 wire \vgademo.plane_dx_div.r[20] ;
 wire \vgademo.plane_dx_div.r[21] ;
 wire \vgademo.plane_dx_div.r[22] ;
 wire \vgademo.plane_dx_div.r[23] ;
 wire \vgademo.plane_dx_div.r[24] ;
 wire \vgademo.plane_dx_div.r[25] ;
 wire \vgademo.plane_u[0] ;
 wire \vgademo.plane_u[10] ;
 wire \vgademo.plane_u[11] ;
 wire \vgademo.plane_u[12] ;
 wire \vgademo.plane_u[13] ;
 wire \vgademo.plane_u[14] ;
 wire \vgademo.plane_u[15] ;
 wire \vgademo.plane_u[16] ;
 wire \vgademo.plane_u[17] ;
 wire \vgademo.plane_u[18] ;
 wire \vgademo.plane_u[19] ;
 wire \vgademo.plane_u[1] ;
 wire \vgademo.plane_u[20] ;
 wire \vgademo.plane_u[21] ;
 wire \vgademo.plane_u[2] ;
 wire \vgademo.plane_u[3] ;
 wire \vgademo.plane_u[4] ;
 wire \vgademo.plane_u[5] ;
 wire \vgademo.plane_u[6] ;
 wire \vgademo.plane_u[7] ;
 wire \vgademo.plane_u[8] ;
 wire \vgademo.plane_u[9] ;
 wire \vgademo.scanline_audio_sample[0] ;
 wire \vgademo.scanline_audio_sample[1] ;
 wire \vgademo.scanline_audio_sample[2] ;
 wire \vgademo.scanline_audio_sample[3] ;
 wire \vgademo.scanline_audio_sample[4] ;
 wire \vgademo.scanline_audio_sample[5] ;
 wire \vgademo.scanline_audio_sample[6] ;
 wire \vgademo.soundtrack.noise_lfsr[0] ;
 wire \vgademo.soundtrack.noise_lfsr[10] ;
 wire \vgademo.soundtrack.noise_lfsr[11] ;
 wire \vgademo.soundtrack.noise_lfsr[12] ;
 wire \vgademo.soundtrack.noise_lfsr[13] ;
 wire \vgademo.soundtrack.noise_lfsr[14] ;
 wire \vgademo.soundtrack.noise_lfsr[1] ;
 wire \vgademo.soundtrack.noise_lfsr[2] ;
 wire \vgademo.soundtrack.noise_lfsr[3] ;
 wire \vgademo.soundtrack.noise_lfsr[4] ;
 wire \vgademo.soundtrack.noise_lfsr[5] ;
 wire \vgademo.soundtrack.noise_lfsr[6] ;
 wire \vgademo.soundtrack.noise_lfsr[7] ;
 wire \vgademo.soundtrack.noise_lfsr[8] ;
 wire \vgademo.soundtrack.noise_lfsr[9] ;
 wire \vgademo.soundtrack.pulse_osc_p[0] ;
 wire \vgademo.soundtrack.pulse_osc_p[10] ;
 wire \vgademo.soundtrack.pulse_osc_p[11] ;
 wire \vgademo.soundtrack.pulse_osc_p[12] ;
 wire \vgademo.soundtrack.pulse_osc_p[13] ;
 wire \vgademo.soundtrack.pulse_osc_p[1] ;
 wire \vgademo.soundtrack.pulse_osc_p[2] ;
 wire \vgademo.soundtrack.pulse_osc_p[3] ;
 wire \vgademo.soundtrack.pulse_osc_p[4] ;
 wire \vgademo.soundtrack.pulse_osc_p[5] ;
 wire \vgademo.soundtrack.pulse_osc_p[6] ;
 wire \vgademo.soundtrack.pulse_osc_p[7] ;
 wire \vgademo.soundtrack.pulse_osc_p[8] ;
 wire \vgademo.soundtrack.pulse_osc_p[9] ;
 wire \vgademo.soundtrack.pulse_vol[0] ;
 wire \vgademo.soundtrack.pulse_vol[1] ;
 wire \vgademo.soundtrack.pulse_vol[2] ;
 wire \vgademo.soundtrack.pulse_vol[3] ;
 wire \vgademo.soundtrack.sample_div[0] ;
 wire \vgademo.soundtrack.sample_div[1] ;
 wire \vgademo.soundtrack.sample_div[2] ;
 wire \vgademo.soundtrack.sample_div[3] ;
 wire \vgademo.soundtrack.sample_div[4] ;
 wire \vgademo.soundtrack.sample_div[5] ;
 wire \vgademo.soundtrack.sample_div[6] ;
 wire \vgademo.soundtrack.sample_div[7] ;
 wire \vgademo.soundtrack.sample_div[8] ;
 wire \vgademo.soundtrack.sample_div[9] ;
 wire \vgademo.soundtrack.sample_div_[0] ;
 wire \vgademo.soundtrack.sample_div_[1] ;
 wire \vgademo.soundtrack.sample_div_[2] ;
 wire \vgademo.soundtrack.sample_div_[3] ;
 wire \vgademo.soundtrack.sample_div_[4] ;
 wire \vgademo.soundtrack.sample_div_[5] ;
 wire \vgademo.soundtrack.sample_div_[6] ;
 wire \vgademo.soundtrack.sample_div_[7] ;
 wire \vgademo.soundtrack.sample_div_[8] ;
 wire \vgademo.soundtrack.sample_div_[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[9] ;
 wire \vgademo.soundtrack.tick_div[0] ;
 wire \vgademo.soundtrack.tick_div[1] ;
 wire \vgademo.soundtrack.tick_div[2] ;
 wire \vgademo.soundtrack.tick_div[3] ;
 wire \vgademo.soundtrack.tick_div[4] ;
 wire \vgademo.soundtrack.tick_div[5] ;
 wire \vgademo.soundtrack.tick_div[6] ;
 wire \vgademo.soundtrack.tick_div[7] ;
 wire \vgademo.soundtrack.tick_div_[0] ;
 wire \vgademo.soundtrack.tri_osc_i[0] ;
 wire \vgademo.soundtrack.tri_osc_i[1] ;
 wire \vgademo.soundtrack.tri_osc_i[2] ;
 wire \vgademo.soundtrack.tri_osc_i[3] ;
 wire \vgademo.soundtrack.tri_osc_i[4] ;
 wire \vgademo.soundtrack.tri_osc_i[5] ;
 wire \vgademo.soundtrack.tri_osc_i[6] ;
 wire \vgademo.soundtrack.tri_osc_i[7] ;
 wire \vgademo.soundtrack.tri_osc_i[8] ;
 wire \vgademo.soundtrack.tri_osc_p[0] ;
 wire \vgademo.soundtrack.tri_osc_p[10] ;
 wire \vgademo.soundtrack.tri_osc_p[11] ;
 wire \vgademo.soundtrack.tri_osc_p[12] ;
 wire \vgademo.soundtrack.tri_osc_p[13] ;
 wire \vgademo.soundtrack.tri_osc_p[14] ;
 wire \vgademo.soundtrack.tri_osc_p[15] ;
 wire \vgademo.soundtrack.tri_osc_p[1] ;
 wire \vgademo.soundtrack.tri_osc_p[2] ;
 wire \vgademo.soundtrack.tri_osc_p[3] ;
 wire \vgademo.soundtrack.tri_osc_p[4] ;
 wire \vgademo.soundtrack.tri_osc_p[5] ;
 wire \vgademo.soundtrack.tri_osc_p[6] ;
 wire \vgademo.soundtrack.tri_osc_p[7] ;
 wire \vgademo.soundtrack.tri_osc_p[8] ;
 wire \vgademo.soundtrack.tri_osc_p[9] ;
 wire \vgademo.v_count[2] ;
 wire \vgademo.v_count[3] ;
 wire \vgademo.v_count[4] ;
 wire \vgademo.v_count[5] ;
 wire \vgademo.v_count[6] ;
 wire \vgademo.v_count[7] ;
 wire \vgademo.v_count[8] ;
 wire \vgademo.v_count[9] ;
 wire \vgademo.vsync ;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;

 sg13g2_inv_1 _3810_ (.Y(_3163_),
    .A(net211));
 sg13g2_inv_2 _3811_ (.Y(_3164_),
    .A(net351));
 sg13g2_inv_1 _3812_ (.Y(_3165_),
    .A(net531));
 sg13g2_inv_1 _3813_ (.Y(_3166_),
    .A(net544));
 sg13g2_inv_1 _3814_ (.Y(_3167_),
    .A(\vgademo.linelfsr[10] ));
 sg13g2_inv_1 _3815_ (.Y(_3168_),
    .A(\vgademo.linelfsr[6] ));
 sg13g2_inv_1 _3816_ (.Y(_3169_),
    .A(\vgademo.linelfsr[2] ));
 sg13g2_inv_2 _3817_ (.Y(_3170_),
    .A(net1151));
 sg13g2_inv_1 _3818_ (.Y(_3171_),
    .A(net512));
 sg13g2_inv_4 _3819_ (.A(net416),
    .Y(_3172_));
 sg13g2_inv_1 _3820_ (.Y(_3173_),
    .A(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_inv_1 _3821_ (.Y(_3174_),
    .A(net254));
 sg13g2_inv_1 _3822_ (.Y(_3175_),
    .A(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_inv_1 _3823_ (.Y(_3176_),
    .A(\vgademo.audio_beat_out[2] ));
 sg13g2_inv_2 _3824_ (.Y(_3177_),
    .A(net1137));
 sg13g2_inv_1 _3825_ (.Y(_3178_),
    .A(net1143));
 sg13g2_inv_1 _3826_ (.Y(_3179_),
    .A(net1145));
 sg13g2_inv_1 _3827_ (.Y(_3180_),
    .A(net1134));
 sg13g2_inv_1 _3828_ (.Y(_3181_),
    .A(net1132));
 sg13g2_inv_4 _3829_ (.A(_0059_),
    .Y(_3182_));
 sg13g2_inv_2 _3830_ (.Y(_3183_),
    .A(\vgademo.bayer_j[1] ));
 sg13g2_inv_2 _3831_ (.Y(_3184_),
    .A(\vgademo.bayer_j[0] ));
 sg13g2_inv_2 _3832_ (.Y(_3185_),
    .A(\vgademo.v_count[5] ));
 sg13g2_inv_1 _3833_ (.Y(_3186_),
    .A(net1061));
 sg13g2_inv_1 _3834_ (.Y(_3187_),
    .A(\vgademo.v_count[8] ));
 sg13g2_inv_1 _3835_ (.Y(_3188_),
    .A(net1096));
 sg13g2_inv_1 _3836_ (.Y(_3189_),
    .A(net1098));
 sg13g2_inv_1 _3837_ (.Y(_3190_),
    .A(net1094));
 sg13g2_inv_1 _3838_ (.Y(_3191_),
    .A(net1095));
 sg13g2_inv_4 _3839_ (.A(\vgademo.h_count[5] ),
    .Y(_3192_));
 sg13g2_inv_2 _3840_ (.Y(_3193_),
    .A(\vgademo.h_count[4] ));
 sg13g2_inv_1 _3841_ (.Y(_3194_),
    .A(\vgademo.h_count[7] ));
 sg13g2_inv_2 _3842_ (.Y(_3195_),
    .A(\vgademo.h_count[9] ));
 sg13g2_inv_2 _3843_ (.Y(_3196_),
    .A(net1067));
 sg13g2_inv_2 _3844_ (.Y(_3197_),
    .A(net1068));
 sg13g2_inv_2 _3845_ (.Y(_3198_),
    .A(net1076));
 sg13g2_inv_1 _3846_ (.Y(_3199_),
    .A(net1078));
 sg13g2_inv_2 _3847_ (.Y(_3200_),
    .A(net1081));
 sg13g2_inv_2 _3848_ (.Y(_3201_),
    .A(net1087));
 sg13g2_inv_1 _3849_ (.Y(_3202_),
    .A(_0063_));
 sg13g2_inv_1 _3850_ (.Y(_3203_),
    .A(net458));
 sg13g2_inv_2 _3851_ (.Y(_3204_),
    .A(_0068_));
 sg13g2_inv_1 _3852_ (.Y(_3205_),
    .A(net391));
 sg13g2_inv_1 _3853_ (.Y(_3206_),
    .A(net359));
 sg13g2_inv_1 _3854_ (.Y(_3207_),
    .A(net455));
 sg13g2_inv_1 _3855_ (.Y(_3208_),
    .A(\vgademo.plane_dx_div.r[20] ));
 sg13g2_inv_1 _3856_ (.Y(_3209_),
    .A(_0014_));
 sg13g2_inv_1 _3857_ (.Y(_3210_),
    .A(_0016_));
 sg13g2_inv_1 _3858_ (.Y(_3211_),
    .A(net383));
 sg13g2_inv_1 _3859_ (.Y(_3212_),
    .A(_0019_));
 sg13g2_inv_1 _3860_ (.Y(_3213_),
    .A(_0018_));
 sg13g2_inv_1 _3861_ (.Y(_3214_),
    .A(net298));
 sg13g2_inv_1 _3862_ (.Y(_3215_),
    .A(_0020_));
 sg13g2_inv_1 _3863_ (.Y(_3216_),
    .A(net397));
 sg13g2_inv_1 _3864_ (.Y(_3217_),
    .A(net282));
 sg13g2_inv_1 _3865_ (.Y(_3218_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ));
 sg13g2_inv_1 _3866_ (.Y(_3219_),
    .A(net567));
 sg13g2_inv_1 _3867_ (.Y(_3220_),
    .A(net509));
 sg13g2_inv_1 _3868_ (.Y(_3221_),
    .A(net445));
 sg13g2_inv_1 _3869_ (.Y(_3222_),
    .A(\vgademo.soundtrack.pulse_vol[0] ));
 sg13g2_inv_2 _3870_ (.Y(_3223_),
    .A(net1101));
 sg13g2_inv_2 _3871_ (.Y(_3224_),
    .A(net1114));
 sg13g2_inv_1 _3872_ (.Y(_3225_),
    .A(net1107));
 sg13g2_inv_2 _3873_ (.Y(_3226_),
    .A(net1111));
 sg13g2_inv_1 _3874_ (.Y(_3227_),
    .A(net307));
 sg13g2_inv_1 _3875_ (.Y(_3228_),
    .A(\vgademo.b_sin[8] ));
 sg13g2_inv_1 _3876_ (.Y(_3229_),
    .A(\vgademo.b_sin[9] ));
 sg13g2_inv_1 _3877_ (.Y(_3230_),
    .A(\vgademo.b_sin[10] ));
 sg13g2_inv_1 _3878_ (.Y(_3231_),
    .A(net515));
 sg13g2_inv_2 _3879_ (.Y(_3232_),
    .A(net1051));
 sg13g2_inv_1 _3880_ (.Y(_3233_),
    .A(net496));
 sg13g2_inv_2 _3881_ (.Y(_3234_),
    .A(net469));
 sg13g2_inv_1 _3882_ (.Y(_3235_),
    .A(\vgademo.b_cos[7] ));
 sg13g2_inv_1 _3883_ (.Y(_3236_),
    .A(net461));
 sg13g2_inv_2 _3884_ (.Y(_3237_),
    .A(\vgademo.b_cos[8] ));
 sg13g2_inv_2 _3885_ (.Y(_3238_),
    .A(net1055));
 sg13g2_inv_1 _3886_ (.Y(_3239_),
    .A(net1054));
 sg13g2_inv_1 _3887_ (.Y(_3240_),
    .A(net324));
 sg13g2_inv_1 _3888_ (.Y(_3241_),
    .A(net311));
 sg13g2_inv_1 _3889_ (.Y(_3242_),
    .A(net553));
 sg13g2_inv_1 _3890_ (.Y(_3243_),
    .A(\vgademo.a_sin[11] ));
 sg13g2_inv_1 _3891_ (.Y(_3244_),
    .A(net497));
 sg13g2_inv_1 _3892_ (.Y(_3245_),
    .A(net1057));
 sg13g2_inv_1 _3893_ (.Y(_3246_),
    .A(net354));
 sg13g2_inv_2 _3894_ (.Y(_3247_),
    .A(net472));
 sg13g2_inv_1 _3895_ (.Y(_3248_),
    .A(\vgademo.plane_du[4] ));
 sg13g2_inv_1 _3896_ (.Y(_3249_),
    .A(net420));
 sg13g2_inv_2 _3897_ (.Y(_3250_),
    .A(net545));
 sg13g2_inv_1 _3898_ (.Y(_3251_),
    .A(_0022_));
 sg13g2_inv_1 _3899_ (.Y(_3252_),
    .A(net297));
 sg13g2_inv_1 _3900_ (.Y(_3253_),
    .A(net365));
 sg13g2_inv_1 _3901_ (.Y(_3254_),
    .A(\vgademo.plane_du[7] ));
 sg13g2_inv_1 _3902_ (.Y(_3255_),
    .A(net396));
 sg13g2_inv_2 _3903_ (.Y(_3256_),
    .A(\vgademo.plane_du[8] ));
 sg13g2_inv_1 _3904_ (.Y(_3257_),
    .A(_0025_));
 sg13g2_inv_1 _3905_ (.Y(_3258_),
    .A(net446));
 sg13g2_inv_2 _3906_ (.Y(_3259_),
    .A(\vgademo.plane_du[9] ));
 sg13g2_inv_1 _3907_ (.Y(_3260_),
    .A(net374));
 sg13g2_inv_1 _3908_ (.Y(_3261_),
    .A(net342));
 sg13g2_inv_1 _3909_ (.Y(_3262_),
    .A(net482));
 sg13g2_inv_1 _3910_ (.Y(_3263_),
    .A(net502));
 sg13g2_inv_1 _3911_ (.Y(_3264_),
    .A(net508));
 sg13g2_inv_1 _3912_ (.Y(_3265_),
    .A(net414));
 sg13g2_inv_1 _3913_ (.Y(_3266_),
    .A(net266));
 sg13g2_inv_2 _3914_ (.Y(_3267_),
    .A(net303));
 sg13g2_inv_1 _3915_ (.Y(_3268_),
    .A(\vgademo.linelfsr[5] ));
 sg13g2_inv_1 _3916_ (.Y(_3269_),
    .A(\vgademo.soundtrack.pulse_osc_p[13] ));
 sg13g2_inv_1 _3917_ (.Y(_3270_),
    .A(net366));
 sg13g2_inv_1 _3918_ (.Y(_3271_),
    .A(net398));
 sg13g2_inv_1 _3919_ (.Y(_3272_),
    .A(net448));
 sg13g2_inv_1 _3920_ (.Y(_3273_),
    .A(net538));
 sg13g2_inv_1 _3921_ (.Y(_3274_),
    .A(net527));
 sg13g2_inv_1 _3922_ (.Y(_3275_),
    .A(net218));
 sg13g2_inv_1 _3923_ (.Y(_3276_),
    .A(net361));
 sg13g2_inv_1 _3924_ (.Y(_3277_),
    .A(net323));
 sg13g2_inv_1 _3925_ (.Y(_3278_),
    .A(net372));
 sg13g2_inv_1 _3926_ (.Y(_3279_),
    .A(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_inv_1 _3927_ (.Y(_3280_),
    .A(net350));
 sg13g2_inv_1 _3928_ (.Y(_3281_),
    .A(net563));
 sg13g2_inv_1 _3929_ (.Y(_3282_),
    .A(net312));
 sg13g2_nand2_2 _3930_ (.Y(_3283_),
    .A(\vgademo.h_count[7] ),
    .B(\vgademo.h_count[6] ));
 sg13g2_nor3_2 _3931_ (.A(_3192_),
    .B(_3193_),
    .C(_3283_),
    .Y(_3284_));
 sg13g2_nor4_2 _3932_ (.A(net1096),
    .B(net1098),
    .C(net1094),
    .Y(_3285_),
    .D(_3191_));
 sg13g2_inv_1 _3933_ (.Y(_3286_),
    .A(_3285_));
 sg13g2_nor2_1 _3934_ (.A(\vgademo.h_count[9] ),
    .B(_0060_),
    .Y(_3287_));
 sg13g2_and4_1 _3935_ (.A(\vgademo.h_count[8] ),
    .B(_3284_),
    .C(_3285_),
    .D(_3287_),
    .X(_3288_));
 sg13g2_nand4_1 _3936_ (.B(_3284_),
    .C(_3285_),
    .A(\vgademo.h_count[8] ),
    .Y(_3289_),
    .D(_3287_));
 sg13g2_nor2_1 _3937_ (.A(net166),
    .B(net1035),
    .Y(_0000_));
 sg13g2_nand2_2 _3938_ (.Y(_3290_),
    .A(net1097),
    .B(net1098));
 sg13g2_xor2_1 _3939_ (.B(net1098),
    .A(net1097),
    .X(_0002_));
 sg13g2_and2_1 _3940_ (.A(net536),
    .B(_3290_),
    .X(_3291_));
 sg13g2_nor2_1 _3941_ (.A(net536),
    .B(_3290_),
    .Y(_3292_));
 sg13g2_nor3_1 _3942_ (.A(net1035),
    .B(_3291_),
    .C(_3292_),
    .Y(_0003_));
 sg13g2_xor2_1 _3943_ (.B(_3292_),
    .A(net321),
    .X(_3293_));
 sg13g2_nor2_1 _3944_ (.A(net1035),
    .B(net322),
    .Y(_0004_));
 sg13g2_nor3_2 _3945_ (.A(_3190_),
    .B(_3191_),
    .C(_3290_),
    .Y(_3294_));
 sg13g2_nand2_1 _3946_ (.Y(_3295_),
    .A(\vgademo.h_count[4] ),
    .B(_3294_));
 sg13g2_o21ai_1 _3947_ (.B1(net1033),
    .Y(_3296_),
    .A1(net417),
    .A2(_3294_));
 sg13g2_nor2b_1 _3948_ (.A(_3296_),
    .B_N(_3295_),
    .Y(_0005_));
 sg13g2_o21ai_1 _3949_ (.B1(net1033),
    .Y(_3297_),
    .A1(net300),
    .A2(_3295_));
 sg13g2_a21oi_1 _3950_ (.A1(net300),
    .A2(_3295_),
    .Y(_0006_),
    .B1(_3297_));
 sg13g2_nand3_1 _3951_ (.B(\vgademo.h_count[4] ),
    .C(_3294_),
    .A(\vgademo.h_count[5] ),
    .Y(_3298_));
 sg13g2_nor2_1 _3952_ (.A(net575),
    .B(_3298_),
    .Y(_3299_));
 sg13g2_a21oi_1 _3953_ (.A1(net575),
    .A2(_3298_),
    .Y(_3300_),
    .B1(net1035));
 sg13g2_nor2b_1 _3954_ (.A(_3299_),
    .B_N(_3300_),
    .Y(_0007_));
 sg13g2_nor3_1 _3955_ (.A(_0035_),
    .B(net558),
    .C(_3298_),
    .Y(_3301_));
 sg13g2_nor2b_1 _3956_ (.A(_3299_),
    .B_N(net558),
    .Y(_3302_));
 sg13g2_nor3_1 _3957_ (.A(net1035),
    .B(_3301_),
    .C(net559),
    .Y(_0008_));
 sg13g2_or2_1 _3958_ (.X(_3303_),
    .B(_3298_),
    .A(_3283_));
 sg13g2_nor2_1 _3959_ (.A(net562),
    .B(_3303_),
    .Y(_3304_));
 sg13g2_a21oi_1 _3960_ (.A1(net562),
    .A2(_3303_),
    .Y(_3305_),
    .B1(net1035));
 sg13g2_nor2b_1 _3961_ (.A(_3304_),
    .B_N(_3305_),
    .Y(_0009_));
 sg13g2_nor3_1 _3962_ (.A(_0037_),
    .B(net385),
    .C(_3303_),
    .Y(_3306_));
 sg13g2_nor2b_1 _3963_ (.A(_3304_),
    .B_N(net385),
    .Y(_3307_));
 sg13g2_nor3_1 _3964_ (.A(net1035),
    .B(_3306_),
    .C(net386),
    .Y(_0010_));
 sg13g2_nand2_1 _3965_ (.Y(_3308_),
    .A(\vgademo.h_count[9] ),
    .B(\vgademo.h_count[8] ));
 sg13g2_or2_1 _3966_ (.X(_3309_),
    .B(_3308_),
    .A(_3303_));
 sg13g2_a21oi_1 _3967_ (.A1(net1092),
    .A2(_3309_),
    .Y(_3310_),
    .B1(net1035));
 sg13g2_o21ai_1 _3968_ (.B1(_3310_),
    .Y(_3311_),
    .A1(net1092),
    .A2(_3309_));
 sg13g2_inv_1 _3969_ (.Y(_0001_),
    .A(_3311_));
 sg13g2_nor2_2 _3970_ (.A(\vgademo.v_count[8] ),
    .B(net1059),
    .Y(_3312_));
 sg13g2_nand2_1 _3971_ (.Y(_3313_),
    .A(\vgademo.v_count[7] ),
    .B(net1061));
 sg13g2_nor3_2 _3972_ (.A(_0062_),
    .B(_3312_),
    .C(_3313_),
    .Y(_3314_));
 sg13g2_nand2b_1 _3973_ (.Y(_3315_),
    .B(\vgademo.v_count[8] ),
    .A_N(\vgademo.v_count[9] ));
 sg13g2_or4_1 _3974_ (.A(net1062),
    .B(_3185_),
    .C(_3313_),
    .D(_3315_),
    .X(_3316_));
 sg13g2_nand2_1 _3975_ (.Y(_3317_),
    .A(net476),
    .B(net1064));
 sg13g2_nor3_1 _3976_ (.A(net1065),
    .B(_3316_),
    .C(_3317_),
    .Y(_3318_));
 sg13g2_o21ai_1 _3977_ (.B1(_3318_),
    .Y(_0012_),
    .A1(_3184_),
    .A2(_3314_));
 sg13g2_nor2_2 _3978_ (.A(\vgademo.h_count[9] ),
    .B(\vgademo.h_count[8] ),
    .Y(_3319_));
 sg13g2_nand2b_1 _3979_ (.Y(_3320_),
    .B(_3319_),
    .A_N(_3284_));
 sg13g2_nand3_1 _3980_ (.B(_3191_),
    .C(_3290_),
    .A(_3190_),
    .Y(_3321_));
 sg13g2_nor3_1 _3981_ (.A(_3192_),
    .B(\vgademo.h_count[4] ),
    .C(_3283_),
    .Y(_3322_));
 sg13g2_a22oi_1 _3982_ (.Y(_3323_),
    .B1(_3321_),
    .B2(_3322_),
    .A2(_3320_),
    .A1(\vgademo.h_count[10] ));
 sg13g2_nor2_1 _3983_ (.A(net1096),
    .B(net1095),
    .Y(_3324_));
 sg13g2_nand2_1 _3984_ (.Y(_3325_),
    .A(net1094),
    .B(\vgademo.h_count[4] ));
 sg13g2_nor2_1 _3985_ (.A(\vgademo.h_count[5] ),
    .B(\vgademo.h_count[6] ),
    .Y(_3326_));
 sg13g2_o21ai_1 _3986_ (.B1(_3326_),
    .Y(_3327_),
    .A1(_3324_),
    .A2(_3325_));
 sg13g2_nand3_1 _3987_ (.B(\vgademo.h_count[8] ),
    .C(_3327_),
    .A(\vgademo.h_count[7] ),
    .Y(_3328_));
 sg13g2_nor2b_1 _3988_ (.A(\vgademo.h_count[9] ),
    .B_N(\vgademo.h_count[10] ),
    .Y(_3329_));
 sg13g2_nor3_2 _3989_ (.A(\vgademo.h_count[9] ),
    .B(\vgademo.h_count[8] ),
    .C(net1092),
    .Y(_3330_));
 sg13g2_nor3_1 _3990_ (.A(net1094),
    .B(net1095),
    .C(\vgademo.h_count[10] ),
    .Y(_3331_));
 sg13g2_a22oi_1 _3991_ (.Y(_3332_),
    .B1(_3330_),
    .B2(_3331_),
    .A2(_3329_),
    .A1(_3328_));
 sg13g2_or2_2 _3992_ (.X(_0011_),
    .B(_3332_),
    .A(_3323_));
 sg13g2_nand2b_1 _3993_ (.Y(_3333_),
    .B(net1103),
    .A_N(net1104));
 sg13g2_nor2_1 _3994_ (.A(_3181_),
    .B(net1131),
    .Y(_3334_));
 sg13g2_nand2b_2 _3995_ (.Y(_3335_),
    .B(net1132),
    .A_N(net1131));
 sg13g2_nor2_2 _3996_ (.A(net1139),
    .B(net1134),
    .Y(_3336_));
 sg13g2_nand2_2 _3997_ (.Y(_3337_),
    .A(_3177_),
    .B(net1047));
 sg13g2_or2_1 _3998_ (.X(_3338_),
    .B(net1145),
    .A(net1147));
 sg13g2_nand2_1 _3999_ (.Y(_3339_),
    .A(net1147),
    .B(net1140));
 sg13g2_nand2_2 _4000_ (.Y(_3340_),
    .A(net1140),
    .B(net1144));
 sg13g2_nand2_1 _4001_ (.Y(_3341_),
    .A(_3339_),
    .B(_3340_));
 sg13g2_nand3_1 _4002_ (.B(_3339_),
    .C(_3340_),
    .A(_3336_),
    .Y(_3342_));
 sg13g2_nor2_2 _4003_ (.A(net1140),
    .B(net1144),
    .Y(_3343_));
 sg13g2_nor2_1 _4004_ (.A(net1137),
    .B(_3343_),
    .Y(_3344_));
 sg13g2_nor2b_2 _4005_ (.A(net1134),
    .B_N(net1139),
    .Y(_3345_));
 sg13g2_nor2_1 _4006_ (.A(\vgademo.audio_songpos[1] ),
    .B(net1049),
    .Y(_3346_));
 sg13g2_nand2b_2 _4007_ (.Y(_3347_),
    .B(net1140),
    .A_N(net1147));
 sg13g2_nand2_1 _4008_ (.Y(_3348_),
    .A(_3345_),
    .B(_3347_));
 sg13g2_nor2_2 _4009_ (.A(net1150),
    .B(net1147),
    .Y(_3349_));
 sg13g2_nand2b_1 _4010_ (.Y(_3350_),
    .B(net1151),
    .A_N(net1145));
 sg13g2_a21oi_1 _4011_ (.A1(_3345_),
    .A2(_3350_),
    .Y(_3351_),
    .B1(_3349_));
 sg13g2_nor2_1 _4012_ (.A(net1144),
    .B(_3347_),
    .Y(_3352_));
 sg13g2_nand3b_1 _4013_ (.B(_3348_),
    .C(_3351_),
    .Y(_3353_),
    .A_N(_3344_));
 sg13g2_nand2_1 _4014_ (.Y(_3354_),
    .A(_3342_),
    .B(_3353_));
 sg13g2_a21oi_1 _4015_ (.A1(_3342_),
    .A2(_3353_),
    .Y(_3355_),
    .B1(_3335_));
 sg13g2_nor2b_1 _4016_ (.A(net1150),
    .B_N(net1147),
    .Y(_3356_));
 sg13g2_nor2_1 _4017_ (.A(_3170_),
    .B(net1048),
    .Y(_3357_));
 sg13g2_and2_1 _4018_ (.A(net1148),
    .B(net1145),
    .X(_3358_));
 sg13g2_nand2_2 _4019_ (.Y(_3359_),
    .A(\vgademo.audio_songpos[1] ),
    .B(net1145));
 sg13g2_nand2_1 _4020_ (.Y(_3360_),
    .A(net1141),
    .B(_3359_));
 sg13g2_o21ai_1 _4021_ (.B1(net1141),
    .Y(_3361_),
    .A1(net1150),
    .A2(_3359_));
 sg13g2_and2_1 _4022_ (.A(net1151),
    .B(net1149),
    .X(_3362_));
 sg13g2_nand2_1 _4023_ (.Y(_3363_),
    .A(net1150),
    .B(net1148));
 sg13g2_xor2_1 _4024_ (.B(net1149),
    .A(net1151),
    .X(_3364_));
 sg13g2_xnor2_1 _4025_ (.Y(_3365_),
    .A(net1150),
    .B(net1149));
 sg13g2_nor2b_2 _4026_ (.A(net1149),
    .B_N(net1151),
    .Y(_3366_));
 sg13g2_a221oi_1 _4027_ (.B2(_3179_),
    .C1(net1048),
    .B1(_3365_),
    .A1(_3170_),
    .Y(_3367_),
    .A2(_3358_));
 sg13g2_and2_1 _4028_ (.A(_3343_),
    .B(_3365_),
    .X(_3368_));
 sg13g2_o21ai_1 _4029_ (.B1(net1139),
    .Y(_3369_),
    .A1(_3367_),
    .A2(_3368_));
 sg13g2_o21ai_1 _4030_ (.B1(net1048),
    .Y(_3370_),
    .A1(_3179_),
    .A2(_3364_));
 sg13g2_nand3_1 _4031_ (.B(_3338_),
    .C(_3350_),
    .A(_3177_),
    .Y(_3371_));
 sg13g2_a21o_1 _4032_ (.A2(_3370_),
    .A1(_3361_),
    .B1(_3371_),
    .X(_3372_));
 sg13g2_nand3_1 _4033_ (.B(_3369_),
    .C(_3372_),
    .A(net1135),
    .Y(_3373_));
 sg13g2_nor2b_1 _4034_ (.A(net1143),
    .B_N(net1149),
    .Y(_3374_));
 sg13g2_nor2_1 _4035_ (.A(net1150),
    .B(net1145),
    .Y(_3375_));
 sg13g2_nor3_1 _4036_ (.A(_3366_),
    .B(_3374_),
    .C(_3375_),
    .Y(_3376_));
 sg13g2_o21ai_1 _4037_ (.B1(_3336_),
    .Y(_3377_),
    .A1(_3343_),
    .A2(_3376_));
 sg13g2_nor2b_2 _4038_ (.A(net1144),
    .B_N(net1148),
    .Y(_3378_));
 sg13g2_nand2b_2 _4039_ (.Y(_3379_),
    .B(net1147),
    .A_N(net1144));
 sg13g2_o21ai_1 _4040_ (.B1(_3356_),
    .Y(_3380_),
    .A1(net1048),
    .A2(_3379_));
 sg13g2_nand3_1 _4041_ (.B(net1140),
    .C(_3378_),
    .A(net1150),
    .Y(_3381_));
 sg13g2_nand3_1 _4042_ (.B(_3380_),
    .C(_3381_),
    .A(_3345_),
    .Y(_3382_));
 sg13g2_nand2_2 _4043_ (.Y(_3383_),
    .A(net1132),
    .B(\vgademo.audio_songpos[7] ));
 sg13g2_and4_1 _4044_ (.A(net1133),
    .B(net1131),
    .C(_3377_),
    .D(_3382_),
    .X(_3384_));
 sg13g2_a21o_1 _4045_ (.A2(_3384_),
    .A1(_3373_),
    .B1(_3355_),
    .X(_3385_));
 sg13g2_a221oi_1 _4046_ (.B2(_3384_),
    .C1(_3269_),
    .B1(_3373_),
    .A1(_3334_),
    .Y(_3386_),
    .A2(_3354_));
 sg13g2_a21o_2 _4047_ (.A2(_3385_),
    .A1(\vgademo.soundtrack.pulse_osc_p[12] ),
    .B1(_3386_),
    .X(_3387_));
 sg13g2_a21oi_1 _4048_ (.A1(\vgademo.soundtrack.pulse_osc_p[12] ),
    .A2(_3385_),
    .Y(_3388_),
    .B1(_3386_));
 sg13g2_nor2_2 _4049_ (.A(_3222_),
    .B(_3387_),
    .Y(_3389_));
 sg13g2_a21oi_2 _4050_ (.B1(_3333_),
    .Y(_3390_),
    .A2(_3388_),
    .A1(\vgademo.soundtrack.pulse_vol[0] ));
 sg13g2_mux2_1 _4051_ (.A0(\vgademo.soundtrack.noise_lfsr[10] ),
    .A1(\vgademo.soundtrack.noise_lfsr[11] ),
    .S(net1116),
    .X(_3391_));
 sg13g2_nand2_1 _4052_ (.Y(_3392_),
    .A(net1112),
    .B(_3391_));
 sg13g2_nand2b_1 _4053_ (.Y(_3393_),
    .B(net1117),
    .A_N(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_o21ai_1 _4054_ (.B1(_3393_),
    .Y(_3394_),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .A2(net1117));
 sg13g2_o21ai_1 _4055_ (.B1(_3392_),
    .Y(_3395_),
    .A1(net1112),
    .A2(_3394_));
 sg13g2_nor2_1 _4056_ (.A(net1108),
    .B(_3395_),
    .Y(_3396_));
 sg13g2_nand3b_1 _4057_ (.B(\vgademo.soundtrack.noise_lfsr[12] ),
    .C(net1043),
    .Y(_3397_),
    .A_N(net1116));
 sg13g2_a21oi_1 _4058_ (.A1(net1108),
    .A2(_3397_),
    .Y(_3398_),
    .B1(_3396_));
 sg13g2_nor2_1 _4059_ (.A(net1117),
    .B(_0039_),
    .Y(_3399_));
 sg13g2_a21oi_1 _4060_ (.A1(net1117),
    .A2(\vgademo.soundtrack.noise_lfsr[5] ),
    .Y(_3400_),
    .B1(_3399_));
 sg13g2_nor2_1 _4061_ (.A(net1112),
    .B(_3400_),
    .Y(_3401_));
 sg13g2_mux2_1 _4062_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(\vgademo.soundtrack.noise_lfsr[7] ),
    .S(net1117),
    .X(_3402_));
 sg13g2_a21oi_1 _4063_ (.A1(net1112),
    .A2(_3402_),
    .Y(_3403_),
    .B1(_3401_));
 sg13g2_nor2_1 _4064_ (.A(\vgademo.soundtrack.noise_lfsr[2] ),
    .B(net1115),
    .Y(_3404_));
 sg13g2_nor2b_1 _4065_ (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .B_N(net1115),
    .Y(_3405_));
 sg13g2_mux4_1 _4066_ (.S0(net1115),
    .A0(\vgademo.soundtrack.noise_lfsr[0] ),
    .A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(\vgademo.soundtrack.noise_lfsr[2] ),
    .A3(\vgademo.soundtrack.noise_lfsr[3] ),
    .S1(net1113),
    .X(_3406_));
 sg13g2_nand2_1 _4067_ (.Y(_3407_),
    .A(net1105),
    .B(_3398_));
 sg13g2_a21oi_1 _4068_ (.A1(net1109),
    .A2(_3403_),
    .Y(_3408_),
    .B1(net1106));
 sg13g2_o21ai_1 _4069_ (.B1(_3408_),
    .Y(_3409_),
    .A1(net1109),
    .A2(_3406_));
 sg13g2_nand2_1 _4070_ (.Y(_3410_),
    .A(_3407_),
    .B(_3409_));
 sg13g2_nand3_1 _4071_ (.B(_3390_),
    .C(_3410_),
    .A(net1101),
    .Y(_3411_));
 sg13g2_a21oi_1 _4072_ (.A1(net1101),
    .A2(_3390_),
    .Y(_3412_),
    .B1(_3410_));
 sg13g2_a21o_1 _4073_ (.A2(_3390_),
    .A1(net1101),
    .B1(_3410_),
    .X(_3413_));
 sg13g2_and2_1 _4074_ (.A(_3411_),
    .B(_3413_),
    .X(_3414_));
 sg13g2_xnor2_1 _4075_ (.Y(_3415_),
    .A(net1100),
    .B(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_xnor2_1 _4076_ (.Y(_3416_),
    .A(_3414_),
    .B(_3415_));
 sg13g2_and2_1 _4077_ (.A(net214),
    .B(_3416_),
    .X(_3417_));
 sg13g2_xor2_1 _4078_ (.B(_3416_),
    .A(net214),
    .X(\vgademo.soundtrack.sigma_delta_accum_[0] ));
 sg13g2_o21ai_1 _4079_ (.B1(_3411_),
    .Y(_3418_),
    .A1(_3412_),
    .A2(_3415_));
 sg13g2_nand2_2 _4080_ (.Y(_3419_),
    .A(net1104),
    .B(net1103));
 sg13g2_nor2_2 _4081_ (.A(_3223_),
    .B(_3419_),
    .Y(_3420_));
 sg13g2_xnor2_1 _4082_ (.Y(_3421_),
    .A(_3223_),
    .B(_3419_));
 sg13g2_xnor2_1 _4083_ (.Y(_3422_),
    .A(net1104),
    .B(net1103));
 sg13g2_inv_1 _4084_ (.Y(_3423_),
    .A(_3422_));
 sg13g2_and2_1 _4085_ (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .B(\vgademo.soundtrack.pulse_vol[0] ),
    .X(_3424_));
 sg13g2_nor2_1 _4086_ (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .B(\vgademo.soundtrack.pulse_vol[0] ),
    .Y(_3425_));
 sg13g2_nor2_1 _4087_ (.A(_3424_),
    .B(_3425_),
    .Y(_3426_));
 sg13g2_a221oi_1 _4088_ (.B2(_3385_),
    .C1(_3386_),
    .B1(\vgademo.soundtrack.pulse_osc_p[12] ),
    .A1(net1104),
    .Y(_3427_),
    .A2(\vgademo.soundtrack.pulse_vol[0] ));
 sg13g2_or2_2 _4089_ (.X(_3428_),
    .B(_3427_),
    .A(_3426_));
 sg13g2_nor4_1 _4090_ (.A(_3421_),
    .B(_3422_),
    .C(_3426_),
    .D(_3427_),
    .Y(_3429_));
 sg13g2_mux2_1 _4091_ (.A0(\vgademo.soundtrack.noise_lfsr[7] ),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .S(net1117),
    .X(_3430_));
 sg13g2_mux2_1 _4092_ (.A0(\vgademo.soundtrack.noise_lfsr[5] ),
    .A1(\vgademo.soundtrack.noise_lfsr[6] ),
    .S(net1117),
    .X(_3431_));
 sg13g2_mux2_1 _4093_ (.A0(_3430_),
    .A1(_3431_),
    .S(net1043),
    .X(_3432_));
 sg13g2_inv_1 _4094_ (.Y(_3433_),
    .A(_3432_));
 sg13g2_nor2_1 _4095_ (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .B(net1115),
    .Y(_3434_));
 sg13g2_a21oi_1 _4096_ (.A1(net1115),
    .A2(_0039_),
    .Y(_3435_),
    .B1(_3434_));
 sg13g2_nand2b_1 _4097_ (.Y(_3436_),
    .B(net1115),
    .A_N(\vgademo.soundtrack.noise_lfsr[2] ));
 sg13g2_o21ai_1 _4098_ (.B1(_3436_),
    .Y(_3437_),
    .A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(net1115));
 sg13g2_nor2b_1 _4099_ (.A(net1116),
    .B_N(\vgademo.soundtrack.noise_lfsr[9] ),
    .Y(_3438_));
 sg13g2_a21oi_1 _4100_ (.A1(net1116),
    .A2(\vgademo.soundtrack.noise_lfsr[10] ),
    .Y(_3439_),
    .B1(_3438_));
 sg13g2_mux2_1 _4101_ (.A0(\vgademo.soundtrack.noise_lfsr[11] ),
    .A1(\vgademo.soundtrack.noise_lfsr[12] ),
    .S(net1115),
    .X(_3440_));
 sg13g2_nor2_1 _4102_ (.A(net1043),
    .B(_3440_),
    .Y(_3441_));
 sg13g2_a21oi_1 _4103_ (.A1(net1043),
    .A2(_3439_),
    .Y(_3442_),
    .B1(_3441_));
 sg13g2_and2_1 _4104_ (.A(_3226_),
    .B(_3442_),
    .X(_3443_));
 sg13g2_a21oi_1 _4105_ (.A1(net1112),
    .A2(_3435_),
    .Y(_3444_),
    .B1(net1109));
 sg13g2_o21ai_1 _4106_ (.B1(_3444_),
    .Y(_3445_),
    .A1(net1112),
    .A2(_3437_));
 sg13g2_a21oi_1 _4107_ (.A1(net1110),
    .A2(_3433_),
    .Y(_3446_),
    .B1(net1105));
 sg13g2_a22oi_1 _4108_ (.Y(_3447_),
    .B1(_3445_),
    .B2(_3446_),
    .A2(_3443_),
    .A1(net1105));
 sg13g2_or4_1 _4109_ (.A(_3421_),
    .B(_3422_),
    .C(_3428_),
    .D(_3447_),
    .X(_3448_));
 sg13g2_xor2_1 _4110_ (.B(_3447_),
    .A(_3429_),
    .X(_3449_));
 sg13g2_xnor2_1 _4111_ (.Y(_3450_),
    .A(net1099),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_xnor2_1 _4112_ (.Y(_3451_),
    .A(_3449_),
    .B(_3450_));
 sg13g2_nand2b_1 _4113_ (.Y(_3452_),
    .B(_3418_),
    .A_N(_3451_));
 sg13g2_xor2_1 _4114_ (.B(_3451_),
    .A(_3418_),
    .X(_3453_));
 sg13g2_nor2_1 _4115_ (.A(_3273_),
    .B(_3453_),
    .Y(_3454_));
 sg13g2_nand2_1 _4116_ (.Y(_3455_),
    .A(_3273_),
    .B(_3453_));
 sg13g2_nand2b_1 _4117_ (.Y(_3456_),
    .B(_3455_),
    .A_N(_3454_));
 sg13g2_xnor2_1 _4118_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[1] ),
    .A(_3417_),
    .B(_3456_));
 sg13g2_a21oi_1 _4119_ (.A1(_3417_),
    .A2(_3455_),
    .Y(_3457_),
    .B1(_3454_));
 sg13g2_o21ai_1 _4120_ (.B1(_3448_),
    .Y(_3458_),
    .A1(_3449_),
    .A2(_3450_));
 sg13g2_nor2b_1 _4121_ (.A(net1103),
    .B_N(net1104),
    .Y(_3459_));
 sg13g2_o21ai_1 _4122_ (.B1(_3459_),
    .Y(_3460_),
    .A1(_3222_),
    .A2(_3387_));
 sg13g2_nand2_1 _4123_ (.Y(_3461_),
    .A(net1044),
    .B(_3402_));
 sg13g2_o21ai_1 _4124_ (.B1(_3461_),
    .Y(_3462_),
    .A1(net1044),
    .A2(_3394_));
 sg13g2_o21ai_1 _4125_ (.B1(net1044),
    .Y(_3463_),
    .A1(_3404_),
    .A2(_3405_));
 sg13g2_a21oi_1 _4126_ (.A1(net1112),
    .A2(_3400_),
    .Y(_3464_),
    .B1(net1109));
 sg13g2_a221oi_1 _4127_ (.B2(_3464_),
    .C1(net1106),
    .B1(_3463_),
    .A1(net1109),
    .Y(_3465_),
    .A2(_3462_));
 sg13g2_nor2_1 _4128_ (.A(net1043),
    .B(net1116),
    .Y(_3466_));
 sg13g2_a22oi_1 _4129_ (.Y(_3467_),
    .B1(_3466_),
    .B2(\vgademo.soundtrack.noise_lfsr[12] ),
    .A2(_3391_),
    .A1(net1043));
 sg13g2_or2_1 _4130_ (.X(_3468_),
    .B(_3467_),
    .A(net1108));
 sg13g2_a21o_1 _4131_ (.A2(_3468_),
    .A1(net1105),
    .B1(_3465_),
    .X(_0365_));
 sg13g2_or3_1 _4132_ (.A(_3223_),
    .B(_3460_),
    .C(_0365_),
    .X(_0366_));
 sg13g2_o21ai_1 _4133_ (.B1(_0365_),
    .Y(_0367_),
    .A1(_3223_),
    .A2(_3460_));
 sg13g2_xor2_1 _4134_ (.B(\vgademo.soundtrack.tri_osc_p[3] ),
    .A(net1099),
    .X(_0368_));
 sg13g2_nand3_1 _4135_ (.B(_0367_),
    .C(_0368_),
    .A(_0366_),
    .Y(_0369_));
 sg13g2_a21o_1 _4136_ (.A2(_0367_),
    .A1(_0366_),
    .B1(_0368_),
    .X(_0370_));
 sg13g2_and3_1 _4137_ (.X(_0371_),
    .A(_3458_),
    .B(_0369_),
    .C(_0370_));
 sg13g2_nand3_1 _4138_ (.B(_0369_),
    .C(_0370_),
    .A(_3458_),
    .Y(_0372_));
 sg13g2_a21oi_1 _4139_ (.A1(_0369_),
    .A2(_0370_),
    .Y(_0373_),
    .B1(_3458_));
 sg13g2_or3_1 _4140_ (.A(_3452_),
    .B(_0371_),
    .C(_0373_),
    .X(_0374_));
 sg13g2_o21ai_1 _4141_ (.B1(_3452_),
    .Y(_0375_),
    .A1(_0371_),
    .A2(_0373_));
 sg13g2_and3_1 _4142_ (.X(_0376_),
    .A(net549),
    .B(_0374_),
    .C(_0375_));
 sg13g2_nand3_1 _4143_ (.B(_0374_),
    .C(_0375_),
    .A(\vgademo.soundtrack.sigma_delta_accum[2] ),
    .Y(_0377_));
 sg13g2_a21oi_1 _4144_ (.A1(_0374_),
    .A2(_0375_),
    .Y(_0378_),
    .B1(net549));
 sg13g2_nor2_1 _4145_ (.A(_0376_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_xnor2_1 _4146_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .A(_3457_),
    .B(_0379_));
 sg13g2_o21ai_1 _4147_ (.B1(_0377_),
    .Y(_0380_),
    .A1(_3457_),
    .A2(_0378_));
 sg13g2_o21ai_1 _4148_ (.B1(_0372_),
    .Y(_0381_),
    .A1(_3452_),
    .A2(_0373_));
 sg13g2_nand2_1 _4149_ (.Y(_0382_),
    .A(_0366_),
    .B(_0369_));
 sg13g2_nor3_1 _4150_ (.A(net1103),
    .B(_3424_),
    .C(_3425_),
    .Y(_0383_));
 sg13g2_o21ai_1 _4151_ (.B1(_0383_),
    .Y(_0384_),
    .A1(\vgademo.soundtrack.pulse_vol[0] ),
    .A2(_3387_));
 sg13g2_nor2_1 _4152_ (.A(_3421_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_nor2_1 _4153_ (.A(net1113),
    .B(_3430_),
    .Y(_0386_));
 sg13g2_a21oi_1 _4154_ (.A1(net1113),
    .A2(_3439_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_nand2_1 _4155_ (.Y(_0388_),
    .A(net1112),
    .B(_3431_));
 sg13g2_a21oi_1 _4156_ (.A1(net1043),
    .A2(_3435_),
    .Y(_0389_),
    .B1(net1108));
 sg13g2_o21ai_1 _4157_ (.B1(net1042),
    .Y(_0390_),
    .A1(_3226_),
    .A2(_0387_));
 sg13g2_a21oi_1 _4158_ (.A1(_0388_),
    .A2(_0389_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_nand2_1 _4159_ (.Y(_0392_),
    .A(net1043),
    .B(_3440_));
 sg13g2_nor2_1 _4160_ (.A(net1110),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_a21oi_2 _4161_ (.B1(_0391_),
    .Y(_0394_),
    .A2(_0393_),
    .A1(net1105));
 sg13g2_nor3_1 _4162_ (.A(_3421_),
    .B(_0384_),
    .C(_0394_),
    .Y(_0395_));
 sg13g2_xnor2_1 _4163_ (.Y(_0396_),
    .A(_0385_),
    .B(_0394_));
 sg13g2_xor2_1 _4164_ (.B(\vgademo.soundtrack.tri_osc_p[4] ),
    .A(net1099),
    .X(_0397_));
 sg13g2_xor2_1 _4165_ (.B(_0397_),
    .A(_0396_),
    .X(_0398_));
 sg13g2_and2_1 _4166_ (.A(_0382_),
    .B(_0398_),
    .X(_0399_));
 sg13g2_or2_1 _4167_ (.X(_0400_),
    .B(_0398_),
    .A(_0382_));
 sg13g2_xor2_1 _4168_ (.B(_0398_),
    .A(_0382_),
    .X(_0401_));
 sg13g2_xnor2_1 _4169_ (.Y(_0402_),
    .A(_0381_),
    .B(_0401_));
 sg13g2_nor2_1 _4170_ (.A(_3274_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_xnor2_1 _4171_ (.Y(_0404_),
    .A(net527),
    .B(_0402_));
 sg13g2_xor2_1 _4172_ (.B(_0404_),
    .A(_0380_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[3] ));
 sg13g2_a21oi_1 _4173_ (.A1(_0380_),
    .A2(_0404_),
    .Y(_0405_),
    .B1(_0403_));
 sg13g2_a21o_1 _4174_ (.A2(_0400_),
    .A1(_0381_),
    .B1(_0399_),
    .X(_0406_));
 sg13g2_a21oi_1 _4175_ (.A1(_0396_),
    .A2(_0397_),
    .Y(_0407_),
    .B1(_0395_));
 sg13g2_or4_1 _4176_ (.A(net1104),
    .B(net1103),
    .C(_3223_),
    .D(_3389_),
    .X(_0408_));
 sg13g2_o21ai_1 _4177_ (.B1(net1105),
    .Y(_0409_),
    .A1(net1108),
    .A2(_3397_));
 sg13g2_a21oi_1 _4178_ (.A1(net1109),
    .A2(_3395_),
    .Y(_0410_),
    .B1(net1105));
 sg13g2_o21ai_1 _4179_ (.B1(_0410_),
    .Y(_0411_),
    .A1(net1108),
    .A2(_3403_));
 sg13g2_nand2_1 _4180_ (.Y(_0412_),
    .A(_0409_),
    .B(_0411_));
 sg13g2_xor2_1 _4181_ (.B(_0412_),
    .A(_0408_),
    .X(_0413_));
 sg13g2_xnor2_1 _4182_ (.Y(_0414_),
    .A(net1099),
    .B(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_nand2b_1 _4183_ (.Y(_0415_),
    .B(_0413_),
    .A_N(_0414_));
 sg13g2_xor2_1 _4184_ (.B(_0414_),
    .A(_0413_),
    .X(_0416_));
 sg13g2_nor2_1 _4185_ (.A(_0407_),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_xor2_1 _4186_ (.B(_0416_),
    .A(_0407_),
    .X(_0418_));
 sg13g2_xor2_1 _4187_ (.B(_0418_),
    .A(_0406_),
    .X(_0419_));
 sg13g2_nand2_1 _4188_ (.Y(_0420_),
    .A(net533),
    .B(_0419_));
 sg13g2_xnor2_1 _4189_ (.Y(_0421_),
    .A(net533),
    .B(_0419_));
 sg13g2_xor2_1 _4190_ (.B(_0421_),
    .A(_0405_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[4] ));
 sg13g2_o21ai_1 _4191_ (.B1(_0420_),
    .Y(_0422_),
    .A1(_0405_),
    .A2(_0421_));
 sg13g2_a21oi_1 _4192_ (.A1(_0406_),
    .A2(_0418_),
    .Y(_0423_),
    .B1(_0417_));
 sg13g2_o21ai_1 _4193_ (.B1(_0415_),
    .Y(_0424_),
    .A1(_0408_),
    .A2(_0412_));
 sg13g2_nor3_2 _4194_ (.A(_3421_),
    .B(_3423_),
    .C(_3428_),
    .Y(_0425_));
 sg13g2_o21ai_1 _4195_ (.B1(net1042),
    .Y(_0426_),
    .A1(_3226_),
    .A2(_3442_));
 sg13g2_a21oi_2 _4196_ (.B1(_0426_),
    .Y(_0427_),
    .A2(_3433_),
    .A1(_3226_));
 sg13g2_nand2_1 _4197_ (.Y(_0428_),
    .A(_0425_),
    .B(_0427_));
 sg13g2_xnor2_1 _4198_ (.Y(_0429_),
    .A(_0425_),
    .B(_0427_));
 sg13g2_xor2_1 _4199_ (.B(\vgademo.soundtrack.tri_osc_p[6] ),
    .A(net1099),
    .X(_0430_));
 sg13g2_inv_1 _4200_ (.Y(_0431_),
    .A(_0430_));
 sg13g2_xnor2_1 _4201_ (.Y(_0432_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_nand2_1 _4202_ (.Y(_0433_),
    .A(_0424_),
    .B(_0432_));
 sg13g2_xnor2_1 _4203_ (.Y(_0434_),
    .A(_0424_),
    .B(_0432_));
 sg13g2_xor2_1 _4204_ (.B(_0434_),
    .A(_0423_),
    .X(_0435_));
 sg13g2_and2_1 _4205_ (.A(net570),
    .B(_0435_),
    .X(_0436_));
 sg13g2_or2_1 _4206_ (.X(_0437_),
    .B(_0435_),
    .A(net570));
 sg13g2_nand2b_1 _4207_ (.Y(_0438_),
    .B(_0437_),
    .A_N(_0436_));
 sg13g2_xnor2_1 _4208_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[5] ),
    .A(_0422_),
    .B(_0438_));
 sg13g2_a21oi_1 _4209_ (.A1(_0422_),
    .A2(_0437_),
    .Y(_0439_),
    .B1(_0436_));
 sg13g2_o21ai_1 _4210_ (.B1(_0433_),
    .Y(_0440_),
    .A1(_0423_),
    .A2(_0434_));
 sg13g2_o21ai_1 _4211_ (.B1(_0428_),
    .Y(_0441_),
    .A1(_0429_),
    .A2(_0431_));
 sg13g2_nor3_2 _4212_ (.A(net1101),
    .B(_3389_),
    .C(_3419_),
    .Y(_0442_));
 sg13g2_a21oi_1 _4213_ (.A1(net1109),
    .A2(_3467_),
    .Y(_0443_),
    .B1(net1105));
 sg13g2_o21ai_1 _4214_ (.B1(_0443_),
    .Y(_0444_),
    .A1(net1108),
    .A2(_3462_));
 sg13g2_inv_1 _4215_ (.Y(_0445_),
    .A(_0444_));
 sg13g2_nand2_1 _4216_ (.Y(_0446_),
    .A(_0442_),
    .B(_0445_));
 sg13g2_xnor2_1 _4217_ (.Y(_0447_),
    .A(_0442_),
    .B(_0445_));
 sg13g2_xnor2_1 _4218_ (.Y(_0448_),
    .A(net1099),
    .B(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_xnor2_1 _4219_ (.Y(_0449_),
    .A(_0447_),
    .B(_0448_));
 sg13g2_nor2b_1 _4220_ (.A(_0449_),
    .B_N(_0441_),
    .Y(_0450_));
 sg13g2_xor2_1 _4221_ (.B(_0449_),
    .A(_0441_),
    .X(_0451_));
 sg13g2_inv_1 _4222_ (.Y(_0452_),
    .A(_0451_));
 sg13g2_xnor2_1 _4223_ (.Y(_0453_),
    .A(_0440_),
    .B(_0451_));
 sg13g2_nand2_1 _4224_ (.Y(_0454_),
    .A(\vgademo.soundtrack.sigma_delta_accum[6] ),
    .B(_0453_));
 sg13g2_xnor2_1 _4225_ (.Y(_0455_),
    .A(net520),
    .B(_0453_));
 sg13g2_xor2_1 _4226_ (.B(_0455_),
    .A(_0439_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[6] ));
 sg13g2_o21ai_1 _4227_ (.B1(_0454_),
    .Y(_0456_),
    .A1(_0439_),
    .A2(_0455_));
 sg13g2_a21oi_1 _4228_ (.A1(_0440_),
    .A2(_0452_),
    .Y(_0457_),
    .B1(_0450_));
 sg13g2_o21ai_1 _4229_ (.B1(_0446_),
    .Y(_0458_),
    .A1(_0447_),
    .A2(_0448_));
 sg13g2_o21ai_1 _4230_ (.B1(net1042),
    .Y(_0459_),
    .A1(net1110),
    .A2(_0387_));
 sg13g2_a21oi_1 _4231_ (.A1(net1108),
    .A2(_0392_),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_nor2_1 _4232_ (.A(net1101),
    .B(_3333_),
    .Y(_0461_));
 sg13g2_nor3_1 _4233_ (.A(\vgademo.soundtrack.pulse_vol[0] ),
    .B(net1101),
    .C(_3419_),
    .Y(_0462_));
 sg13g2_a22oi_1 _4234_ (.Y(_0463_),
    .B1(_0462_),
    .B2(_3387_),
    .A2(_0461_),
    .A1(\vgademo.soundtrack.pulse_vol[0] ));
 sg13g2_nor2b_1 _4235_ (.A(_0463_),
    .B_N(_0460_),
    .Y(_0464_));
 sg13g2_xnor2_1 _4236_ (.Y(_0465_),
    .A(_0460_),
    .B(_0463_));
 sg13g2_xor2_1 _4237_ (.B(\vgademo.soundtrack.tri_osc_p[8] ),
    .A(net1099),
    .X(_0466_));
 sg13g2_xor2_1 _4238_ (.B(_0466_),
    .A(_0465_),
    .X(_0467_));
 sg13g2_nand2_1 _4239_ (.Y(_0468_),
    .A(_0458_),
    .B(_0467_));
 sg13g2_xnor2_1 _4240_ (.Y(_0469_),
    .A(_0458_),
    .B(_0467_));
 sg13g2_xor2_1 _4241_ (.B(_0469_),
    .A(_0457_),
    .X(_0470_));
 sg13g2_xnor2_1 _4242_ (.Y(_0471_),
    .A(net499),
    .B(_0470_));
 sg13g2_nor2b_1 _4243_ (.A(_0471_),
    .B_N(_0456_),
    .Y(_0472_));
 sg13g2_xnor2_1 _4244_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .A(_0456_),
    .B(_0471_));
 sg13g2_a21oi_1 _4245_ (.A1(net499),
    .A2(_0470_),
    .Y(_0473_),
    .B1(_0472_));
 sg13g2_o21ai_1 _4246_ (.B1(_0468_),
    .Y(_0474_),
    .A1(_0457_),
    .A2(_0469_));
 sg13g2_a21oi_1 _4247_ (.A1(_0465_),
    .A2(_0466_),
    .Y(_0475_),
    .B1(_0464_));
 sg13g2_and2_1 _4248_ (.A(_3223_),
    .B(_3390_),
    .X(_0476_));
 sg13g2_and2_1 _4249_ (.A(net1042),
    .B(_3398_),
    .X(_0477_));
 sg13g2_nand2_1 _4250_ (.Y(_0478_),
    .A(_0476_),
    .B(_0477_));
 sg13g2_xnor2_1 _4251_ (.Y(_0479_),
    .A(_0476_),
    .B(_0477_));
 sg13g2_xnor2_1 _4252_ (.Y(_0480_),
    .A(net1099),
    .B(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_xnor2_1 _4253_ (.Y(_0481_),
    .A(_0479_),
    .B(_0480_));
 sg13g2_nor2_1 _4254_ (.A(_0475_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_xor2_1 _4255_ (.B(_0481_),
    .A(_0475_),
    .X(_0483_));
 sg13g2_xor2_1 _4256_ (.B(_0483_),
    .A(_0474_),
    .X(_0484_));
 sg13g2_nand2_1 _4257_ (.Y(_0485_),
    .A(\vgademo.soundtrack.sigma_delta_accum[8] ),
    .B(_0484_));
 sg13g2_xnor2_1 _4258_ (.Y(_0486_),
    .A(net529),
    .B(_0484_));
 sg13g2_xor2_1 _4259_ (.B(_0486_),
    .A(_0473_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[8] ));
 sg13g2_o21ai_1 _4260_ (.B1(_0485_),
    .Y(_0487_),
    .A1(_0473_),
    .A2(_0486_));
 sg13g2_a21oi_2 _4261_ (.B1(_0482_),
    .Y(_0488_),
    .A2(_0483_),
    .A1(_0474_));
 sg13g2_o21ai_1 _4262_ (.B1(_0478_),
    .Y(_0489_),
    .A1(_0479_),
    .A2(_0480_));
 sg13g2_nor3_2 _4263_ (.A(net1102),
    .B(_3422_),
    .C(_3428_),
    .Y(_0490_));
 sg13g2_nand2_1 _4264_ (.Y(_0491_),
    .A(net1042),
    .B(_3443_));
 sg13g2_nand3_1 _4265_ (.B(_3443_),
    .C(_0490_),
    .A(net1042),
    .Y(_0492_));
 sg13g2_xor2_1 _4266_ (.B(_0491_),
    .A(_0490_),
    .X(_0493_));
 sg13g2_xnor2_1 _4267_ (.Y(_0494_),
    .A(net1100),
    .B(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_xor2_1 _4268_ (.B(_0494_),
    .A(_0493_),
    .X(_0495_));
 sg13g2_nand2_1 _4269_ (.Y(_0496_),
    .A(_0489_),
    .B(_0495_));
 sg13g2_xnor2_1 _4270_ (.Y(_0497_),
    .A(_0489_),
    .B(_0495_));
 sg13g2_xor2_1 _4271_ (.B(_0497_),
    .A(_0488_),
    .X(_0498_));
 sg13g2_xnor2_1 _4272_ (.Y(_0499_),
    .A(net525),
    .B(_0498_));
 sg13g2_nor2b_1 _4273_ (.A(_0499_),
    .B_N(_0487_),
    .Y(_0500_));
 sg13g2_xnor2_1 _4274_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .A(_0487_),
    .B(_0499_));
 sg13g2_a21o_1 _4275_ (.A2(_0498_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[9] ),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_o21ai_1 _4276_ (.B1(_0496_),
    .Y(_0502_),
    .A1(_0488_),
    .A2(_0497_));
 sg13g2_o21ai_1 _4277_ (.B1(_0492_),
    .Y(_0503_),
    .A1(_0493_),
    .A2(_0494_));
 sg13g2_nor2_1 _4278_ (.A(net1101),
    .B(_3460_),
    .Y(_0504_));
 sg13g2_nor2_1 _4279_ (.A(net1106),
    .B(_3468_),
    .Y(_0505_));
 sg13g2_nand2_1 _4280_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_xnor2_1 _4281_ (.Y(_0507_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_xnor2_1 _4282_ (.Y(_0508_),
    .A(net1100),
    .B(\vgademo.soundtrack.tri_osc_p[11] ));
 sg13g2_xnor2_1 _4283_ (.Y(_0509_),
    .A(_0507_),
    .B(_0508_));
 sg13g2_inv_1 _4284_ (.Y(_0510_),
    .A(_0509_));
 sg13g2_xor2_1 _4285_ (.B(_0509_),
    .A(_0503_),
    .X(_0511_));
 sg13g2_nor2b_1 _4286_ (.A(_0511_),
    .B_N(_0502_),
    .Y(_0512_));
 sg13g2_xnor2_1 _4287_ (.Y(_0513_),
    .A(_0502_),
    .B(_0511_));
 sg13g2_xnor2_1 _4288_ (.Y(_0514_),
    .A(net510),
    .B(_0513_));
 sg13g2_nor2b_1 _4289_ (.A(_0514_),
    .B_N(_0501_),
    .Y(_0515_));
 sg13g2_xnor2_1 _4290_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .A(_0501_),
    .B(_0514_));
 sg13g2_a21o_1 _4291_ (.A2(_0513_),
    .A1(net510),
    .B1(_0515_),
    .X(_0516_));
 sg13g2_a21oi_1 _4292_ (.A1(_0503_),
    .A2(_0510_),
    .Y(_0517_),
    .B1(_0512_));
 sg13g2_o21ai_1 _4293_ (.B1(_0506_),
    .Y(_0518_),
    .A1(_0507_),
    .A2(_0508_));
 sg13g2_nand2b_1 _4294_ (.Y(_0519_),
    .B(_3421_),
    .A_N(_0384_));
 sg13g2_nand2_1 _4295_ (.Y(_0520_),
    .A(net1042),
    .B(_0393_));
 sg13g2_nor2_1 _4296_ (.A(_0519_),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_xor2_1 _4297_ (.B(_0520_),
    .A(_0519_),
    .X(_0522_));
 sg13g2_xor2_1 _4298_ (.B(\vgademo.soundtrack.tri_osc_p[12] ),
    .A(net1100),
    .X(_0523_));
 sg13g2_xnor2_1 _4299_ (.Y(_0524_),
    .A(_0522_),
    .B(_0523_));
 sg13g2_nand2b_1 _4300_ (.Y(_0525_),
    .B(_0518_),
    .A_N(_0524_));
 sg13g2_xor2_1 _4301_ (.B(_0524_),
    .A(_0518_),
    .X(_0526_));
 sg13g2_xor2_1 _4302_ (.B(_0526_),
    .A(_0517_),
    .X(_0527_));
 sg13g2_xnor2_1 _4303_ (.Y(_0528_),
    .A(net513),
    .B(_0527_));
 sg13g2_nor2b_1 _4304_ (.A(_0528_),
    .B_N(_0516_),
    .Y(_0529_));
 sg13g2_xnor2_1 _4305_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .A(_0516_),
    .B(_0528_));
 sg13g2_a21o_1 _4306_ (.A2(_0527_),
    .A1(net513),
    .B1(_0529_),
    .X(_0530_));
 sg13g2_o21ai_1 _4307_ (.B1(_0525_),
    .Y(_0531_),
    .A1(_0517_),
    .A2(_0526_));
 sg13g2_a21oi_1 _4308_ (.A1(_0522_),
    .A2(_0523_),
    .Y(_0532_),
    .B1(_0521_));
 sg13g2_nor4_2 _4309_ (.A(net1104),
    .B(net1103),
    .C(net1102),
    .Y(_0533_),
    .D(_3389_));
 sg13g2_nor3_1 _4310_ (.A(net1106),
    .B(net1110),
    .C(_3397_),
    .Y(_0534_));
 sg13g2_nand2_1 _4311_ (.Y(_0535_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_xnor2_1 _4312_ (.Y(_0536_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_xor2_1 _4313_ (.B(\vgademo.soundtrack.tri_osc_p[13] ),
    .A(net1100),
    .X(_0537_));
 sg13g2_inv_1 _4314_ (.Y(_0538_),
    .A(_0537_));
 sg13g2_xnor2_1 _4315_ (.Y(_0539_),
    .A(_0536_),
    .B(_0538_));
 sg13g2_nor2_1 _4316_ (.A(_0532_),
    .B(_0539_),
    .Y(_0540_));
 sg13g2_nand2_1 _4317_ (.Y(_0541_),
    .A(_0532_),
    .B(_0539_));
 sg13g2_nand2b_1 _4318_ (.Y(_0542_),
    .B(_0541_),
    .A_N(_0540_));
 sg13g2_xnor2_1 _4319_ (.Y(_0543_),
    .A(_0531_),
    .B(_0542_));
 sg13g2_xnor2_1 _4320_ (.Y(_0544_),
    .A(net514),
    .B(_0543_));
 sg13g2_nor2b_1 _4321_ (.A(_0544_),
    .B_N(_0530_),
    .Y(_0545_));
 sg13g2_xnor2_1 _4322_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .A(_0530_),
    .B(_0544_));
 sg13g2_a21o_1 _4323_ (.A2(_0543_),
    .A1(net514),
    .B1(_0545_),
    .X(_0546_));
 sg13g2_a21o_1 _4324_ (.A2(_0541_),
    .A1(_0531_),
    .B1(_0540_),
    .X(_0547_));
 sg13g2_o21ai_1 _4325_ (.B1(_0535_),
    .Y(_0548_),
    .A1(_0536_),
    .A2(_0538_));
 sg13g2_inv_1 _4326_ (.Y(_0549_),
    .A(_0548_));
 sg13g2_nor4_2 _4327_ (.A(net1104),
    .B(\vgademo.soundtrack.pulse_vol[2] ),
    .C(net1102),
    .Y(_0550_),
    .D(_3428_));
 sg13g2_nand2b_1 _4328_ (.Y(_0551_),
    .B(net366),
    .A_N(net1100));
 sg13g2_xnor2_1 _4329_ (.Y(_0552_),
    .A(\vgademo.soundtrack.tri_osc_p[14] ),
    .B(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_nand2b_1 _4330_ (.Y(_0553_),
    .B(_0552_),
    .A_N(_0550_));
 sg13g2_xnor2_1 _4331_ (.Y(_0554_),
    .A(_0550_),
    .B(_0552_));
 sg13g2_xnor2_1 _4332_ (.Y(_0555_),
    .A(_0548_),
    .B(_0554_));
 sg13g2_nand2_1 _4333_ (.Y(_0556_),
    .A(_0547_),
    .B(_0555_));
 sg13g2_xor2_1 _4334_ (.B(_0555_),
    .A(_0547_),
    .X(_0557_));
 sg13g2_xnor2_1 _4335_ (.Y(_0558_),
    .A(net519),
    .B(_0557_));
 sg13g2_nor2b_1 _4336_ (.A(_0558_),
    .B_N(_0546_),
    .Y(_0559_));
 sg13g2_xnor2_1 _4337_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .A(_0546_),
    .B(_0558_));
 sg13g2_a21o_1 _4338_ (.A2(_0557_),
    .A1(net519),
    .B1(_0559_),
    .X(_0560_));
 sg13g2_o21ai_1 _4339_ (.B1(_0556_),
    .Y(_0561_),
    .A1(_0549_),
    .A2(_0554_));
 sg13g2_or2_1 _4340_ (.X(_0562_),
    .B(_0561_),
    .A(_0553_));
 sg13g2_xnor2_1 _4341_ (.Y(_0563_),
    .A(_0553_),
    .B(_0561_));
 sg13g2_and2_1 _4342_ (.A(net561),
    .B(_0563_),
    .X(_0564_));
 sg13g2_xor2_1 _4343_ (.B(_0563_),
    .A(net561),
    .X(_0565_));
 sg13g2_xor2_1 _4344_ (.B(_0565_),
    .A(_0560_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[14] ));
 sg13g2_a21o_1 _4345_ (.A2(_0565_),
    .A1(_0560_),
    .B1(_0564_),
    .X(_0566_));
 sg13g2_and2_1 _4346_ (.A(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .B(_0562_),
    .X(_0567_));
 sg13g2_xor2_1 _4347_ (.B(_0562_),
    .A(net576),
    .X(_0568_));
 sg13g2_xor2_1 _4348_ (.B(_0568_),
    .A(_0566_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[15] ));
 sg13g2_xor2_1 _4349_ (.B(net258),
    .A(\vgademo.soundtrack.sample_div[0] ),
    .X(\vgademo.soundtrack.sample_div_[1] ));
 sg13g2_nand3_1 _4350_ (.B(net465),
    .C(net258),
    .A(\vgademo.soundtrack.sample_div[0] ),
    .Y(_0569_));
 sg13g2_a21o_1 _4351_ (.A2(net258),
    .A1(\vgademo.soundtrack.sample_div[0] ),
    .B1(net465),
    .X(_0570_));
 sg13g2_and2_1 _4352_ (.A(_0569_),
    .B(net466),
    .X(\vgademo.soundtrack.sample_div_[2] ));
 sg13g2_nor2_1 _4353_ (.A(_3174_),
    .B(_0569_),
    .Y(_0571_));
 sg13g2_xnor2_1 _4354_ (.Y(\vgademo.soundtrack.sample_div_[3] ),
    .A(net254),
    .B(_0569_));
 sg13g2_and2_1 _4355_ (.A(net215),
    .B(_0571_),
    .X(_0572_));
 sg13g2_xor2_1 _4356_ (.B(_0571_),
    .A(net215),
    .X(\vgademo.soundtrack.sample_div_[4] ));
 sg13g2_xor2_1 _4357_ (.B(_0572_),
    .A(net273),
    .X(\vgademo.soundtrack.sample_div_[5] ));
 sg13g2_nand3_1 _4358_ (.B(net273),
    .C(_0572_),
    .A(net459),
    .Y(_0573_));
 sg13g2_a21o_1 _4359_ (.A2(_0572_),
    .A1(net273),
    .B1(net459),
    .X(_0574_));
 sg13g2_and2_1 _4360_ (.A(_0573_),
    .B(_0574_),
    .X(\vgademo.soundtrack.sample_div_[6] ));
 sg13g2_nor2_1 _4361_ (.A(_3173_),
    .B(_0573_),
    .Y(_0575_));
 sg13g2_xnor2_1 _4362_ (.Y(\vgademo.soundtrack.sample_div_[7] ),
    .A(net228),
    .B(_0573_));
 sg13g2_and2_1 _4363_ (.A(\vgademo.soundtrack.sample_div[8] ),
    .B(_0575_),
    .X(_0576_));
 sg13g2_xor2_1 _4364_ (.B(_0575_),
    .A(net224),
    .X(\vgademo.soundtrack.sample_div_[8] ));
 sg13g2_and2_1 _4365_ (.A(net284),
    .B(_0576_),
    .X(_0577_));
 sg13g2_nand2_1 _4366_ (.Y(_0578_),
    .A(net284),
    .B(_0576_));
 sg13g2_xor2_1 _4367_ (.B(_0576_),
    .A(net284),
    .X(\vgademo.soundtrack.sample_div_[9] ));
 sg13g2_nor4_2 _4368_ (.A(\vgademo.h_count[5] ),
    .B(\vgademo.h_count[4] ),
    .C(_3283_),
    .Y(_0579_),
    .D(_3286_));
 sg13g2_and2_1 _4369_ (.A(_3330_),
    .B(_0579_),
    .X(_0580_));
 sg13g2_nand2_1 _4370_ (.Y(_0581_),
    .A(_3330_),
    .B(_0579_));
 sg13g2_and2_2 _4371_ (.A(net1174),
    .B(net1034),
    .X(_0582_));
 sg13g2_nand2_1 _4372_ (.Y(_0583_),
    .A(net1174),
    .B(net1034));
 sg13g2_nor2_1 _4373_ (.A(net1006),
    .B(net1025),
    .Y(_0584_));
 sg13g2_nor3_1 _4374_ (.A(net1060),
    .B(net1061),
    .C(\vgademo.v_count[8] ),
    .Y(_0585_));
 sg13g2_nand2_1 _4375_ (.Y(_0586_),
    .A(net1059),
    .B(_0585_));
 sg13g2_nand2_2 _4376_ (.Y(_0587_),
    .A(_3183_),
    .B(_3184_));
 sg13g2_nand2_1 _4377_ (.Y(_0588_),
    .A(net1064),
    .B(net1065));
 sg13g2_nor4_1 _4378_ (.A(net1062),
    .B(\vgademo.v_count[5] ),
    .C(_0587_),
    .D(_0588_),
    .Y(_0589_));
 sg13g2_nand2b_2 _4379_ (.Y(_0590_),
    .B(_0589_),
    .A_N(_0586_));
 sg13g2_nand2b_1 _4380_ (.Y(_0591_),
    .B(_3185_),
    .A_N(_0588_));
 sg13g2_nor4_2 _4381_ (.A(net1062),
    .B(_0586_),
    .C(_0587_),
    .Y(_0592_),
    .D(_0591_));
 sg13g2_and2_1 _4382_ (.A(net1036),
    .B(_0592_),
    .X(_0593_));
 sg13g2_nand2_1 _4383_ (.Y(_0594_),
    .A(net1036),
    .B(_0592_));
 sg13g2_nor2_1 _4384_ (.A(net1033),
    .B(_0590_),
    .Y(_0595_));
 sg13g2_a21o_1 _4385_ (.A2(net999),
    .A1(net1162),
    .B1(net987),
    .X(_0596_));
 sg13g2_a21oi_1 _4386_ (.A1(net1154),
    .A2(net974),
    .Y(_0597_),
    .B1(net1156));
 sg13g2_nand2b_1 _4387_ (.Y(_0598_),
    .B(net1011),
    .A_N(net1157));
 sg13g2_a21o_1 _4388_ (.A2(net1154),
    .A1(net1156),
    .B1(net1000),
    .X(_0599_));
 sg13g2_a21oi_1 _4389_ (.A1(net974),
    .A2(_0599_),
    .Y(_0111_),
    .B1(_0597_));
 sg13g2_nor2_1 _4390_ (.A(net1153),
    .B(net976),
    .Y(_0600_));
 sg13g2_nor2_1 _4391_ (.A(net537),
    .B(net1000),
    .Y(_0601_));
 sg13g2_a21oi_1 _4392_ (.A1(net976),
    .A2(_0601_),
    .Y(_0112_),
    .B1(_0600_));
 sg13g2_nand3_1 _4393_ (.B(net1011),
    .C(net975),
    .A(net370),
    .Y(_0602_));
 sg13g2_o21ai_1 _4394_ (.B1(_0602_),
    .Y(_0113_),
    .A1(_3169_),
    .A2(net975));
 sg13g2_nor2_1 _4395_ (.A(net370),
    .B(net975),
    .Y(_0603_));
 sg13g2_xor2_1 _4396_ (.B(net395),
    .A(net1157),
    .X(_0604_));
 sg13g2_nor2_1 _4397_ (.A(net1000),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_a21oi_1 _4398_ (.A1(net975),
    .A2(_0605_),
    .Y(_0114_),
    .B1(_0603_));
 sg13g2_nor2_1 _4399_ (.A(net395),
    .B(net975),
    .Y(_0606_));
 sg13g2_xor2_1 _4400_ (.B(net412),
    .A(net1157),
    .X(_0607_));
 sg13g2_nor2_1 _4401_ (.A(net1000),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_a21oi_1 _4402_ (.A1(net975),
    .A2(_0608_),
    .Y(_0115_),
    .B1(_0606_));
 sg13g2_nor2_1 _4403_ (.A(net412),
    .B(net975),
    .Y(_0609_));
 sg13g2_nor2_1 _4404_ (.A(net319),
    .B(net1000),
    .Y(_0610_));
 sg13g2_a21oi_1 _4405_ (.A1(net975),
    .A2(_0610_),
    .Y(_0116_),
    .B1(_0609_));
 sg13g2_nor2_1 _4406_ (.A(net319),
    .B(net974),
    .Y(_0611_));
 sg13g2_xor2_1 _4407_ (.B(\vgademo.linelfsr[7] ),
    .A(net1155),
    .X(_0612_));
 sg13g2_nor2_1 _4408_ (.A(net1000),
    .B(_0612_),
    .Y(_0613_));
 sg13g2_a21oi_1 _4409_ (.A1(net976),
    .A2(_0613_),
    .Y(_0117_),
    .B1(_0611_));
 sg13g2_nor2_1 _4410_ (.A(net368),
    .B(net974),
    .Y(_0614_));
 sg13g2_nor2_1 _4411_ (.A(\vgademo.linelfsr[8] ),
    .B(net1000),
    .Y(_0615_));
 sg13g2_a21oi_1 _4412_ (.A1(net974),
    .A2(_0615_),
    .Y(_0118_),
    .B1(_0614_));
 sg13g2_nor2_1 _4413_ (.A(net376),
    .B(net974),
    .Y(_0616_));
 sg13g2_xor2_1 _4414_ (.B(\vgademo.linelfsr[9] ),
    .A(net1156),
    .X(_0617_));
 sg13g2_nand2_1 _4415_ (.Y(_0618_),
    .A(net1011),
    .B(_0617_));
 sg13g2_a21oi_1 _4416_ (.A1(net974),
    .A2(_0618_),
    .Y(_0119_),
    .B1(_0616_));
 sg13g2_nor2_1 _4417_ (.A(net403),
    .B(net974),
    .Y(_0619_));
 sg13g2_nor2_1 _4418_ (.A(\vgademo.linelfsr[10] ),
    .B(net1000),
    .Y(_0620_));
 sg13g2_a21oi_1 _4419_ (.A1(net976),
    .A2(_0620_),
    .Y(_0120_),
    .B1(_0619_));
 sg13g2_nand3_1 _4420_ (.B(net1011),
    .C(net977),
    .A(net401),
    .Y(_0621_));
 sg13g2_o21ai_1 _4421_ (.B1(_0621_),
    .Y(_0121_),
    .A1(_3167_),
    .A2(net977));
 sg13g2_nor2_1 _4422_ (.A(net401),
    .B(net977),
    .Y(_0622_));
 sg13g2_nor2_1 _4423_ (.A(net409),
    .B(net1007),
    .Y(_0623_));
 sg13g2_a21oi_1 _4424_ (.A1(net977),
    .A2(_0623_),
    .Y(_0122_),
    .B1(_0622_));
 sg13g2_mux2_1 _4425_ (.A0(net409),
    .A1(_0598_),
    .S(net977),
    .X(_0123_));
 sg13g2_nand3_1 _4426_ (.B(net489),
    .C(net981),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0624_));
 sg13g2_nand4_1 _4427_ (.B(net242),
    .C(\vgademo.soundtrack.tick_div[1] ),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0625_),
    .D(net980));
 sg13g2_nor2_1 _4428_ (.A(_3175_),
    .B(_0625_),
    .Y(_0626_));
 sg13g2_and2_1 _4429_ (.A(net226),
    .B(_0626_),
    .X(_0627_));
 sg13g2_and3_1 _4430_ (.X(_0628_),
    .A(net199),
    .B(\vgademo.soundtrack.tick_div[5] ),
    .C(_0627_));
 sg13g2_and2_1 _4431_ (.A(\vgademo.soundtrack.tick_div[7] ),
    .B(_0628_),
    .X(_0629_));
 sg13g2_or2_1 _4432_ (.X(_0630_),
    .B(\vgademo.audio_beat_out[0] ),
    .A(\vgademo.audio_beat_out[1] ));
 sg13g2_nor4_2 _4433_ (.A(\vgademo.audio_beat_out[3] ),
    .B(\vgademo.audio_beat_out[2] ),
    .C(\vgademo.audio_beat_out[4] ),
    .Y(_0631_),
    .D(_0630_));
 sg13g2_or4_1 _4434_ (.A(\vgademo.audio_beat_out[3] ),
    .B(\vgademo.audio_beat_out[2] ),
    .C(\vgademo.audio_beat_out[4] ),
    .D(_0630_),
    .X(_0632_));
 sg13g2_nand2_1 _4435_ (.Y(_0633_),
    .A(net949),
    .B(net1039));
 sg13g2_nand3_1 _4436_ (.B(net950),
    .C(net1039),
    .A(_3170_),
    .Y(_0634_));
 sg13g2_mux2_1 _4437_ (.A0(net1151),
    .A1(net271),
    .S(net945),
    .X(_0124_));
 sg13g2_nand2_1 _4438_ (.Y(_0635_),
    .A(net191),
    .B(net946));
 sg13g2_o21ai_1 _4439_ (.B1(_0635_),
    .Y(_0125_),
    .A1(_3364_),
    .A2(net946));
 sg13g2_nor2_1 _4440_ (.A(_3170_),
    .B(_3179_),
    .Y(_0636_));
 sg13g2_nand2_2 _4441_ (.Y(_0637_),
    .A(net1146),
    .B(_3362_));
 sg13g2_nor2_1 _4442_ (.A(net1146),
    .B(_3362_),
    .Y(_0638_));
 sg13g2_nor2b_1 _4443_ (.A(_0638_),
    .B_N(_0637_),
    .Y(_0639_));
 sg13g2_nand2_1 _4444_ (.Y(_0640_),
    .A(net185),
    .B(net945));
 sg13g2_o21ai_1 _4445_ (.B1(_0640_),
    .Y(_0126_),
    .A1(net945),
    .A2(_0639_));
 sg13g2_xnor2_1 _4446_ (.Y(_0641_),
    .A(net1049),
    .B(_0637_));
 sg13g2_xnor2_1 _4447_ (.Y(_0642_),
    .A(net1143),
    .B(_0637_));
 sg13g2_nand2_1 _4448_ (.Y(_0643_),
    .A(net213),
    .B(net944));
 sg13g2_o21ai_1 _4449_ (.B1(_0643_),
    .Y(_0127_),
    .A1(net944),
    .A2(_0642_));
 sg13g2_nand2_2 _4450_ (.Y(_0644_),
    .A(net1137),
    .B(net1141));
 sg13g2_nor2_2 _4451_ (.A(_0637_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_nor2_1 _4452_ (.A(_3340_),
    .B(_3363_),
    .Y(_0646_));
 sg13g2_nor2_2 _4453_ (.A(net1139),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_nor2_1 _4454_ (.A(_0645_),
    .B(_0647_),
    .Y(_0648_));
 sg13g2_nand2_1 _4455_ (.Y(_0649_),
    .A(net195),
    .B(net945));
 sg13g2_o21ai_1 _4456_ (.B1(_0649_),
    .Y(_0128_),
    .A1(net944),
    .A2(net1017));
 sg13g2_nand3_1 _4457_ (.B(net1141),
    .C(net1135),
    .A(net1138),
    .Y(_0650_));
 sg13g2_nor2_1 _4458_ (.A(_0637_),
    .B(_0650_),
    .Y(_0651_));
 sg13g2_xnor2_1 _4459_ (.Y(_0652_),
    .A(net1046),
    .B(_0645_));
 sg13g2_nand2_1 _4460_ (.Y(_0653_),
    .A(net208),
    .B(net944));
 sg13g2_o21ai_1 _4461_ (.B1(_0653_),
    .Y(_0129_),
    .A1(net944),
    .A2(_0652_));
 sg13g2_nand2_1 _4462_ (.Y(_0654_),
    .A(net1132),
    .B(_0651_));
 sg13g2_xnor2_1 _4463_ (.Y(_0655_),
    .A(net1132),
    .B(_0651_));
 sg13g2_mux2_1 _4464_ (.A0(_0655_),
    .A1(net276),
    .S(net944),
    .X(_0130_));
 sg13g2_xnor2_1 _4465_ (.Y(_0656_),
    .A(\vgademo.audio_songpos[7] ),
    .B(_0654_));
 sg13g2_nand2_1 _4466_ (.Y(_0657_),
    .A(net189),
    .B(net944));
 sg13g2_o21ai_1 _4467_ (.B1(_0657_),
    .Y(_0131_),
    .A1(net944),
    .A2(_0656_));
 sg13g2_nor2_1 _4468_ (.A(\vgademo.plane_dx_div.i[1] ),
    .B(net327),
    .Y(_0658_));
 sg13g2_nor4_2 _4469_ (.A(net405),
    .B(net477),
    .C(net543),
    .Y(_0659_),
    .D(net327));
 sg13g2_nor4_2 _4470_ (.A(_3192_),
    .B(_3193_),
    .C(_3194_),
    .Y(_0660_),
    .D(\vgademo.h_count[6] ));
 sg13g2_and3_1 _4471_ (.X(_0661_),
    .A(_3285_),
    .B(_3330_),
    .C(_0660_));
 sg13g2_and3_2 _4472_ (.X(_0662_),
    .A(_3285_),
    .B(_3330_),
    .C(_0660_));
 sg13g2_nand3_1 _4473_ (.B(_3330_),
    .C(_0660_),
    .A(_3285_),
    .Y(_0663_));
 sg13g2_nor2_1 _4474_ (.A(_0659_),
    .B(net1032),
    .Y(_0664_));
 sg13g2_nor2b_2 _4475_ (.A(net1032),
    .B_N(_0659_),
    .Y(_0665_));
 sg13g2_nand2_2 _4476_ (.Y(_0666_),
    .A(_0659_),
    .B(_0663_));
 sg13g2_a22oi_1 _4477_ (.Y(_0132_),
    .B1(_0665_),
    .B2(_3165_),
    .A2(_0664_),
    .A1(_3166_));
 sg13g2_a22oi_1 _4478_ (.Y(_0667_),
    .B1(net1013),
    .B2(\vgademo.plane_dx[2] ),
    .A2(net1015),
    .A1(net531));
 sg13g2_inv_1 _4479_ (.Y(_0133_),
    .A(net532));
 sg13g2_a22oi_1 _4480_ (.Y(_0668_),
    .B1(_0665_),
    .B2(net1130),
    .A2(net1015),
    .A1(\vgademo.plane_dx[2] ));
 sg13g2_inv_1 _4481_ (.Y(_0134_),
    .A(net524));
 sg13g2_a22oi_1 _4482_ (.Y(_0669_),
    .B1(_0665_),
    .B2(net206),
    .A2(net1015),
    .A1(\vgademo.plane_dx[3] ));
 sg13g2_inv_1 _4483_ (.Y(_0135_),
    .A(net207));
 sg13g2_a22oi_1 _4484_ (.Y(_0670_),
    .B1(net1013),
    .B2(net1127),
    .A2(net1015),
    .A1(net206));
 sg13g2_inv_1 _4485_ (.Y(_0136_),
    .A(_0670_));
 sg13g2_a22oi_1 _4486_ (.Y(_0671_),
    .B1(net1013),
    .B2(net421),
    .A2(net1015),
    .A1(net1128));
 sg13g2_inv_1 _4487_ (.Y(_0137_),
    .A(_0671_));
 sg13g2_a22oi_1 _4488_ (.Y(_0672_),
    .B1(net1012),
    .B2(net1125),
    .A2(net1014),
    .A1(net1126));
 sg13g2_inv_1 _4489_ (.Y(_0138_),
    .A(_0672_));
 sg13g2_a22oi_1 _4490_ (.Y(_0673_),
    .B1(net1012),
    .B2(net1123),
    .A2(net1014),
    .A1(net1125));
 sg13g2_inv_1 _4491_ (.Y(_0139_),
    .A(_0673_));
 sg13g2_a22oi_1 _4492_ (.Y(_0674_),
    .B1(net1012),
    .B2(net1122),
    .A2(net1014),
    .A1(net1123));
 sg13g2_inv_1 _4493_ (.Y(_0140_),
    .A(net540));
 sg13g2_a22oi_1 _4494_ (.Y(_0675_),
    .B1(net1012),
    .B2(net1119),
    .A2(net1014),
    .A1(net1121));
 sg13g2_inv_1 _4495_ (.Y(_0141_),
    .A(_0675_));
 sg13g2_o21ai_1 _4496_ (.B1(_0666_),
    .Y(_0676_),
    .A1(net217),
    .A2(_0662_));
 sg13g2_inv_1 _4497_ (.Y(_0142_),
    .A(_0676_));
 sg13g2_and2_1 _4498_ (.A(\vgademo.plane_dx_div.i[1] ),
    .B(net327),
    .X(_0677_));
 sg13g2_nor3_1 _4499_ (.A(net328),
    .B(net1032),
    .C(_0677_),
    .Y(_0143_));
 sg13g2_nand2_1 _4500_ (.Y(_0678_),
    .A(net477),
    .B(_0677_));
 sg13g2_o21ai_1 _4501_ (.B1(_0663_),
    .Y(_0679_),
    .A1(net477),
    .A2(_0677_));
 sg13g2_nor2b_1 _4502_ (.A(net478),
    .B_N(_0678_),
    .Y(_0144_));
 sg13g2_xor2_1 _4503_ (.B(_0678_),
    .A(net405),
    .X(_0680_));
 sg13g2_nor2_1 _4504_ (.A(net1032),
    .B(net406),
    .Y(_0145_));
 sg13g2_nand2_2 _4505_ (.Y(_0681_),
    .A(net949),
    .B(net1038));
 sg13g2_a21oi_1 _4506_ (.A1(net950),
    .A2(_0632_),
    .Y(_0682_),
    .B1(net318));
 sg13g2_a21oi_1 _4507_ (.A1(net318),
    .A2(net950),
    .Y(_0146_),
    .B1(_0682_));
 sg13g2_and3_1 _4508_ (.X(_0683_),
    .A(net375),
    .B(net318),
    .C(net949));
 sg13g2_nand3_1 _4509_ (.B(net318),
    .C(net949),
    .A(net375),
    .Y(_0684_));
 sg13g2_a21oi_1 _4510_ (.A1(net318),
    .A2(net949),
    .Y(_0685_),
    .B1(net375));
 sg13g2_o21ai_1 _4511_ (.B1(_0634_),
    .Y(_0147_),
    .A1(_0683_),
    .A2(_0685_));
 sg13g2_nor2_1 _4512_ (.A(_0061_),
    .B(_0684_),
    .Y(_0686_));
 sg13g2_o21ai_1 _4513_ (.B1(net946),
    .Y(_0687_),
    .A1(net550),
    .A2(_0684_));
 sg13g2_mux2_1 _4514_ (.A0(_3176_),
    .A1(net550),
    .S(net950),
    .X(_0688_));
 sg13g2_a21oi_1 _4515_ (.A1(_0684_),
    .A2(_0688_),
    .Y(_0148_),
    .B1(_0687_));
 sg13g2_o21ai_1 _4516_ (.B1(_0634_),
    .Y(_0689_),
    .A1(net407),
    .A2(_0687_));
 sg13g2_a21oi_1 _4517_ (.A1(net407),
    .A2(_0686_),
    .Y(_0149_),
    .B1(_0689_));
 sg13g2_nand3_1 _4518_ (.B(\vgademo.audio_beat_out[2] ),
    .C(_0683_),
    .A(net407),
    .Y(_0690_));
 sg13g2_xor2_1 _4519_ (.B(_0690_),
    .A(net505),
    .X(_0691_));
 sg13g2_nand2_1 _4520_ (.Y(_0150_),
    .A(_0634_),
    .B(net506));
 sg13g2_o21ai_1 _4521_ (.B1(_0642_),
    .Y(_0692_),
    .A1(net1146),
    .A2(_3364_));
 sg13g2_nor2_1 _4522_ (.A(net1143),
    .B(_3362_),
    .Y(_0693_));
 sg13g2_a21oi_1 _4523_ (.A1(_3359_),
    .A2(_0693_),
    .Y(_0694_),
    .B1(_0652_));
 sg13g2_nand2_1 _4524_ (.Y(_0695_),
    .A(_0692_),
    .B(_0694_));
 sg13g2_nor2_1 _4525_ (.A(net1047),
    .B(net1133),
    .Y(_0696_));
 sg13g2_nor3_1 _4526_ (.A(_0645_),
    .B(_0647_),
    .C(_0696_),
    .Y(_0697_));
 sg13g2_nor2_2 _4527_ (.A(net1140),
    .B(_3179_),
    .Y(_0698_));
 sg13g2_nand2_1 _4528_ (.Y(_0699_),
    .A(net1048),
    .B(net1145));
 sg13g2_a21oi_1 _4529_ (.A1(_3356_),
    .A2(_0698_),
    .Y(_0700_),
    .B1(net1047));
 sg13g2_nand2b_1 _4530_ (.Y(_0701_),
    .B(net1016),
    .A_N(_0700_));
 sg13g2_a22oi_1 _4531_ (.Y(_0702_),
    .B1(_0701_),
    .B2(_3363_),
    .A2(_0697_),
    .A1(_0695_));
 sg13g2_o21ai_1 _4532_ (.B1(net949),
    .Y(_0703_),
    .A1(net1038),
    .A2(_0702_));
 sg13g2_nor3_2 _4533_ (.A(net460),
    .B(\vgademo.audio_kick_frames[0] ),
    .C(_3182_),
    .Y(_0704_));
 sg13g2_or3_1 _4534_ (.A(\vgademo.audio_kick_frames[1] ),
    .B(\vgademo.audio_kick_frames[0] ),
    .C(_3182_),
    .X(_0705_));
 sg13g2_nand2b_2 _4535_ (.Y(_0706_),
    .B(net1144),
    .A_N(net1147));
 sg13g2_and2_1 _4536_ (.A(_3379_),
    .B(_0706_),
    .X(_0707_));
 sg13g2_nand2_1 _4537_ (.Y(_0708_),
    .A(_3379_),
    .B(_0706_));
 sg13g2_a221oi_1 _4538_ (.B2(net1137),
    .C1(net1047),
    .B1(_0708_),
    .A1(_3344_),
    .Y(_0709_),
    .A2(_3347_));
 sg13g2_a21oi_1 _4539_ (.A1(net1048),
    .A2(_0708_),
    .Y(_0710_),
    .B1(_3337_));
 sg13g2_nor2_1 _4540_ (.A(net1141),
    .B(_3359_),
    .Y(_0711_));
 sg13g2_nor2_1 _4541_ (.A(_3348_),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_nor3_2 _4542_ (.A(_0709_),
    .B(_0710_),
    .C(_0712_),
    .Y(_0713_));
 sg13g2_and2_1 _4543_ (.A(_0704_),
    .B(_0713_),
    .X(_0714_));
 sg13g2_nor2_1 _4544_ (.A(_3177_),
    .B(net1141),
    .Y(_0715_));
 sg13g2_nand2_1 _4545_ (.Y(_0716_),
    .A(net1139),
    .B(net1048));
 sg13g2_nor2_1 _4546_ (.A(_3378_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_and2_1 _4547_ (.A(net1147),
    .B(_3340_),
    .X(_0718_));
 sg13g2_a21oi_2 _4548_ (.B1(net1047),
    .Y(_0719_),
    .A2(_0718_),
    .A1(_3344_));
 sg13g2_nand2b_1 _4549_ (.Y(_0720_),
    .B(_3379_),
    .A_N(_0644_));
 sg13g2_nand2b_1 _4550_ (.Y(_0721_),
    .B(_0715_),
    .A_N(_0706_));
 sg13g2_a21oi_1 _4551_ (.A1(_3177_),
    .A2(_3379_),
    .Y(_0722_),
    .B1(net1134));
 sg13g2_a22oi_1 _4552_ (.Y(_0723_),
    .B1(_0721_),
    .B2(_0722_),
    .A2(_0720_),
    .A1(_0719_));
 sg13g2_a22oi_1 _4553_ (.Y(_0724_),
    .B1(_0723_),
    .B2(_3336_),
    .A2(_0717_),
    .A1(net1134));
 sg13g2_nor2_1 _4554_ (.A(net1037),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_nand2b_1 _4555_ (.Y(_0726_),
    .B(\vgademo.soundtrack.tri_osc_i[3] ),
    .A_N(\vgademo.soundtrack.tri_osc_i[0] ));
 sg13g2_xor2_1 _4556_ (.B(\vgademo.soundtrack.tri_osc_i[3] ),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(_0727_));
 sg13g2_nor2_1 _4557_ (.A(net1039),
    .B(net1037),
    .Y(_0728_));
 sg13g2_o21ai_1 _4558_ (.B1(net1038),
    .Y(_0729_),
    .A1(_0704_),
    .A2(_0727_));
 sg13g2_nor4_1 _4559_ (.A(net942),
    .B(_0714_),
    .C(_0725_),
    .D(_0729_),
    .Y(_0730_));
 sg13g2_a21o_1 _4560_ (.A2(net942),
    .A1(net429),
    .B1(_0730_),
    .X(_0151_));
 sg13g2_nand2_1 _4561_ (.Y(_0731_),
    .A(net430),
    .B(net942));
 sg13g2_o21ai_1 _4562_ (.B1(_3345_),
    .Y(_0732_),
    .A1(net1144),
    .A2(_3347_));
 sg13g2_o21ai_1 _4563_ (.B1(_0732_),
    .Y(_0733_),
    .A1(net1047),
    .A2(_0717_));
 sg13g2_nand2_1 _4564_ (.Y(_0734_),
    .A(_0723_),
    .B(_0733_));
 sg13g2_inv_1 _4565_ (.Y(_0735_),
    .A(_0734_));
 sg13g2_nor2_2 _4566_ (.A(net1037),
    .B(_0713_),
    .Y(_0736_));
 sg13g2_nor2b_1 _4567_ (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[1] ),
    .Y(_0737_));
 sg13g2_xnor2_1 _4568_ (.Y(_0738_),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .B(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_xor2_1 _4569_ (.B(_0738_),
    .A(_0726_),
    .X(_0739_));
 sg13g2_a22oi_1 _4570_ (.Y(_0740_),
    .B1(_0735_),
    .B2(_0736_),
    .A2(_0725_),
    .A1(_0713_));
 sg13g2_o21ai_1 _4571_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0704_),
    .A2(_0739_));
 sg13g2_o21ai_1 _4572_ (.B1(_0731_),
    .Y(_0152_),
    .A1(_0681_),
    .A2(_0741_));
 sg13g2_nor2_1 _4573_ (.A(_0715_),
    .B(_0723_),
    .Y(_0742_));
 sg13g2_nand2_1 _4574_ (.Y(_0743_),
    .A(_0719_),
    .B(_0742_));
 sg13g2_a21oi_1 _4575_ (.A1(_0726_),
    .A2(_0738_),
    .Y(_0744_),
    .B1(_0737_));
 sg13g2_nor2b_1 _4576_ (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[2] ),
    .Y(_0745_));
 sg13g2_xnor2_1 _4577_ (.Y(_0746_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_nor2b_1 _4578_ (.A(_0744_),
    .B_N(_0746_),
    .Y(_0747_));
 sg13g2_xor2_1 _4579_ (.B(_0746_),
    .A(_0744_),
    .X(_0748_));
 sg13g2_a21oi_1 _4580_ (.A1(_0713_),
    .A2(_0734_),
    .Y(_0749_),
    .B1(net1037));
 sg13g2_a221oi_1 _4581_ (.B2(_0743_),
    .C1(_0681_),
    .B1(_0749_),
    .A1(net1037),
    .Y(_0750_),
    .A2(_0748_));
 sg13g2_a21o_1 _4582_ (.A2(net942),
    .A1(net454),
    .B1(_0750_),
    .X(_0153_));
 sg13g2_nand2_1 _4583_ (.Y(_0751_),
    .A(net516),
    .B(net942));
 sg13g2_o21ai_1 _4584_ (.B1(_0719_),
    .Y(_0752_),
    .A1(_3379_),
    .A2(_0716_));
 sg13g2_o21ai_1 _4585_ (.B1(_0752_),
    .Y(_0753_),
    .A1(net1134),
    .A2(_0721_));
 sg13g2_nand2b_1 _4586_ (.Y(_0754_),
    .B(_0733_),
    .A_N(_0753_));
 sg13g2_inv_1 _4587_ (.Y(_0755_),
    .A(_0754_));
 sg13g2_mux2_1 _4588_ (.A0(_0723_),
    .A1(_0742_),
    .S(_0754_),
    .X(_0756_));
 sg13g2_xnor2_1 _4589_ (.Y(_0757_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_o21ai_1 _4590_ (.B1(_0757_),
    .Y(_0758_),
    .A1(_0745_),
    .A2(_0747_));
 sg13g2_or3_1 _4591_ (.A(_0745_),
    .B(_0747_),
    .C(_0757_),
    .X(_0759_));
 sg13g2_a21oi_1 _4592_ (.A1(_0758_),
    .A2(_0759_),
    .Y(_0760_),
    .B1(_0704_));
 sg13g2_a22oi_1 _4593_ (.Y(_0761_),
    .B1(_0756_),
    .B2(_0736_),
    .A2(_0743_),
    .A1(_0714_));
 sg13g2_nand3_1 _4594_ (.B(net1038),
    .C(_0761_),
    .A(net949),
    .Y(_0762_));
 sg13g2_o21ai_1 _4595_ (.B1(_0751_),
    .Y(_0154_),
    .A1(_0760_),
    .A2(_0762_));
 sg13g2_nand2_1 _4596_ (.Y(_0763_),
    .A(net495),
    .B(net943));
 sg13g2_o21ai_1 _4597_ (.B1(_0758_),
    .Y(_0764_),
    .A1(_3218_),
    .A2(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_nor2b_1 _4598_ (.A(\vgademo.soundtrack.tri_osc_i[7] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[4] ),
    .Y(_0765_));
 sg13g2_xnor2_1 _4599_ (.Y(_0766_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(\vgademo.soundtrack.tri_osc_i[7] ));
 sg13g2_xor2_1 _4600_ (.B(_0766_),
    .A(_0764_),
    .X(_0767_));
 sg13g2_o21ai_1 _4601_ (.B1(_0733_),
    .Y(_0768_),
    .A1(_0723_),
    .A2(_0753_));
 sg13g2_inv_1 _4602_ (.Y(_0769_),
    .A(_0768_));
 sg13g2_a22oi_1 _4603_ (.Y(_0770_),
    .B1(_0769_),
    .B2(_0736_),
    .A2(_0756_),
    .A1(_0714_));
 sg13g2_o21ai_1 _4604_ (.B1(_0770_),
    .Y(_0771_),
    .A1(_0704_),
    .A2(_0767_));
 sg13g2_o21ai_1 _4605_ (.B1(_0763_),
    .Y(_0155_),
    .A1(_0681_),
    .A2(_0771_));
 sg13g2_nor2_1 _4606_ (.A(_0713_),
    .B(_0723_),
    .Y(_0772_));
 sg13g2_a221oi_1 _4607_ (.B2(_0754_),
    .C1(net1037),
    .B1(_0772_),
    .A1(_0713_),
    .Y(_0773_),
    .A2(_0768_));
 sg13g2_a21o_1 _4608_ (.A2(_0766_),
    .A1(_0764_),
    .B1(_0765_),
    .X(_0774_));
 sg13g2_nor2b_1 _4609_ (.A(\vgademo.soundtrack.tri_osc_i[8] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[5] ),
    .Y(_0775_));
 sg13g2_nand2b_1 _4610_ (.Y(_0776_),
    .B(\vgademo.soundtrack.tri_osc_i[8] ),
    .A_N(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_nand2b_1 _4611_ (.Y(_0777_),
    .B(_0776_),
    .A_N(_0775_));
 sg13g2_o21ai_1 _4612_ (.B1(_0705_),
    .Y(_0778_),
    .A1(_0774_),
    .A2(_0777_));
 sg13g2_a21oi_1 _4613_ (.A1(_0774_),
    .A2(_0777_),
    .Y(_0779_),
    .B1(_0778_));
 sg13g2_nor3_1 _4614_ (.A(_0681_),
    .B(_0773_),
    .C(_0779_),
    .Y(_0780_));
 sg13g2_a21o_1 _4615_ (.A2(net943),
    .A1(net568),
    .B1(_0780_),
    .X(_0156_));
 sg13g2_a21oi_1 _4616_ (.A1(_0774_),
    .A2(_0776_),
    .Y(_0781_),
    .B1(_0775_));
 sg13g2_and2_1 _4617_ (.A(_3219_),
    .B(_0781_),
    .X(_0782_));
 sg13g2_xnor2_1 _4618_ (.Y(_0783_),
    .A(_3219_),
    .B(_0781_));
 sg13g2_nand2_1 _4619_ (.Y(_0784_),
    .A(_0713_),
    .B(_0755_));
 sg13g2_nor2_1 _4620_ (.A(net1037),
    .B(_0723_),
    .Y(_0785_));
 sg13g2_a221oi_1 _4621_ (.B2(_0785_),
    .C1(_0681_),
    .B1(_0784_),
    .A1(net1037),
    .Y(_0786_),
    .A2(_0783_));
 sg13g2_a21oi_1 _4622_ (.A1(_3219_),
    .A2(net942),
    .Y(_0157_),
    .B1(_0786_));
 sg13g2_xnor2_1 _4623_ (.Y(_0787_),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .B(_0782_));
 sg13g2_nor2_1 _4624_ (.A(_0704_),
    .B(_0787_),
    .Y(_0788_));
 sg13g2_nor2_1 _4625_ (.A(_0736_),
    .B(_0785_),
    .Y(_0789_));
 sg13g2_nor2_1 _4626_ (.A(_0772_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_nor3_1 _4627_ (.A(_0681_),
    .B(_0788_),
    .C(_0790_),
    .Y(_0791_));
 sg13g2_a21oi_1 _4628_ (.A1(_3220_),
    .A2(net942),
    .Y(_0158_),
    .B1(_0791_));
 sg13g2_a21oi_1 _4629_ (.A1(_3220_),
    .A2(_0782_),
    .Y(_0792_),
    .B1(_3221_));
 sg13g2_o21ai_1 _4630_ (.B1(_0789_),
    .Y(_0793_),
    .A1(_0704_),
    .A2(_0792_));
 sg13g2_nor2b_1 _4631_ (.A(_0681_),
    .B_N(_0793_),
    .Y(_0794_));
 sg13g2_a21oi_1 _4632_ (.A1(_3221_),
    .A2(net942),
    .Y(_0159_),
    .B1(_0794_));
 sg13g2_nor2_1 _4633_ (.A(net1166),
    .B(net248),
    .Y(_0795_));
 sg13g2_a21oi_2 _4634_ (.B1(_0567_),
    .Y(_0796_),
    .A2(_0568_),
    .A1(_0566_));
 sg13g2_a21oi_1 _4635_ (.A1(net1166),
    .A2(_0796_),
    .Y(_0160_),
    .B1(_0795_));
 sg13g2_mux2_1 _4636_ (.A0(\vgademo.soundtrack.tick_div[0] ),
    .A1(net175),
    .S(net980),
    .X(_0161_));
 sg13g2_a21o_1 _4637_ (.A2(net980),
    .A1(\vgademo.soundtrack.tick_div[0] ),
    .B1(net489),
    .X(_0797_));
 sg13g2_and2_1 _4638_ (.A(_0624_),
    .B(net490),
    .X(_0162_));
 sg13g2_xnor2_1 _4639_ (.Y(_0163_),
    .A(net242),
    .B(_0624_));
 sg13g2_xnor2_1 _4640_ (.Y(_0164_),
    .A(net252),
    .B(_0625_));
 sg13g2_xor2_1 _4641_ (.B(_0626_),
    .A(net226),
    .X(_0165_));
 sg13g2_xor2_1 _4642_ (.B(_0627_),
    .A(net264),
    .X(_0166_));
 sg13g2_a21oi_1 _4643_ (.A1(\vgademo.soundtrack.tick_div[5] ),
    .A2(_0627_),
    .Y(_0798_),
    .B1(net199));
 sg13g2_nor2_1 _4644_ (.A(_0628_),
    .B(net200),
    .Y(_0167_));
 sg13g2_xor2_1 _4645_ (.B(_0628_),
    .A(net220),
    .X(_0168_));
 sg13g2_nand2_1 _4646_ (.Y(_0799_),
    .A(_0093_),
    .B(net978));
 sg13g2_o21ai_1 _4647_ (.B1(_0799_),
    .Y(_0169_),
    .A1(net169),
    .A2(net978));
 sg13g2_nand2_1 _4648_ (.Y(_0800_),
    .A(net186),
    .B(net978));
 sg13g2_o21ai_1 _4649_ (.B1(net187),
    .Y(_0170_),
    .A1(\vgademo.soundtrack.noise_lfsr[2] ),
    .A2(net978));
 sg13g2_nand2_1 _4650_ (.Y(_0801_),
    .A(net192),
    .B(net978));
 sg13g2_o21ai_1 _4651_ (.B1(net193),
    .Y(_0171_),
    .A1(\vgademo.soundtrack.noise_lfsr[3] ),
    .A2(net978));
 sg13g2_mux2_1 _4652_ (.A0(net222),
    .A1(_0039_),
    .S(net981),
    .X(_0172_));
 sg13g2_mux2_1 _4653_ (.A0(net240),
    .A1(\vgademo.soundtrack.noise_lfsr[5] ),
    .S(net980),
    .X(_0173_));
 sg13g2_mux2_1 _4654_ (.A0(_0097_),
    .A1(net173),
    .S(net980),
    .X(_0174_));
 sg13g2_mux2_1 _4655_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(net260),
    .S(net980),
    .X(_0175_));
 sg13g2_mux2_1 _4656_ (.A0(_0098_),
    .A1(net177),
    .S(net980),
    .X(_0176_));
 sg13g2_mux2_1 _4657_ (.A0(net330),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net980),
    .X(_0177_));
 sg13g2_mux2_1 _4658_ (.A0(net204),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net979),
    .X(_0178_));
 sg13g2_nand2_1 _4659_ (.Y(_0802_),
    .A(_0099_),
    .B(net979));
 sg13g2_o21ai_1 _4660_ (.B1(_0802_),
    .Y(_0179_),
    .A1(net167),
    .A2(net979));
 sg13g2_nand2_1 _4661_ (.Y(_0803_),
    .A(net196),
    .B(net979));
 sg13g2_o21ai_1 _4662_ (.B1(net197),
    .Y(_0180_),
    .A1(\vgademo.soundtrack.noise_lfsr[12] ),
    .A2(net978));
 sg13g2_mux2_1 _4663_ (.A0(_0101_),
    .A1(net171),
    .S(net981),
    .X(_0181_));
 sg13g2_xor2_1 _4664_ (.B(\vgademo.soundtrack.noise_lfsr[14] ),
    .A(\vgademo.soundtrack.noise_lfsr[0] ),
    .X(_0804_));
 sg13g2_mux2_1 _4665_ (.A0(net244),
    .A1(_0804_),
    .S(net981),
    .X(_0182_));
 sg13g2_mux2_1 _4666_ (.A0(net292),
    .A1(\vgademo.soundtrack.noise_lfsr[14] ),
    .S(net978),
    .X(_0183_));
 sg13g2_nand3_1 _4667_ (.B(_3364_),
    .C(_3379_),
    .A(net1140),
    .Y(_0805_));
 sg13g2_nand3_1 _4668_ (.B(net1133),
    .C(_0805_),
    .A(net1135),
    .Y(_0806_));
 sg13g2_nand2_1 _4669_ (.Y(_0807_),
    .A(net1016),
    .B(_0806_));
 sg13g2_o21ai_1 _4670_ (.B1(_0696_),
    .Y(_0808_),
    .A1(net1150),
    .A2(_3340_));
 sg13g2_o21ai_1 _4671_ (.B1(_0808_),
    .Y(_0809_),
    .A1(net1135),
    .A2(_3352_));
 sg13g2_a22oi_1 _4672_ (.Y(_0810_),
    .B1(_0809_),
    .B2(net1016),
    .A2(_0807_),
    .A1(_0706_));
 sg13g2_nor3_2 _4673_ (.A(net1046),
    .B(_0645_),
    .C(_0647_),
    .Y(_0811_));
 sg13g2_nand4_1 _4674_ (.B(net1133),
    .C(_0805_),
    .A(net1142),
    .Y(_0812_),
    .D(_0811_));
 sg13g2_o21ai_1 _4675_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_3366_),
    .A2(_0810_));
 sg13g2_and2_1 _4676_ (.A(net1039),
    .B(_0813_),
    .X(_0814_));
 sg13g2_a21o_2 _4677_ (.A2(_0684_),
    .A1(net946),
    .B1(_0814_),
    .X(_0815_));
 sg13g2_nand3_1 _4678_ (.B(net1118),
    .C(net1111),
    .A(net1114),
    .Y(_0816_));
 sg13g2_or2_1 _4679_ (.X(_0817_),
    .B(_0816_),
    .A(net1042));
 sg13g2_a21oi_1 _4680_ (.A1(net1118),
    .A2(_0817_),
    .Y(_0818_),
    .B1(net1039));
 sg13g2_nand2_1 _4681_ (.Y(_0819_),
    .A(net183),
    .B(_0815_));
 sg13g2_o21ai_1 _4682_ (.B1(_0819_),
    .Y(_0184_),
    .A1(_0815_),
    .A2(_0818_));
 sg13g2_xnor2_1 _4683_ (.Y(_0820_),
    .A(net1114),
    .B(net1118));
 sg13g2_a21oi_1 _4684_ (.A1(_0817_),
    .A2(_0820_),
    .Y(_0821_),
    .B1(_0631_));
 sg13g2_nand2_1 _4685_ (.Y(_0822_),
    .A(net181),
    .B(_0815_));
 sg13g2_o21ai_1 _4686_ (.B1(_0822_),
    .Y(_0185_),
    .A1(_0815_),
    .A2(_0821_));
 sg13g2_nor2_1 _4687_ (.A(net1107),
    .B(_0816_),
    .Y(_0823_));
 sg13g2_a21oi_1 _4688_ (.A1(net1114),
    .A2(net1118),
    .Y(_0824_),
    .B1(net1111));
 sg13g2_nor4_1 _4689_ (.A(net1039),
    .B(_0684_),
    .C(_0823_),
    .D(_0824_),
    .Y(_0825_));
 sg13g2_a21oi_1 _4690_ (.A1(_3163_),
    .A2(_0815_),
    .Y(_0186_),
    .B1(_0825_));
 sg13g2_a21oi_1 _4691_ (.A1(_3225_),
    .A2(_0816_),
    .Y(_0826_),
    .B1(net1039));
 sg13g2_nand2_1 _4692_ (.Y(_0827_),
    .A(net179),
    .B(_0815_));
 sg13g2_o21ai_1 _4693_ (.B1(_0827_),
    .Y(_0187_),
    .A1(_0815_),
    .A2(_0826_));
 sg13g2_and2_1 _4694_ (.A(net1160),
    .B(net982),
    .X(_0828_));
 sg13g2_nand2_2 _4695_ (.Y(_0829_),
    .A(net1160),
    .B(net982));
 sg13g2_a21oi_1 _4696_ (.A1(_0696_),
    .A2(_0715_),
    .Y(_0830_),
    .B1(\vgademo.audio_beat_out[2] ));
 sg13g2_a22oi_1 _4697_ (.Y(_0831_),
    .B1(_0707_),
    .B2(_3357_),
    .A2(_3364_),
    .A1(_3343_));
 sg13g2_or2_1 _4698_ (.X(_0832_),
    .B(_0831_),
    .A(net1137));
 sg13g2_a21oi_1 _4699_ (.A1(net1141),
    .A2(_0637_),
    .Y(_0833_),
    .B1(_3177_));
 sg13g2_nor2_1 _4700_ (.A(net1046),
    .B(_0833_),
    .Y(_0834_));
 sg13g2_nor3_1 _4701_ (.A(net1142),
    .B(_3378_),
    .C(_0636_),
    .Y(_0835_));
 sg13g2_o21ai_1 _4702_ (.B1(_3345_),
    .Y(_0836_),
    .A1(_3341_),
    .A2(_0835_));
 sg13g2_nor2_1 _4703_ (.A(net1148),
    .B(_0636_),
    .Y(_0837_));
 sg13g2_a21oi_1 _4704_ (.A1(net1140),
    .A2(_3363_),
    .Y(_0838_),
    .B1(_0837_));
 sg13g2_nor2_1 _4705_ (.A(_3352_),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_o21ai_1 _4706_ (.B1(_0836_),
    .Y(_0840_),
    .A1(_3337_),
    .A2(_0839_));
 sg13g2_a21oi_1 _4707_ (.A1(_0832_),
    .A2(_0834_),
    .Y(_0841_),
    .B1(_0840_));
 sg13g2_nand2b_1 _4708_ (.Y(_0842_),
    .B(net1131),
    .A_N(_0841_));
 sg13g2_nand3b_1 _4709_ (.B(net1134),
    .C(_0644_),
    .Y(_0843_),
    .A_N(_0647_));
 sg13g2_nor2b_1 _4710_ (.A(net1131),
    .B_N(_0843_),
    .Y(_0844_));
 sg13g2_o21ai_1 _4711_ (.B1(_3345_),
    .Y(_0845_),
    .A1(_3352_),
    .A2(_0698_));
 sg13g2_o21ai_1 _4712_ (.B1(_3336_),
    .Y(_0846_),
    .A1(net1048),
    .A2(_0707_));
 sg13g2_nand3_1 _4713_ (.B(_0845_),
    .C(_0846_),
    .A(_0844_),
    .Y(_0847_));
 sg13g2_nand3_1 _4714_ (.B(_0842_),
    .C(_0847_),
    .A(net1132),
    .Y(_0848_));
 sg13g2_a21oi_1 _4715_ (.A1(_3360_),
    .A2(_3370_),
    .Y(_0849_),
    .B1(_0638_));
 sg13g2_nor2_1 _4716_ (.A(net1138),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_o21ai_1 _4717_ (.B1(_0639_),
    .Y(_0851_),
    .A1(_3346_),
    .A2(_3374_));
 sg13g2_a21oi_1 _4718_ (.A1(net1138),
    .A2(_0851_),
    .Y(_0852_),
    .B1(_0850_));
 sg13g2_o21ai_1 _4719_ (.B1(_3336_),
    .Y(_0853_),
    .A1(_3170_),
    .A2(net1142));
 sg13g2_nor2_1 _4720_ (.A(_0706_),
    .B(_0853_),
    .Y(_0854_));
 sg13g2_nor2_1 _4721_ (.A(_3383_),
    .B(_0854_),
    .Y(_0855_));
 sg13g2_o21ai_1 _4722_ (.B1(_0855_),
    .Y(_0856_),
    .A1(net1046),
    .A2(_0852_));
 sg13g2_o21ai_1 _4723_ (.B1(net1138),
    .Y(_0857_),
    .A1(_3349_),
    .A2(_0698_));
 sg13g2_nand2b_1 _4724_ (.Y(_0858_),
    .B(_0857_),
    .A_N(_0647_));
 sg13g2_a21oi_1 _4725_ (.A1(net1135),
    .A2(_0858_),
    .Y(_0859_),
    .B1(_3335_));
 sg13g2_a221oi_1 _4726_ (.B2(_0859_),
    .C1(_3176_),
    .B1(_0845_),
    .A1(net1046),
    .Y(_0860_),
    .A2(_3181_));
 sg13g2_a22oi_1 _4727_ (.Y(_0861_),
    .B1(_0856_),
    .B2(_0860_),
    .A2(_0848_),
    .A1(_0830_));
 sg13g2_inv_1 _4728_ (.Y(_0862_),
    .A(net959));
 sg13g2_nor3_1 _4729_ (.A(net1135),
    .B(_3378_),
    .C(_0646_),
    .Y(_0863_));
 sg13g2_a21oi_1 _4730_ (.A1(_3370_),
    .A2(_0863_),
    .Y(_0864_),
    .B1(_3336_));
 sg13g2_nand3_1 _4731_ (.B(_3361_),
    .C(_0699_),
    .A(net1046),
    .Y(_0865_));
 sg13g2_nand3_1 _4732_ (.B(_0859_),
    .C(_0865_),
    .A(_3337_),
    .Y(_0866_));
 sg13g2_nand3b_1 _4733_ (.B(_3347_),
    .C(net1137),
    .Y(_0867_),
    .A_N(_3343_));
 sg13g2_nand3_1 _4734_ (.B(_0849_),
    .C(_0867_),
    .A(net1135),
    .Y(_0868_));
 sg13g2_o21ai_1 _4735_ (.B1(_0868_),
    .Y(_0869_),
    .A1(_0647_),
    .A2(_0864_));
 sg13g2_inv_1 _4736_ (.Y(_0870_),
    .A(_0869_));
 sg13g2_o21ai_1 _4737_ (.B1(_0866_),
    .Y(_0871_),
    .A1(_3383_),
    .A2(_0870_));
 sg13g2_nor2_1 _4738_ (.A(_0839_),
    .B(_0864_),
    .Y(_0872_));
 sg13g2_a21oi_1 _4739_ (.A1(net1144),
    .A2(_3356_),
    .Y(_0873_),
    .B1(_0716_));
 sg13g2_a21oi_1 _4740_ (.A1(net1134),
    .A2(_0873_),
    .Y(_0874_),
    .B1(_0872_));
 sg13g2_nand3_1 _4741_ (.B(_3336_),
    .C(_0708_),
    .A(net1141),
    .Y(_0875_));
 sg13g2_a221oi_1 _4742_ (.B2(_0844_),
    .C1(_3181_),
    .B1(_0875_),
    .A1(net1131),
    .Y(_0876_),
    .A2(_0874_));
 sg13g2_o21ai_1 _4743_ (.B1(_0830_),
    .Y(_0877_),
    .A1(net1132),
    .A2(_3337_));
 sg13g2_nor2_1 _4744_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_a21oi_2 _4745_ (.B1(_0878_),
    .Y(_0879_),
    .A2(_0871_),
    .A1(\vgademo.audio_beat_out[2] ));
 sg13g2_o21ai_1 _4746_ (.B1(_0650_),
    .Y(_0880_),
    .A1(_3181_),
    .A2(_0845_));
 sg13g2_nor4_1 _4747_ (.A(net1046),
    .B(_3383_),
    .C(_0850_),
    .D(_0873_),
    .Y(_0881_));
 sg13g2_a21oi_1 _4748_ (.A1(_3383_),
    .A2(_0880_),
    .Y(_0882_),
    .B1(_0881_));
 sg13g2_nor2_1 _4749_ (.A(net1046),
    .B(_0832_),
    .Y(_0883_));
 sg13g2_a21oi_1 _4750_ (.A1(net1137),
    .A2(_0700_),
    .Y(_0884_),
    .B1(_3383_));
 sg13g2_nand2_1 _4751_ (.Y(_0885_),
    .A(_0836_),
    .B(_0884_));
 sg13g2_o21ai_1 _4752_ (.B1(net1137),
    .Y(_0886_),
    .A1(_3341_),
    .A2(_3343_));
 sg13g2_nor2_1 _4753_ (.A(_3335_),
    .B(_0811_),
    .Y(_0887_));
 sg13g2_a221oi_1 _4754_ (.B2(_0887_),
    .C1(\vgademo.audio_beat_out[2] ),
    .B1(_0886_),
    .A1(_3177_),
    .Y(_0888_),
    .A2(_3181_));
 sg13g2_o21ai_1 _4755_ (.B1(_0888_),
    .Y(_0889_),
    .A1(_0883_),
    .A2(_0885_));
 sg13g2_o21ai_1 _4756_ (.B1(_0889_),
    .Y(_0890_),
    .A1(_3176_),
    .A2(_0882_));
 sg13g2_inv_1 _4757_ (.Y(_0891_),
    .A(_0890_));
 sg13g2_a21oi_2 _4758_ (.B1(net959),
    .Y(_0892_),
    .A2(_0891_),
    .A1(_0879_));
 sg13g2_nand2_1 _4759_ (.Y(_0893_),
    .A(_0879_),
    .B(_0890_));
 sg13g2_nand2_1 _4760_ (.Y(_0894_),
    .A(net959),
    .B(_0893_));
 sg13g2_nand2b_1 _4761_ (.Y(_0895_),
    .B(_0894_),
    .A_N(_0892_));
 sg13g2_nand2_1 _4762_ (.Y(_0896_),
    .A(net964),
    .B(_0895_));
 sg13g2_xnor2_1 _4763_ (.Y(_0188_),
    .A(net270),
    .B(_0896_));
 sg13g2_or2_1 _4764_ (.X(_0897_),
    .B(_0892_),
    .A(_0041_));
 sg13g2_xnor2_1 _4765_ (.Y(_0898_),
    .A(_0041_),
    .B(_0892_));
 sg13g2_inv_1 _4766_ (.Y(_0899_),
    .A(_0898_));
 sg13g2_nand3_1 _4767_ (.B(_0895_),
    .C(_0899_),
    .A(net270),
    .Y(_0900_));
 sg13g2_a21o_1 _4768_ (.A2(_0895_),
    .A1(\vgademo.soundtrack.pulse_osc_p[0] ),
    .B1(_0899_),
    .X(_0901_));
 sg13g2_nand3_1 _4769_ (.B(_0900_),
    .C(_0901_),
    .A(net964),
    .Y(_0902_));
 sg13g2_o21ai_1 _4770_ (.B1(_0902_),
    .Y(_0189_),
    .A1(_3275_),
    .A2(net964));
 sg13g2_nand2b_1 _4771_ (.Y(_0903_),
    .B(_0890_),
    .A_N(_0879_));
 sg13g2_mux2_1 _4772_ (.A0(_0893_),
    .A1(_0903_),
    .S(net959),
    .X(_0904_));
 sg13g2_nor2_1 _4773_ (.A(_3276_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_xnor2_1 _4774_ (.Y(_0906_),
    .A(_3276_),
    .B(_0904_));
 sg13g2_a21oi_1 _4775_ (.A1(_0897_),
    .A2(_0900_),
    .Y(_0907_),
    .B1(_0906_));
 sg13g2_nand3_1 _4776_ (.B(_0900_),
    .C(_0906_),
    .A(_0897_),
    .Y(_0908_));
 sg13g2_nand3b_1 _4777_ (.B(_0908_),
    .C(net964),
    .Y(_0909_),
    .A_N(_0907_));
 sg13g2_o21ai_1 _4778_ (.B1(_0909_),
    .Y(_0190_),
    .A1(_3276_),
    .A2(net964));
 sg13g2_nor2_1 _4779_ (.A(_0879_),
    .B(_0890_),
    .Y(_0910_));
 sg13g2_mux2_1 _4780_ (.A0(_0894_),
    .A1(net959),
    .S(_0910_),
    .X(_0911_));
 sg13g2_nand2_1 _4781_ (.Y(_0912_),
    .A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .B(_0911_));
 sg13g2_xnor2_1 _4782_ (.Y(_0913_),
    .A(_3277_),
    .B(_0911_));
 sg13g2_o21ai_1 _4783_ (.B1(_0913_),
    .Y(_0914_),
    .A1(_0905_),
    .A2(_0907_));
 sg13g2_or3_1 _4784_ (.A(_0905_),
    .B(_0907_),
    .C(_0913_),
    .X(_0915_));
 sg13g2_a21oi_1 _4785_ (.A1(_0914_),
    .A2(_0915_),
    .Y(_0916_),
    .B1(_0829_));
 sg13g2_a21oi_1 _4786_ (.A1(_3277_),
    .A2(_0829_),
    .Y(_0191_),
    .B1(_0916_));
 sg13g2_nor2b_1 _4787_ (.A(_0892_),
    .B_N(_0903_),
    .Y(_0917_));
 sg13g2_and2_1 _4788_ (.A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .B(_0917_),
    .X(_0918_));
 sg13g2_xnor2_1 _4789_ (.Y(_0919_),
    .A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .B(_0917_));
 sg13g2_a21oi_1 _4790_ (.A1(_0912_),
    .A2(_0914_),
    .Y(_0920_),
    .B1(_0919_));
 sg13g2_nand3_1 _4791_ (.B(_0914_),
    .C(_0919_),
    .A(_0912_),
    .Y(_0921_));
 sg13g2_nand2_1 _4792_ (.Y(_0922_),
    .A(net964),
    .B(_0921_));
 sg13g2_nand2_1 _4793_ (.Y(_0923_),
    .A(net316),
    .B(_0829_));
 sg13g2_o21ai_1 _4794_ (.B1(_0923_),
    .Y(_0192_),
    .A1(_0920_),
    .A2(_0922_));
 sg13g2_a21oi_1 _4795_ (.A1(_0862_),
    .A2(_0893_),
    .Y(_0924_),
    .B1(_0910_));
 sg13g2_nand2_1 _4796_ (.Y(_0925_),
    .A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .B(_0924_));
 sg13g2_xnor2_1 _4797_ (.Y(_0926_),
    .A(_3278_),
    .B(_0924_));
 sg13g2_o21ai_1 _4798_ (.B1(_0926_),
    .Y(_0927_),
    .A1(_0918_),
    .A2(_0920_));
 sg13g2_or3_1 _4799_ (.A(_0918_),
    .B(_0920_),
    .C(_0926_),
    .X(_0928_));
 sg13g2_nand3_1 _4800_ (.B(_0927_),
    .C(_0928_),
    .A(net965),
    .Y(_0929_));
 sg13g2_o21ai_1 _4801_ (.B1(_0929_),
    .Y(_0193_),
    .A1(_3278_),
    .A2(net964));
 sg13g2_xnor2_1 _4802_ (.Y(_0930_),
    .A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .B(net959));
 sg13g2_a21oi_1 _4803_ (.A1(_0925_),
    .A2(_0927_),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_and3_1 _4804_ (.X(_0932_),
    .A(_0925_),
    .B(_0927_),
    .C(_0930_));
 sg13g2_nor3_1 _4805_ (.A(_0829_),
    .B(_0931_),
    .C(_0932_),
    .Y(_0933_));
 sg13g2_a21o_1 _4806_ (.A2(_0829_),
    .A1(net345),
    .B1(_0933_),
    .X(_0194_));
 sg13g2_nor2_1 _4807_ (.A(net315),
    .B(net965),
    .Y(_0934_));
 sg13g2_a21o_1 _4808_ (.A2(_0861_),
    .A1(net583),
    .B1(_0931_),
    .X(_0935_));
 sg13g2_nor2_1 _4809_ (.A(_3279_),
    .B(_0861_),
    .Y(_0936_));
 sg13g2_xnor2_1 _4810_ (.Y(_0937_),
    .A(net315),
    .B(net959));
 sg13g2_xnor2_1 _4811_ (.Y(_0938_),
    .A(_0935_),
    .B(_0937_));
 sg13g2_a21oi_1 _4812_ (.A1(net965),
    .A2(_0938_),
    .Y(_0195_),
    .B1(_0934_));
 sg13g2_o21ai_1 _4813_ (.B1(net964),
    .Y(_0939_),
    .A1(_0935_),
    .A2(_0936_));
 sg13g2_a21oi_2 _4814_ (.B1(_0939_),
    .Y(_0940_),
    .A2(net959),
    .A1(_3279_));
 sg13g2_xor2_1 _4815_ (.B(_0940_),
    .A(net267),
    .X(_0196_));
 sg13g2_a21oi_1 _4816_ (.A1(\vgademo.soundtrack.pulse_osc_p[8] ),
    .A2(_0940_),
    .Y(_0941_),
    .B1(net230));
 sg13g2_and3_1 _4817_ (.X(_0942_),
    .A(\vgademo.soundtrack.pulse_osc_p[8] ),
    .B(net230),
    .C(_0940_));
 sg13g2_nor2_1 _4818_ (.A(net231),
    .B(_0942_),
    .Y(_0197_));
 sg13g2_and2_1 _4819_ (.A(net209),
    .B(_0942_),
    .X(_0943_));
 sg13g2_xor2_1 _4820_ (.B(_0942_),
    .A(net209),
    .X(_0198_));
 sg13g2_xor2_1 _4821_ (.B(_0943_),
    .A(net269),
    .X(_0199_));
 sg13g2_nand3_1 _4822_ (.B(net269),
    .C(_0943_),
    .A(net548),
    .Y(_0944_));
 sg13g2_a21o_1 _4823_ (.A2(_0943_),
    .A1(net269),
    .B1(net548),
    .X(_0945_));
 sg13g2_and2_1 _4824_ (.A(_0944_),
    .B(_0945_),
    .X(_0200_));
 sg13g2_xnor2_1 _4825_ (.Y(_0201_),
    .A(net238),
    .B(_0944_));
 sg13g2_nor3_1 _4826_ (.A(\vgademo.audio_kick_frames[0] ),
    .B(net943),
    .C(_0728_),
    .Y(_0946_));
 sg13g2_a21o_1 _4827_ (.A2(_0681_),
    .A1(\vgademo.audio_kick_frames[0] ),
    .B1(_0946_),
    .X(_0202_));
 sg13g2_nand2b_1 _4828_ (.Y(_0947_),
    .B(_0946_),
    .A_N(net460));
 sg13g2_nand3_1 _4829_ (.B(net1039),
    .C(_0702_),
    .A(net949),
    .Y(_0948_));
 sg13g2_o21ai_1 _4830_ (.B1(net460),
    .Y(_0949_),
    .A1(\vgademo.audio_kick_frames[0] ),
    .A2(net943));
 sg13g2_nand3_1 _4831_ (.B(_0948_),
    .C(_0949_),
    .A(_0947_),
    .Y(_0203_));
 sg13g2_o21ai_1 _4832_ (.B1(_0948_),
    .Y(_0950_),
    .A1(net280),
    .A2(_0947_));
 sg13g2_a21o_1 _4833_ (.A2(_0947_),
    .A1(net280),
    .B1(_0950_),
    .X(_0204_));
 sg13g2_nand3_1 _4834_ (.B(_3365_),
    .C(_0642_),
    .A(net1146),
    .Y(_0951_));
 sg13g2_a21oi_1 _4835_ (.A1(net1143),
    .A2(_3378_),
    .Y(_0952_),
    .B1(_0693_));
 sg13g2_nor2_1 _4836_ (.A(_3366_),
    .B(_0641_),
    .Y(_0953_));
 sg13g2_or2_1 _4837_ (.X(_0954_),
    .B(_0953_),
    .A(_0693_));
 sg13g2_nand3_1 _4838_ (.B(_0951_),
    .C(_0952_),
    .A(net1017),
    .Y(_0955_));
 sg13g2_o21ai_1 _4839_ (.B1(_0955_),
    .Y(_0956_),
    .A1(net1017),
    .A2(_0954_));
 sg13g2_o21ai_1 _4840_ (.B1(net1017),
    .Y(_0957_),
    .A1(_3365_),
    .A2(_0711_));
 sg13g2_and3_1 _4841_ (.X(_0958_),
    .A(_3360_),
    .B(_3365_),
    .C(_0699_));
 sg13g2_nand2b_1 _4842_ (.Y(_0959_),
    .B(_0837_),
    .A_N(_3375_));
 sg13g2_o21ai_1 _4843_ (.B1(_0642_),
    .Y(_0960_),
    .A1(_3349_),
    .A2(_0698_));
 sg13g2_o21ai_1 _4844_ (.B1(_0957_),
    .Y(_0961_),
    .A1(net1016),
    .A2(_0805_));
 sg13g2_nor3_1 _4845_ (.A(_0656_),
    .B(_0958_),
    .C(_0961_),
    .Y(_0962_));
 sg13g2_a21oi_1 _4846_ (.A1(_3366_),
    .A2(_0698_),
    .Y(_0963_),
    .B1(net1016));
 sg13g2_a22oi_1 _4847_ (.Y(_0964_),
    .B1(_0963_),
    .B2(_0951_),
    .A2(_0959_),
    .A1(net1016));
 sg13g2_a21o_1 _4848_ (.A2(_0964_),
    .A1(_0656_),
    .B1(_0962_),
    .X(_0965_));
 sg13g2_a21oi_1 _4849_ (.A1(_3350_),
    .A2(_3374_),
    .Y(_0966_),
    .B1(net1016));
 sg13g2_a21oi_1 _4850_ (.A1(net1016),
    .A2(_0960_),
    .Y(_0967_),
    .B1(_0966_));
 sg13g2_nand2_1 _4851_ (.Y(_0968_),
    .A(_0656_),
    .B(_0967_));
 sg13g2_o21ai_1 _4852_ (.B1(_0968_),
    .Y(_0969_),
    .A1(_0656_),
    .A2(_0956_));
 sg13g2_mux2_1 _4853_ (.A0(_0969_),
    .A1(_0965_),
    .S(_0652_),
    .X(_0970_));
 sg13g2_nand2_1 _4854_ (.Y(_0971_),
    .A(_3362_),
    .B(_0811_));
 sg13g2_o21ai_1 _4855_ (.B1(_0971_),
    .Y(_0972_),
    .A1(_0811_),
    .A2(_0954_));
 sg13g2_a21oi_1 _4856_ (.A1(_0655_),
    .A2(_0972_),
    .Y(_0973_),
    .B1(net1038));
 sg13g2_o21ai_1 _4857_ (.B1(_0973_),
    .Y(_0974_),
    .A1(_0655_),
    .A2(_0970_));
 sg13g2_nand2_2 _4858_ (.Y(_0975_),
    .A(_0687_),
    .B(_0974_));
 sg13g2_o21ai_1 _4859_ (.B1(net1038),
    .Y(_0976_),
    .A1(_3222_),
    .A2(_3420_));
 sg13g2_mux2_1 _4860_ (.A0(_0976_),
    .A1(net275),
    .S(_0975_),
    .X(_0205_));
 sg13g2_o21ai_1 _4861_ (.B1(net1038),
    .Y(_0977_),
    .A1(_3420_),
    .A2(_3426_));
 sg13g2_mux2_1 _4862_ (.A0(_0977_),
    .A1(net277),
    .S(_0975_),
    .X(_0206_));
 sg13g2_xor2_1 _4863_ (.B(_3424_),
    .A(net1103),
    .X(_0978_));
 sg13g2_o21ai_1 _4864_ (.B1(net1038),
    .Y(_0979_),
    .A1(_3420_),
    .A2(_0978_));
 sg13g2_mux2_1 _4865_ (.A0(_0979_),
    .A1(net274),
    .S(_0975_),
    .X(_0207_));
 sg13g2_a21oi_1 _4866_ (.A1(\vgademo.soundtrack.pulse_vol[2] ),
    .A2(_3424_),
    .Y(_0980_),
    .B1(net1102));
 sg13g2_nor2_1 _4867_ (.A(_0631_),
    .B(_0980_),
    .Y(_0981_));
 sg13g2_nand2_1 _4868_ (.Y(_0982_),
    .A(net202),
    .B(_0975_));
 sg13g2_o21ai_1 _4869_ (.B1(_0982_),
    .Y(_0208_),
    .A1(_0975_),
    .A2(_0981_));
 sg13g2_nand2_1 _4870_ (.Y(_0983_),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B(net965));
 sg13g2_xnor2_1 _4871_ (.Y(_0209_),
    .A(net246),
    .B(_0983_));
 sg13g2_nand2_1 _4872_ (.Y(_0984_),
    .A(net429),
    .B(net246));
 sg13g2_nand2_1 _4873_ (.Y(_0985_),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .B(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_xor2_1 _4874_ (.B(\vgademo.soundtrack.tri_osc_p[1] ),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(_0986_));
 sg13g2_nand2b_1 _4875_ (.Y(_0987_),
    .B(_0986_),
    .A_N(_0984_));
 sg13g2_xnor2_1 _4876_ (.Y(_0988_),
    .A(_0984_),
    .B(_0986_));
 sg13g2_mux2_1 _4877_ (.A0(net468),
    .A1(_0988_),
    .S(net965),
    .X(_0210_));
 sg13g2_nor2_1 _4878_ (.A(net424),
    .B(net967),
    .Y(_0989_));
 sg13g2_nand2_1 _4879_ (.Y(_0990_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(net424));
 sg13g2_xnor2_1 _4880_ (.Y(_0991_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_a21o_1 _4881_ (.A2(_0987_),
    .A1(_0985_),
    .B1(_0991_),
    .X(_0992_));
 sg13g2_nand3_1 _4882_ (.B(_0987_),
    .C(_0991_),
    .A(_0985_),
    .Y(_0993_));
 sg13g2_nand2_1 _4883_ (.Y(_0994_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_a21oi_1 _4884_ (.A1(net967),
    .A2(_0994_),
    .Y(_0211_),
    .B1(_0989_));
 sg13g2_nor2_1 _4885_ (.A(net431),
    .B(net967),
    .Y(_0995_));
 sg13g2_nand2_1 _4886_ (.Y(_0996_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_xnor2_1 _4887_ (.Y(_0997_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_a21o_1 _4888_ (.A2(_0992_),
    .A1(_0990_),
    .B1(_0997_),
    .X(_0998_));
 sg13g2_nand3_1 _4889_ (.B(_0992_),
    .C(_0997_),
    .A(_0990_),
    .Y(_0999_));
 sg13g2_nand2_1 _4890_ (.Y(_1000_),
    .A(_0998_),
    .B(_0999_));
 sg13g2_a21oi_1 _4891_ (.A1(net967),
    .A2(_1000_),
    .Y(_0212_),
    .B1(_0995_));
 sg13g2_nor2_1 _4892_ (.A(net413),
    .B(net966),
    .Y(_1001_));
 sg13g2_xnor2_1 _4893_ (.Y(_1002_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_a21oi_1 _4894_ (.A1(_0996_),
    .A2(_0998_),
    .Y(_1003_),
    .B1(_1002_));
 sg13g2_nand3_1 _4895_ (.B(_0998_),
    .C(_1002_),
    .A(_0996_),
    .Y(_1004_));
 sg13g2_nand2b_1 _4896_ (.Y(_1005_),
    .B(_1004_),
    .A_N(_1003_));
 sg13g2_a21oi_1 _4897_ (.A1(net966),
    .A2(_1005_),
    .Y(_0213_),
    .B1(_1001_));
 sg13g2_nor2_1 _4898_ (.A(net433),
    .B(net966),
    .Y(_1006_));
 sg13g2_a21o_1 _4899_ (.A2(\vgademo.soundtrack.tri_osc_p[4] ),
    .A1(\vgademo.soundtrack.tri_osc_i[4] ),
    .B1(_1003_),
    .X(_1007_));
 sg13g2_nand2_1 _4900_ (.Y(_1008_),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_xor2_1 _4901_ (.B(\vgademo.soundtrack.tri_osc_p[5] ),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(_1009_));
 sg13g2_xnor2_1 _4902_ (.Y(_1010_),
    .A(_1007_),
    .B(_1009_));
 sg13g2_a21oi_1 _4903_ (.A1(net966),
    .A2(_1010_),
    .Y(_0214_),
    .B1(_1006_));
 sg13g2_nor2_1 _4904_ (.A(_3219_),
    .B(_3272_),
    .Y(_1011_));
 sg13g2_xnor2_1 _4905_ (.Y(_1012_),
    .A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_o21ai_1 _4906_ (.B1(_1007_),
    .Y(_1013_),
    .A1(\vgademo.soundtrack.tri_osc_i[5] ),
    .A2(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_nand3_1 _4907_ (.B(_1012_),
    .C(_1013_),
    .A(_1008_),
    .Y(_1014_));
 sg13g2_a21oi_1 _4908_ (.A1(_1008_),
    .A2(_1013_),
    .Y(_1015_),
    .B1(_1012_));
 sg13g2_nand3b_1 _4909_ (.B(net966),
    .C(_1014_),
    .Y(_1016_),
    .A_N(_1015_));
 sg13g2_o21ai_1 _4910_ (.B1(_1016_),
    .Y(_0215_),
    .A1(_3272_),
    .A2(net966));
 sg13g2_nand2_1 _4911_ (.Y(_1017_),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .B(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_xor2_1 _4912_ (.B(\vgademo.soundtrack.tri_osc_p[7] ),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(_1018_));
 sg13g2_or3_1 _4913_ (.A(_1011_),
    .B(_1015_),
    .C(_1018_),
    .X(_1019_));
 sg13g2_o21ai_1 _4914_ (.B1(_1018_),
    .Y(_1020_),
    .A1(_1011_),
    .A2(_1015_));
 sg13g2_nand3_1 _4915_ (.B(_1019_),
    .C(_1020_),
    .A(net967),
    .Y(_1021_));
 sg13g2_o21ai_1 _4916_ (.B1(_1021_),
    .Y(_0216_),
    .A1(_3271_),
    .A2(net966));
 sg13g2_xnor2_1 _4917_ (.Y(_1022_),
    .A(\vgademo.soundtrack.tri_osc_i[8] ),
    .B(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_and3_1 _4918_ (.X(_1023_),
    .A(_1017_),
    .B(_1020_),
    .C(_1022_));
 sg13g2_a21oi_1 _4919_ (.A1(_1017_),
    .A2(_1020_),
    .Y(_1024_),
    .B1(_1022_));
 sg13g2_nor3_1 _4920_ (.A(_0829_),
    .B(_1023_),
    .C(_1024_),
    .Y(_1025_));
 sg13g2_a21o_1 _4921_ (.A2(_0829_),
    .A1(net428),
    .B1(_1025_),
    .X(_0217_));
 sg13g2_a21oi_1 _4922_ (.A1(\vgademo.soundtrack.tri_osc_i[8] ),
    .A2(\vgademo.soundtrack.tri_osc_p[8] ),
    .Y(_1026_),
    .B1(_1024_));
 sg13g2_and3_1 _4923_ (.X(_1027_),
    .A(_0040_),
    .B(net966),
    .C(_1026_));
 sg13g2_nor2_1 _4924_ (.A(net336),
    .B(net967),
    .Y(_1028_));
 sg13g2_nor3_2 _4925_ (.A(_0040_),
    .B(_0829_),
    .C(_1026_),
    .Y(_1029_));
 sg13g2_nor3_1 _4926_ (.A(_1027_),
    .B(_1028_),
    .C(_1029_),
    .Y(_0218_));
 sg13g2_and2_1 _4927_ (.A(\vgademo.soundtrack.tri_osc_p[10] ),
    .B(_1029_),
    .X(_1030_));
 sg13g2_xor2_1 _4928_ (.B(_1029_),
    .A(net309),
    .X(_0219_));
 sg13g2_and2_1 _4929_ (.A(net294),
    .B(_1030_),
    .X(_1031_));
 sg13g2_xor2_1 _4930_ (.B(_1030_),
    .A(net294),
    .X(_0220_));
 sg13g2_xor2_1 _4931_ (.B(_1031_),
    .A(net333),
    .X(_0221_));
 sg13g2_nand3_1 _4932_ (.B(net333),
    .C(_1031_),
    .A(net399),
    .Y(_1032_));
 sg13g2_a21o_1 _4933_ (.A2(_1031_),
    .A1(net333),
    .B1(net399),
    .X(_1033_));
 sg13g2_and2_1 _4934_ (.A(_1032_),
    .B(_1033_),
    .X(_0222_));
 sg13g2_xnor2_1 _4935_ (.Y(_0223_),
    .A(net366),
    .B(_1032_));
 sg13g2_o21ai_1 _4936_ (.B1(net1100),
    .Y(_1034_),
    .A1(_3270_),
    .A2(_1032_));
 sg13g2_o21ai_1 _4937_ (.B1(_1034_),
    .Y(_0224_),
    .A1(_0551_),
    .A2(_1032_));
 sg13g2_and2_1 _4938_ (.A(net1068),
    .B(net1071),
    .X(_1035_));
 sg13g2_nand2_2 _4939_ (.Y(_1036_),
    .A(net1068),
    .B(net1071));
 sg13g2_nor2_2 _4940_ (.A(net1079),
    .B(net1083),
    .Y(_1037_));
 sg13g2_or2_1 _4941_ (.X(_1038_),
    .B(net1084),
    .A(net1079));
 sg13g2_or2_2 _4942_ (.X(_1039_),
    .B(net1086),
    .A(net1083));
 sg13g2_nor3_1 _4943_ (.A(net1079),
    .B(net1083),
    .C(net1086),
    .Y(_1040_));
 sg13g2_or3_1 _4944_ (.A(net1079),
    .B(net1083),
    .C(net1086),
    .X(_1041_));
 sg13g2_nor2_1 _4945_ (.A(net1045),
    .B(_1040_),
    .Y(_1042_));
 sg13g2_a21oi_2 _4946_ (.B1(net1074),
    .Y(_1043_),
    .A2(_1041_),
    .A1(net1077));
 sg13g2_inv_1 _4947_ (.Y(_1044_),
    .A(_1043_));
 sg13g2_and2_1 _4948_ (.A(net1090),
    .B(_1040_),
    .X(_1045_));
 sg13g2_nand3b_1 _4949_ (.B(_3196_),
    .C(_0065_),
    .Y(_1046_),
    .A_N(net1066));
 sg13g2_nor4_2 _4950_ (.A(net1074),
    .B(net1045),
    .C(_1036_),
    .Y(_1047_),
    .D(_1046_));
 sg13g2_nor2_2 _4951_ (.A(\vgademo.a_scrolly[12] ),
    .B(\vgademo.a_scrolly[13] ),
    .Y(_1048_));
 sg13g2_inv_1 _4952_ (.Y(_1049_),
    .A(_1048_));
 sg13g2_nor3_2 _4953_ (.A(net1066),
    .B(\vgademo.a_scrolly[13] ),
    .C(net1067),
    .Y(_1050_));
 sg13g2_o21ai_1 _4954_ (.B1(_1050_),
    .Y(_1051_),
    .A1(_1036_),
    .A2(_1043_));
 sg13g2_a21oi_2 _4955_ (.B1(_1051_),
    .Y(_1052_),
    .A2(_1047_),
    .A1(_1045_));
 sg13g2_a21o_2 _4956_ (.A2(_1047_),
    .A1(_1045_),
    .B1(_1051_),
    .X(_1053_));
 sg13g2_nor2b_1 _4957_ (.A(net1066),
    .B_N(net1067),
    .Y(_1054_));
 sg13g2_nand2b_2 _4958_ (.Y(_1055_),
    .B(\vgademo.a_scrolly[10] ),
    .A_N(net1072));
 sg13g2_nor2_1 _4959_ (.A(net1075),
    .B(net1077),
    .Y(_1056_));
 sg13g2_nand3_1 _4960_ (.B(net1082),
    .C(net1086),
    .A(net1090),
    .Y(_1057_));
 sg13g2_nand2_1 _4961_ (.Y(_1058_),
    .A(_3200_),
    .B(_1057_));
 sg13g2_a221oi_1 _4962_ (.B2(_1057_),
    .C1(_1055_),
    .B1(_3200_),
    .A1(_3198_),
    .Y(_1059_),
    .A2(net1045));
 sg13g2_o21ai_1 _4963_ (.B1(\vgademo.a_scrolly[10] ),
    .Y(_1060_),
    .A1(net1070),
    .A2(net1075));
 sg13g2_inv_1 _4964_ (.Y(_1061_),
    .A(_1060_));
 sg13g2_o21ai_1 _4965_ (.B1(_1054_),
    .Y(_1062_),
    .A1(_1059_),
    .A2(_1061_));
 sg13g2_a21oi_2 _4966_ (.B1(_0065_),
    .Y(_1063_),
    .A2(_1062_),
    .A1(_0066_));
 sg13g2_nand2_2 _4967_ (.Y(_1064_),
    .A(net1066),
    .B(\vgademo.a_scrolly[13] ));
 sg13g2_inv_1 _4968_ (.Y(_1065_),
    .A(_1064_));
 sg13g2_nor2b_1 _4969_ (.A(_1055_),
    .B_N(net1041),
    .Y(_1066_));
 sg13g2_a21oi_1 _4970_ (.A1(net1069),
    .A2(net1072),
    .Y(_1067_),
    .B1(net1067));
 sg13g2_o21ai_1 _4971_ (.B1(_1067_),
    .Y(_1068_),
    .A1(_1055_),
    .A2(net1041));
 sg13g2_a21oi_2 _4972_ (.B1(_1068_),
    .Y(_1069_),
    .A2(_1066_),
    .A1(_1058_));
 sg13g2_a21o_1 _4973_ (.A2(_1066_),
    .A1(_1058_),
    .B1(_1068_),
    .X(_1070_));
 sg13g2_a221oi_1 _4974_ (.B2(_1070_),
    .C1(_0065_),
    .B1(_1065_),
    .A1(_0066_),
    .Y(_1071_),
    .A2(_1062_));
 sg13g2_nor2_1 _4975_ (.A(net1077),
    .B(net1080),
    .Y(_1072_));
 sg13g2_nand3_1 _4976_ (.B(_1040_),
    .C(net1041),
    .A(net1070),
    .Y(_1073_));
 sg13g2_nand2_1 _4977_ (.Y(_1074_),
    .A(net1067),
    .B(net1068));
 sg13g2_nor2_1 _4978_ (.A(_0064_),
    .B(_1074_),
    .Y(_1075_));
 sg13g2_and4_1 _4979_ (.A(_0065_),
    .B(_1035_),
    .C(_1054_),
    .D(_1056_),
    .X(_1076_));
 sg13g2_a22oi_1 _4980_ (.Y(_1077_),
    .B1(_1076_),
    .B2(_1045_),
    .A2(_1075_),
    .A1(_1073_));
 sg13g2_a221oi_1 _4981_ (.B2(_1045_),
    .C1(_1049_),
    .B1(_1076_),
    .A1(_1073_),
    .Y(_1078_),
    .A2(_1075_));
 sg13g2_o21ai_1 _4982_ (.B1(_1053_),
    .Y(_1079_),
    .A1(_1071_),
    .A2(net1028));
 sg13g2_o21ai_1 _4983_ (.B1(\vgademo.bayer_j[0] ),
    .Y(_1080_),
    .A1(_3202_),
    .A2(net995));
 sg13g2_nor3_1 _4984_ (.A(\vgademo.bayer_j[0] ),
    .B(_3202_),
    .C(net995),
    .Y(_1081_));
 sg13g2_nand3b_1 _4985_ (.B(_3184_),
    .C(_0063_),
    .Y(_1082_),
    .A_N(net995));
 sg13g2_nand2_1 _4986_ (.Y(_1083_),
    .A(_1080_),
    .B(_1082_));
 sg13g2_xor2_1 _4987_ (.B(_1083_),
    .A(\vgademo.audio_kick_frames[0] ),
    .X(_1084_));
 sg13g2_nand2_1 _4988_ (.Y(_1085_),
    .A(net1031),
    .B(_1084_));
 sg13g2_o21ai_1 _4989_ (.B1(_1085_),
    .Y(_0225_),
    .A1(_3203_),
    .A2(_0662_));
 sg13g2_o21ai_1 _4990_ (.B1(_1080_),
    .Y(_1086_),
    .A1(\vgademo.audio_kick_frames[0] ),
    .A2(_1081_));
 sg13g2_nor2_1 _4991_ (.A(net1087),
    .B(net1029),
    .Y(_1087_));
 sg13g2_a21oi_2 _4992_ (.B1(_1087_),
    .Y(_1088_),
    .A2(net1029),
    .A1(_3204_));
 sg13g2_nor2_1 _4993_ (.A(net995),
    .B(_1088_),
    .Y(_1089_));
 sg13g2_xnor2_1 _4994_ (.Y(_1090_),
    .A(\vgademo.bayer_j[1] ),
    .B(_1089_));
 sg13g2_xor2_1 _4995_ (.B(_1090_),
    .A(_0067_),
    .X(_1091_));
 sg13g2_nand2_1 _4996_ (.Y(_1092_),
    .A(_1086_),
    .B(_1091_));
 sg13g2_xor2_1 _4997_ (.B(_1091_),
    .A(_1086_),
    .X(_1093_));
 sg13g2_nand2_1 _4998_ (.Y(_1094_),
    .A(net1031),
    .B(_1093_));
 sg13g2_o21ai_1 _4999_ (.B1(_1094_),
    .Y(_0226_),
    .A1(_3205_),
    .A2(_0662_));
 sg13g2_nor2_1 _5000_ (.A(_0071_),
    .B(_1089_),
    .Y(_1095_));
 sg13g2_a21oi_1 _5001_ (.A1(_0067_),
    .A2(_1090_),
    .Y(_1096_),
    .B1(_1095_));
 sg13g2_nand2_1 _5002_ (.Y(_1097_),
    .A(_3201_),
    .B(net1029));
 sg13g2_xnor2_1 _5003_ (.Y(_1098_),
    .A(net1084),
    .B(_1097_));
 sg13g2_nor2_1 _5004_ (.A(net995),
    .B(_1098_),
    .Y(_1099_));
 sg13g2_xnor2_1 _5005_ (.Y(_1100_),
    .A(_0070_),
    .B(_1099_));
 sg13g2_nand2b_1 _5006_ (.Y(_1101_),
    .B(_1100_),
    .A_N(_1096_));
 sg13g2_xor2_1 _5007_ (.B(_1100_),
    .A(_1096_),
    .X(_1102_));
 sg13g2_xnor2_1 _5008_ (.Y(_1103_),
    .A(_3182_),
    .B(_1102_));
 sg13g2_or2_1 _5009_ (.X(_1104_),
    .B(_1103_),
    .A(_1092_));
 sg13g2_xor2_1 _5010_ (.B(_1103_),
    .A(_1092_),
    .X(_1105_));
 sg13g2_mux2_1 _5011_ (.A0(net286),
    .A1(_1105_),
    .S(net1031),
    .X(_0227_));
 sg13g2_o21ai_1 _5012_ (.B1(_1101_),
    .Y(_1106_),
    .A1(_3182_),
    .A2(_1102_));
 sg13g2_nand2_2 _5013_ (.Y(_1107_),
    .A(net1079),
    .B(_1039_));
 sg13g2_nand2_1 _5014_ (.Y(_1108_),
    .A(_1041_),
    .B(_1107_));
 sg13g2_mux2_2 _5015_ (.A0(_0074_),
    .A1(_1108_),
    .S(net1028),
    .X(_1109_));
 sg13g2_or3_1 _5016_ (.A(_3207_),
    .B(_1079_),
    .C(_1109_),
    .X(_1110_));
 sg13g2_o21ai_1 _5017_ (.B1(_3207_),
    .Y(_1111_),
    .A1(_1079_),
    .A2(_1109_));
 sg13g2_and2_1 _5018_ (.A(_1110_),
    .B(_1111_),
    .X(_1112_));
 sg13g2_nor3_1 _5019_ (.A(net1065),
    .B(net995),
    .C(_1098_),
    .Y(_1113_));
 sg13g2_or3_1 _5020_ (.A(net1065),
    .B(net995),
    .C(_1098_),
    .X(_1114_));
 sg13g2_nor2_1 _5021_ (.A(_1112_),
    .B(_1113_),
    .Y(_1115_));
 sg13g2_xnor2_1 _5022_ (.Y(_1116_),
    .A(_1112_),
    .B(_1114_));
 sg13g2_nand2_1 _5023_ (.Y(_1117_),
    .A(_1106_),
    .B(_1116_));
 sg13g2_xnor2_1 _5024_ (.Y(_1118_),
    .A(_1106_),
    .B(_1116_));
 sg13g2_xor2_1 _5025_ (.B(_1118_),
    .A(_1104_),
    .X(_1119_));
 sg13g2_mux2_1 _5026_ (.A0(net373),
    .A1(_1119_),
    .S(net1031),
    .X(_0228_));
 sg13g2_nor2_1 _5027_ (.A(net285),
    .B(net1030),
    .Y(_1120_));
 sg13g2_o21ai_1 _5028_ (.B1(_1117_),
    .Y(_1121_),
    .A1(_1104_),
    .A2(_1118_));
 sg13g2_a221oi_1 _5029_ (.B2(_1048_),
    .C1(_0065_),
    .B1(_1077_),
    .A1(_0066_),
    .Y(_1122_),
    .A2(_1062_));
 sg13g2_xor2_1 _5030_ (.B(net1080),
    .A(net1078),
    .X(_1123_));
 sg13g2_o21ai_1 _5031_ (.B1(_1123_),
    .Y(_1124_),
    .A1(_1064_),
    .A2(_1069_));
 sg13g2_nand2_1 _5032_ (.Y(_1125_),
    .A(_0068_),
    .B(_1037_));
 sg13g2_xnor2_1 _5033_ (.Y(_1126_),
    .A(_0077_),
    .B(_1125_));
 sg13g2_a221oi_1 _5034_ (.B2(net1028),
    .C1(_1052_),
    .B1(_1126_),
    .A1(_1122_),
    .Y(_1127_),
    .A2(_1124_));
 sg13g2_nand2_1 _5035_ (.Y(_1128_),
    .A(_0076_),
    .B(_1127_));
 sg13g2_xnor2_1 _5036_ (.Y(_1129_),
    .A(_0076_),
    .B(_1127_));
 sg13g2_nand2_1 _5037_ (.Y(_1130_),
    .A(_1110_),
    .B(_1129_));
 sg13g2_xnor2_1 _5038_ (.Y(_1131_),
    .A(_1110_),
    .B(_1129_));
 sg13g2_inv_1 _5039_ (.Y(_1132_),
    .A(_1131_));
 sg13g2_xnor2_1 _5040_ (.Y(_1133_),
    .A(_1115_),
    .B(_1132_));
 sg13g2_nor2b_1 _5041_ (.A(_1133_),
    .B_N(_1121_),
    .Y(_1134_));
 sg13g2_xor2_1 _5042_ (.B(_1133_),
    .A(_1121_),
    .X(_1135_));
 sg13g2_a21oi_1 _5043_ (.A1(net1030),
    .A2(_1135_),
    .Y(_0229_),
    .B1(_1120_));
 sg13g2_a21oi_1 _5044_ (.A1(_1115_),
    .A2(_1132_),
    .Y(_1136_),
    .B1(_1134_));
 sg13g2_xor2_1 _5045_ (.B(_1072_),
    .A(_0079_),
    .X(_1137_));
 sg13g2_o21ai_1 _5046_ (.B1(_1137_),
    .Y(_1138_),
    .A1(_1064_),
    .A2(_1069_));
 sg13g2_nand2_1 _5047_ (.Y(_1139_),
    .A(net1078),
    .B(_1125_));
 sg13g2_xor2_1 _5048_ (.B(_1139_),
    .A(_0079_),
    .X(_1140_));
 sg13g2_a22oi_1 _5049_ (.Y(_1141_),
    .B1(_1140_),
    .B2(net1028),
    .A2(_1138_),
    .A1(_1122_));
 sg13g2_nor3_1 _5050_ (.A(_3185_),
    .B(_1052_),
    .C(_1141_),
    .Y(_1142_));
 sg13g2_o21ai_1 _5051_ (.B1(_3185_),
    .Y(_1143_),
    .A1(_1052_),
    .A2(_1141_));
 sg13g2_nand2b_1 _5052_ (.Y(_1144_),
    .B(_1143_),
    .A_N(_1142_));
 sg13g2_nor2_1 _5053_ (.A(_1128_),
    .B(_1144_),
    .Y(_1145_));
 sg13g2_xor2_1 _5054_ (.B(_1144_),
    .A(_1128_),
    .X(_1146_));
 sg13g2_xor2_1 _5055_ (.B(_1146_),
    .A(_1130_),
    .X(_1147_));
 sg13g2_nand2b_1 _5056_ (.Y(_1148_),
    .B(_1147_),
    .A_N(_1136_));
 sg13g2_xnor2_1 _5057_ (.Y(_1149_),
    .A(_1136_),
    .B(_1147_));
 sg13g2_mux2_1 _5058_ (.A0(net410),
    .A1(_1149_),
    .S(net1030),
    .X(_0230_));
 sg13g2_nor2_1 _5059_ (.A(net279),
    .B(net1030),
    .Y(_1150_));
 sg13g2_o21ai_1 _5060_ (.B1(_1148_),
    .Y(_1151_),
    .A1(_1130_),
    .A2(_1146_));
 sg13g2_o21ai_1 _5061_ (.B1(_0062_),
    .Y(_1152_),
    .A1(_1052_),
    .A2(_1141_));
 sg13g2_nand2_1 _5062_ (.Y(_1153_),
    .A(net1074),
    .B(net1077));
 sg13g2_a21oi_2 _5063_ (.B1(_1153_),
    .Y(_1154_),
    .A2(_1037_),
    .A1(_0068_));
 sg13g2_nor2_1 _5064_ (.A(net1071),
    .B(_1154_),
    .Y(_1155_));
 sg13g2_xnor2_1 _5065_ (.Y(_1156_),
    .A(net1071),
    .B(_1154_));
 sg13g2_and2_1 _5066_ (.A(net1028),
    .B(_1156_),
    .X(_1157_));
 sg13g2_nand2_1 _5067_ (.Y(_1158_),
    .A(_0074_),
    .B(net1041));
 sg13g2_nand3b_1 _5068_ (.B(_0074_),
    .C(net1041),
    .Y(_1159_),
    .A_N(net1070));
 sg13g2_xor2_1 _5069_ (.B(_1158_),
    .A(net1073),
    .X(_1160_));
 sg13g2_o21ai_1 _5070_ (.B1(_1160_),
    .Y(_1161_),
    .A1(_1064_),
    .A2(_1069_));
 sg13g2_a21o_1 _5071_ (.A2(_1161_),
    .A1(_1122_),
    .B1(_1157_),
    .X(_1162_));
 sg13g2_and3_1 _5072_ (.X(_1163_),
    .A(\vgademo.v_count[6] ),
    .B(_1053_),
    .C(_1162_));
 sg13g2_a21oi_1 _5073_ (.A1(_1053_),
    .A2(_1162_),
    .Y(_1164_),
    .B1(net1061));
 sg13g2_or2_1 _5074_ (.X(_1165_),
    .B(_1164_),
    .A(_1163_));
 sg13g2_nand2_1 _5075_ (.Y(_1166_),
    .A(_1152_),
    .B(_1165_));
 sg13g2_xnor2_1 _5076_ (.Y(_1167_),
    .A(_1152_),
    .B(_1165_));
 sg13g2_nor2_1 _5077_ (.A(_1145_),
    .B(_1167_),
    .Y(_1168_));
 sg13g2_xor2_1 _5078_ (.B(_1167_),
    .A(_1145_),
    .X(_1169_));
 sg13g2_xnor2_1 _5079_ (.Y(_1170_),
    .A(_1151_),
    .B(_1169_));
 sg13g2_a21oi_1 _5080_ (.A1(net1031),
    .A2(_1170_),
    .Y(_0231_),
    .B1(_1150_));
 sg13g2_a21oi_1 _5081_ (.A1(_1151_),
    .A2(_1169_),
    .Y(_1171_),
    .B1(_1168_));
 sg13g2_inv_1 _5082_ (.Y(_1172_),
    .A(_1171_));
 sg13g2_xor2_1 _5083_ (.B(_1159_),
    .A(_0015_),
    .X(_1173_));
 sg13g2_o21ai_1 _5084_ (.B1(_1173_),
    .Y(_1174_),
    .A1(_1064_),
    .A2(_1069_));
 sg13g2_a21o_2 _5085_ (.A2(_1174_),
    .A1(_1063_),
    .B1(net1028),
    .X(_1175_));
 sg13g2_nor2b_1 _5086_ (.A(_1154_),
    .B_N(_0064_),
    .Y(_1176_));
 sg13g2_xnor2_1 _5087_ (.Y(_1177_),
    .A(_3197_),
    .B(_1176_));
 sg13g2_a21oi_2 _5088_ (.B1(_1052_),
    .Y(_1178_),
    .A2(_1177_),
    .A1(net1029));
 sg13g2_a21oi_2 _5089_ (.B1(_3209_),
    .Y(_1179_),
    .A2(_1178_),
    .A1(_1175_));
 sg13g2_and3_1 _5090_ (.X(_1180_),
    .A(_3209_),
    .B(_1175_),
    .C(_1178_));
 sg13g2_nor2_1 _5091_ (.A(_1179_),
    .B(_1180_),
    .Y(_1181_));
 sg13g2_a21oi_2 _5092_ (.B1(_3210_),
    .Y(_1182_),
    .A2(_1162_),
    .A1(_1053_));
 sg13g2_nor2_1 _5093_ (.A(_1181_),
    .B(_1182_),
    .Y(_1183_));
 sg13g2_xor2_1 _5094_ (.B(_1182_),
    .A(_1181_),
    .X(_1184_));
 sg13g2_nor2b_1 _5095_ (.A(_1166_),
    .B_N(_1184_),
    .Y(_1185_));
 sg13g2_xnor2_1 _5096_ (.Y(_1186_),
    .A(_1166_),
    .B(_1184_));
 sg13g2_xnor2_1 _5097_ (.Y(_1187_),
    .A(_1171_),
    .B(_1186_));
 sg13g2_mux2_1 _5098_ (.A0(net296),
    .A1(_1187_),
    .S(net1031),
    .X(_0232_));
 sg13g2_a21oi_1 _5099_ (.A1(_1172_),
    .A2(_1186_),
    .Y(_1188_),
    .B1(_1185_));
 sg13g2_nand3b_1 _5100_ (.B(net1041),
    .C(_3200_),
    .Y(_1189_),
    .A_N(_1055_));
 sg13g2_a21oi_1 _5101_ (.A1(net1069),
    .A2(_1189_),
    .Y(_1190_),
    .B1(_3212_));
 sg13g2_and3_1 _5102_ (.X(_1191_),
    .A(net1069),
    .B(_3212_),
    .C(_1189_));
 sg13g2_nor3_1 _5103_ (.A(net1028),
    .B(_1190_),
    .C(_1191_),
    .Y(_1192_));
 sg13g2_or2_1 _5104_ (.X(_1193_),
    .B(_1155_),
    .A(_1074_));
 sg13g2_a22oi_1 _5105_ (.Y(_1194_),
    .B1(_1193_),
    .B2(net1028),
    .A2(_1192_),
    .A1(_1071_));
 sg13g2_xnor2_1 _5106_ (.Y(_1195_),
    .A(_3213_),
    .B(_1194_));
 sg13g2_xnor2_1 _5107_ (.Y(_1196_),
    .A(_1179_),
    .B(_1195_));
 sg13g2_xnor2_1 _5108_ (.Y(_1197_),
    .A(_1183_),
    .B(_1196_));
 sg13g2_xor2_1 _5109_ (.B(_1197_),
    .A(_1188_),
    .X(_1198_));
 sg13g2_nand2_1 _5110_ (.Y(_1199_),
    .A(_0662_),
    .B(_1198_));
 sg13g2_o21ai_1 _5111_ (.B1(_1199_),
    .Y(_0233_),
    .A1(_3214_),
    .A2(_0661_));
 sg13g2_nor2_2 _5112_ (.A(net1068),
    .B(net1070),
    .Y(_1200_));
 sg13g2_nand2_1 _5113_ (.Y(_1201_),
    .A(net1090),
    .B(net1079));
 sg13g2_nand3_1 _5114_ (.B(_1200_),
    .C(_1201_),
    .A(net1041),
    .Y(_1202_));
 sg13g2_nand2b_1 _5115_ (.Y(_1203_),
    .B(_1107_),
    .A_N(_1046_));
 sg13g2_nor2_1 _5116_ (.A(net1090),
    .B(net1086),
    .Y(_1204_));
 sg13g2_nand3b_1 _5117_ (.B(_3343_),
    .C(_3349_),
    .Y(_1205_),
    .A_N(net1131));
 sg13g2_nor3_2 _5118_ (.A(net1132),
    .B(_3337_),
    .C(_1205_),
    .Y(_1206_));
 sg13g2_o21ai_1 _5119_ (.B1(_1206_),
    .Y(_1207_),
    .A1(_1202_),
    .A2(_1203_));
 sg13g2_nand2_1 _5120_ (.Y(_1208_),
    .A(_0593_),
    .B(_1207_));
 sg13g2_nand2_1 _5121_ (.Y(_1209_),
    .A(net1088),
    .B(net1020));
 sg13g2_o21ai_1 _5122_ (.B1(_1209_),
    .Y(_0234_),
    .A1(net1088),
    .A2(net994));
 sg13g2_nand2_1 _5123_ (.Y(_1210_),
    .A(net1086),
    .B(net1018));
 sg13g2_xnor2_1 _5124_ (.Y(_1211_),
    .A(net1090),
    .B(net1086));
 sg13g2_o21ai_1 _5125_ (.B1(_1210_),
    .Y(_0235_),
    .A1(net994),
    .A2(_1211_));
 sg13g2_nand2_1 _5126_ (.Y(_1212_),
    .A(net1082),
    .B(net1020));
 sg13g2_a21o_1 _5127_ (.A2(net1085),
    .A1(net1089),
    .B1(net1082),
    .X(_1213_));
 sg13g2_nand2_1 _5128_ (.Y(_1214_),
    .A(_1057_),
    .B(_1213_));
 sg13g2_o21ai_1 _5129_ (.B1(_1212_),
    .Y(_0236_),
    .A1(_1208_),
    .A2(_1214_));
 sg13g2_nand2_1 _5130_ (.Y(_1215_),
    .A(net1080),
    .B(net1018));
 sg13g2_xnor2_1 _5131_ (.Y(_1216_),
    .A(net580),
    .B(_1057_));
 sg13g2_o21ai_1 _5132_ (.B1(_1215_),
    .Y(_0237_),
    .A1(_1208_),
    .A2(_1216_));
 sg13g2_nand2_1 _5133_ (.Y(_1217_),
    .A(net1077),
    .B(net1018));
 sg13g2_nand2_1 _5134_ (.Y(_1218_),
    .A(net1079),
    .B(net1083));
 sg13g2_inv_1 _5135_ (.Y(_1219_),
    .A(_1218_));
 sg13g2_or2_1 _5136_ (.X(_1220_),
    .B(_1057_),
    .A(_3200_));
 sg13g2_nor2_1 _5137_ (.A(_0077_),
    .B(_1220_),
    .Y(_1221_));
 sg13g2_xnor2_1 _5138_ (.Y(_1222_),
    .A(_0077_),
    .B(_1220_));
 sg13g2_o21ai_1 _5139_ (.B1(_1217_),
    .Y(_0238_),
    .A1(net994),
    .A2(_1222_));
 sg13g2_nand2_1 _5140_ (.Y(_1223_),
    .A(net1074),
    .B(net1018));
 sg13g2_xor2_1 _5141_ (.B(_1221_),
    .A(net577),
    .X(_1224_));
 sg13g2_o21ai_1 _5142_ (.B1(_1223_),
    .Y(_0239_),
    .A1(net994),
    .A2(_1224_));
 sg13g2_nand2_1 _5143_ (.Y(_1225_),
    .A(net1071),
    .B(net1018));
 sg13g2_or2_1 _5144_ (.X(_1226_),
    .B(_1220_),
    .A(_1153_));
 sg13g2_nor2_1 _5145_ (.A(_0064_),
    .B(_1226_),
    .Y(_1227_));
 sg13g2_xnor2_1 _5146_ (.Y(_1228_),
    .A(net492),
    .B(_1226_));
 sg13g2_o21ai_1 _5147_ (.B1(_1225_),
    .Y(_0240_),
    .A1(net994),
    .A2(_1228_));
 sg13g2_nand2_1 _5148_ (.Y(_1229_),
    .A(net1068),
    .B(net1018));
 sg13g2_xor2_1 _5149_ (.B(_1227_),
    .A(net470),
    .X(_1230_));
 sg13g2_o21ai_1 _5150_ (.B1(_1229_),
    .Y(_0241_),
    .A1(net994),
    .A2(net471));
 sg13g2_nor2_1 _5151_ (.A(_1036_),
    .B(_1226_),
    .Y(_1231_));
 sg13g2_nor3_1 _5152_ (.A(_0019_),
    .B(_1036_),
    .C(_1226_),
    .Y(_1232_));
 sg13g2_xnor2_1 _5153_ (.Y(_1233_),
    .A(net571),
    .B(_1231_));
 sg13g2_nand3_1 _5154_ (.B(_1207_),
    .C(_1233_),
    .A(net999),
    .Y(_1234_));
 sg13g2_o21ai_1 _5155_ (.B1(_1234_),
    .Y(_0242_),
    .A1(_3196_),
    .A2(net999));
 sg13g2_nand2_1 _5156_ (.Y(_1235_),
    .A(net1066),
    .B(net1018));
 sg13g2_xor2_1 _5157_ (.B(_1232_),
    .A(_0066_),
    .X(_1236_));
 sg13g2_o21ai_1 _5158_ (.B1(_1235_),
    .Y(_0243_),
    .A1(net994),
    .A2(_1236_));
 sg13g2_nand2_1 _5159_ (.Y(_1237_),
    .A(net554),
    .B(net1018));
 sg13g2_nand3_1 _5160_ (.B(\vgademo.a_scrolly[11] ),
    .C(_1231_),
    .A(net1066),
    .Y(_1238_));
 sg13g2_xnor2_1 _5161_ (.Y(_1239_),
    .A(_0065_),
    .B(_1238_));
 sg13g2_o21ai_1 _5162_ (.B1(_1237_),
    .Y(_0244_),
    .A1(net994),
    .A2(_1239_));
 sg13g2_nor2_2 _5163_ (.A(net1033),
    .B(_0592_),
    .Y(_1240_));
 sg13g2_nand2_2 _5164_ (.Y(_1241_),
    .A(net1036),
    .B(_0590_));
 sg13g2_nor2_1 _5165_ (.A(net582),
    .B(_1240_),
    .Y(_1242_));
 sg13g2_nand2_1 _5166_ (.Y(_1243_),
    .A(\vgademo.bayer_j[0] ),
    .B(net1036));
 sg13g2_nor2b_1 _5167_ (.A(_1242_),
    .B_N(_1243_),
    .Y(_0245_));
 sg13g2_xnor2_1 _5168_ (.Y(_0246_),
    .A(net476),
    .B(_1243_));
 sg13g2_nand2_1 _5169_ (.Y(_1244_),
    .A(net256),
    .B(net1034));
 sg13g2_nand2_2 _5170_ (.Y(_1245_),
    .A(\vgademo.bayer_j[1] ),
    .B(\vgademo.bayer_j[0] ));
 sg13g2_nor2_1 _5171_ (.A(_0070_),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_xnor2_1 _5172_ (.Y(_1247_),
    .A(_0070_),
    .B(_1245_));
 sg13g2_o21ai_1 _5173_ (.B1(_1244_),
    .Y(_0247_),
    .A1(_1241_),
    .A2(_1247_));
 sg13g2_nand2_1 _5174_ (.Y(_1248_),
    .A(net1064),
    .B(net1034));
 sg13g2_xnor2_1 _5175_ (.Y(_1249_),
    .A(_3207_),
    .B(_1246_));
 sg13g2_o21ai_1 _5176_ (.B1(_1248_),
    .Y(_0248_),
    .A1(_1241_),
    .A2(net456));
 sg13g2_nand2_1 _5177_ (.Y(_1250_),
    .A(net1063),
    .B(net1033));
 sg13g2_nor2_1 _5178_ (.A(_0588_),
    .B(_1245_),
    .Y(_1251_));
 sg13g2_nor3_1 _5179_ (.A(_0076_),
    .B(_0588_),
    .C(_1245_),
    .Y(_1252_));
 sg13g2_xor2_1 _5180_ (.B(_1251_),
    .A(_0076_),
    .X(_1253_));
 sg13g2_o21ai_1 _5181_ (.B1(_1250_),
    .Y(_0249_),
    .A1(_1241_),
    .A2(_1253_));
 sg13g2_nand2_1 _5182_ (.Y(_1254_),
    .A(net503),
    .B(net1033));
 sg13g2_xor2_1 _5183_ (.B(_1252_),
    .A(_0062_),
    .X(_1255_));
 sg13g2_o21ai_1 _5184_ (.B1(_1254_),
    .Y(_0250_),
    .A1(_1241_),
    .A2(_1255_));
 sg13g2_nand3_1 _5185_ (.B(\vgademo.v_count[5] ),
    .C(_1251_),
    .A(net1062),
    .Y(_1256_));
 sg13g2_nor2_1 _5186_ (.A(_0016_),
    .B(_1256_),
    .Y(_1257_));
 sg13g2_nand2_1 _5187_ (.Y(_1258_),
    .A(net565),
    .B(_1256_));
 sg13g2_nand3b_1 _5188_ (.B(_1258_),
    .C(_1240_),
    .Y(_1259_),
    .A_N(_1257_));
 sg13g2_o21ai_1 _5189_ (.B1(_1259_),
    .Y(_0251_),
    .A1(_3186_),
    .A2(net1036));
 sg13g2_xnor2_1 _5190_ (.Y(_1260_),
    .A(net380),
    .B(_1257_));
 sg13g2_a22oi_1 _5191_ (.Y(_1261_),
    .B1(_1240_),
    .B2(_1260_),
    .A2(net1033),
    .A1(net1060));
 sg13g2_inv_1 _5192_ (.Y(_0252_),
    .A(net381));
 sg13g2_or2_1 _5193_ (.X(_1262_),
    .B(_1256_),
    .A(_3313_));
 sg13g2_nand2_1 _5194_ (.Y(_1263_),
    .A(net452),
    .B(_1262_));
 sg13g2_nand2b_1 _5195_ (.Y(_1264_),
    .B(_3213_),
    .A_N(_1262_));
 sg13g2_nand3_1 _5196_ (.B(_1263_),
    .C(_1264_),
    .A(_1240_),
    .Y(_1265_));
 sg13g2_o21ai_1 _5197_ (.B1(_1265_),
    .Y(_0253_),
    .A1(_3187_),
    .A2(net1036));
 sg13g2_nand2_1 _5198_ (.Y(_1266_),
    .A(net1059),
    .B(net1033));
 sg13g2_xnor2_1 _5199_ (.Y(_1267_),
    .A(net340),
    .B(_1264_));
 sg13g2_o21ai_1 _5200_ (.B1(_1266_),
    .Y(_0254_),
    .A1(_1241_),
    .A2(_1267_));
 sg13g2_nand2_1 _5201_ (.Y(_1268_),
    .A(\vgademo.h_count[5] ),
    .B(_3280_));
 sg13g2_xnor2_1 _5202_ (.Y(_1269_),
    .A(\vgademo.h_count[6] ),
    .B(\vgademo.scanline_audio_sample[6] ));
 sg13g2_nand3_1 _5203_ (.B(_1268_),
    .C(_1269_),
    .A(_0036_),
    .Y(_1270_));
 sg13g2_nor2_1 _5204_ (.A(_3193_),
    .B(\vgademo.scanline_audio_sample[4] ),
    .Y(_1271_));
 sg13g2_nand2_1 _5205_ (.Y(_1272_),
    .A(_3193_),
    .B(\vgademo.scanline_audio_sample[4] ));
 sg13g2_o21ai_1 _5206_ (.B1(_1272_),
    .Y(_1273_),
    .A1(\vgademo.h_count[5] ),
    .A2(_3280_));
 sg13g2_nor3_1 _5207_ (.A(_1270_),
    .B(_1271_),
    .C(_1273_),
    .Y(_1274_));
 sg13g2_nand2_1 _5208_ (.Y(_1275_),
    .A(_3191_),
    .B(\vgademo.scanline_audio_sample[2] ));
 sg13g2_xor2_1 _5209_ (.B(\vgademo.scanline_audio_sample[2] ),
    .A(net1095),
    .X(_1276_));
 sg13g2_inv_1 _5210_ (.Y(_1277_),
    .A(_1276_));
 sg13g2_nand2_1 _5211_ (.Y(_1278_),
    .A(net1093),
    .B(_3281_));
 sg13g2_xnor2_1 _5212_ (.Y(_1279_),
    .A(net1093),
    .B(\vgademo.scanline_audio_sample[3] ));
 sg13g2_nand3_1 _5213_ (.B(_1277_),
    .C(_1279_),
    .A(_1274_),
    .Y(_1280_));
 sg13g2_xor2_1 _5214_ (.B(\vgademo.scanline_audio_sample[1] ),
    .A(net1096),
    .X(_1281_));
 sg13g2_a21oi_1 _5215_ (.A1(net1098),
    .A2(_3282_),
    .Y(_1282_),
    .B1(_1281_));
 sg13g2_a21o_1 _5216_ (.A2(\vgademo.scanline_audio_sample[1] ),
    .A1(_3188_),
    .B1(_1282_),
    .X(_1283_));
 sg13g2_nand2b_1 _5217_ (.Y(_1284_),
    .B(_1283_),
    .A_N(_1280_));
 sg13g2_nor2b_1 _5218_ (.A(_1270_),
    .B_N(_1273_),
    .Y(_1285_));
 sg13g2_nor2_1 _5219_ (.A(\vgademo.h_count[7] ),
    .B(\vgademo.h_count[6] ),
    .Y(_1286_));
 sg13g2_a21oi_1 _5220_ (.A1(\vgademo.scanline_audio_sample[6] ),
    .A2(_1286_),
    .Y(_1287_),
    .B1(_1285_));
 sg13g2_o21ai_1 _5221_ (.B1(_1275_),
    .Y(_1288_),
    .A1(net1093),
    .A2(_3281_));
 sg13g2_nand3_1 _5222_ (.B(_1278_),
    .C(_1288_),
    .A(_1274_),
    .Y(_1289_));
 sg13g2_nand3_1 _5223_ (.B(_1287_),
    .C(_1289_),
    .A(_1284_),
    .Y(_1290_));
 sg13g2_o21ai_1 _5224_ (.B1(_1282_),
    .Y(_1291_),
    .A1(net1098),
    .A2(_3282_));
 sg13g2_nor2_1 _5225_ (.A(_1280_),
    .B(_1291_),
    .Y(_1292_));
 sg13g2_nand2_1 _5226_ (.Y(_1293_),
    .A(net1092),
    .B(_3319_));
 sg13g2_nor2_2 _5227_ (.A(_1292_),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_and2_1 _5228_ (.A(_1290_),
    .B(_1294_),
    .X(_1295_));
 sg13g2_nand2_1 _5229_ (.Y(_1296_),
    .A(_1290_),
    .B(_1294_));
 sg13g2_nor2_1 _5230_ (.A(\vgademo.scanline_audio_sample[3] ),
    .B(\vgademo.scanline_audio_sample[4] ),
    .Y(_1297_));
 sg13g2_nand2_1 _5231_ (.Y(_1298_),
    .A(_0042_),
    .B(_1297_));
 sg13g2_xor2_1 _5232_ (.B(_1298_),
    .A(\vgademo.scanline_audio_sample[6] ),
    .X(_1299_));
 sg13g2_xnor2_1 _5233_ (.Y(_1300_),
    .A(_0035_),
    .B(_1299_));
 sg13g2_xnor2_1 _5234_ (.Y(_1301_),
    .A(_0042_),
    .B(_1297_));
 sg13g2_xor2_1 _5235_ (.B(_1301_),
    .A(_0034_),
    .X(_1302_));
 sg13g2_xor2_1 _5236_ (.B(\vgademo.scanline_audio_sample[4] ),
    .A(\vgademo.scanline_audio_sample[3] ),
    .X(_1303_));
 sg13g2_nor2b_1 _5237_ (.A(_1303_),
    .B_N(_0043_),
    .Y(_1304_));
 sg13g2_xnor2_1 _5238_ (.Y(_1305_),
    .A(_0043_),
    .B(_1303_));
 sg13g2_nand4_1 _5239_ (.B(_1300_),
    .C(_1302_),
    .A(_0036_),
    .Y(_1306_),
    .D(_1305_));
 sg13g2_nor2_1 _5240_ (.A(_1276_),
    .B(_1279_),
    .Y(_1307_));
 sg13g2_nor2_1 _5241_ (.A(_1275_),
    .B(_1279_),
    .Y(_1308_));
 sg13g2_a221oi_1 _5242_ (.B2(_1307_),
    .C1(_1308_),
    .B1(_1283_),
    .A1(_3190_),
    .Y(_1309_),
    .A2(_3281_));
 sg13g2_nor2b_1 _5243_ (.A(_1299_),
    .B_N(_1286_),
    .Y(_1310_));
 sg13g2_a22oi_1 _5244_ (.Y(_1311_),
    .B1(_1302_),
    .B2(_1304_),
    .A2(_1301_),
    .A1(_3192_));
 sg13g2_nand3b_1 _5245_ (.B(_1300_),
    .C(_0036_),
    .Y(_1312_),
    .A_N(_1311_));
 sg13g2_o21ai_1 _5246_ (.B1(_1312_),
    .Y(_1313_),
    .A1(_1306_),
    .A2(_1309_));
 sg13g2_nor2_1 _5247_ (.A(_1291_),
    .B(_1306_),
    .Y(_1314_));
 sg13g2_a21oi_1 _5248_ (.A1(_1307_),
    .A2(_1314_),
    .Y(_1315_),
    .B1(_1293_));
 sg13g2_o21ai_1 _5249_ (.B1(_1315_),
    .Y(_1316_),
    .A1(_1310_),
    .A2(_1313_));
 sg13g2_nor2_2 _5250_ (.A(net961),
    .B(_1316_),
    .Y(_1317_));
 sg13g2_or2_2 _5251_ (.X(_1318_),
    .B(_1316_),
    .A(net961));
 sg13g2_nor4_2 _5252_ (.A(_1163_),
    .B(_1164_),
    .C(_1179_),
    .Y(_1319_),
    .D(_1180_));
 sg13g2_or2_1 _5253_ (.X(_1320_),
    .B(_1195_),
    .A(net1059));
 sg13g2_nor3_1 _5254_ (.A(net1059),
    .B(_1129_),
    .C(_1195_),
    .Y(_1321_));
 sg13g2_nand3b_1 _5255_ (.B(_1319_),
    .C(_1321_),
    .Y(_1322_),
    .A_N(_1144_));
 sg13g2_o21ai_1 _5256_ (.B1(net1065),
    .Y(_1323_),
    .A1(net995),
    .A2(_1098_));
 sg13g2_and4_1 _5257_ (.A(_1110_),
    .B(_1111_),
    .C(_1114_),
    .D(_1323_),
    .X(_1324_));
 sg13g2_and2_1 _5258_ (.A(_0071_),
    .B(_1089_),
    .X(_1325_));
 sg13g2_nand2_1 _5259_ (.Y(_1326_),
    .A(_1090_),
    .B(_1324_));
 sg13g2_nand3_1 _5260_ (.B(_1090_),
    .C(_1324_),
    .A(_1080_),
    .Y(_1327_));
 sg13g2_nor3_1 _5261_ (.A(\vgademo.v_count[3] ),
    .B(_1079_),
    .C(_1109_),
    .Y(_1328_));
 sg13g2_a221oi_1 _5262_ (.B2(_1325_),
    .C1(_1328_),
    .B1(_1324_),
    .A1(_1112_),
    .Y(_1329_),
    .A2(_1113_));
 sg13g2_a21oi_1 _5263_ (.A1(_1327_),
    .A2(_1329_),
    .Y(_1330_),
    .B1(_1322_));
 sg13g2_nand2b_1 _5264_ (.Y(_1331_),
    .B(_3312_),
    .A_N(_1194_));
 sg13g2_nand2b_1 _5265_ (.Y(_1332_),
    .B(_1127_),
    .A_N(net1063));
 sg13g2_a21oi_1 _5266_ (.A1(_1143_),
    .A2(_1332_),
    .Y(_1333_),
    .B1(_1142_));
 sg13g2_a21oi_1 _5267_ (.A1(_1175_),
    .A2(_1178_),
    .Y(_1334_),
    .B1(\vgademo.v_count[7] ));
 sg13g2_a221oi_1 _5268_ (.B2(_1333_),
    .C1(_1334_),
    .B1(_1319_),
    .A1(_1181_),
    .Y(_1335_),
    .A2(_1182_));
 sg13g2_o21ai_1 _5269_ (.B1(_1331_),
    .Y(_1336_),
    .A1(_1320_),
    .A2(_1335_));
 sg13g2_or2_1 _5270_ (.X(_1337_),
    .B(_1336_),
    .A(_1330_));
 sg13g2_or3_1 _5271_ (.A(_1081_),
    .B(_1322_),
    .C(_1327_),
    .X(_1338_));
 sg13g2_or3_2 _5272_ (.A(_1083_),
    .B(_1322_),
    .C(_1326_),
    .X(_1339_));
 sg13g2_and2_1 _5273_ (.A(net958),
    .B(_1338_),
    .X(_1340_));
 sg13g2_o21ai_1 _5274_ (.B1(_1338_),
    .Y(_1341_),
    .A1(_1330_),
    .A2(_1336_));
 sg13g2_mux2_1 _5275_ (.A0(_0076_),
    .A1(_0051_),
    .S(net956),
    .X(_1342_));
 sg13g2_nor2_1 _5276_ (.A(\vgademo.b_cos[9] ),
    .B(_1342_),
    .Y(_1343_));
 sg13g2_nor2_1 _5277_ (.A(_0050_),
    .B(net954),
    .Y(_1344_));
 sg13g2_a21oi_1 _5278_ (.A1(_3207_),
    .A2(net953),
    .Y(_1345_),
    .B1(_1344_));
 sg13g2_nor2_1 _5279_ (.A(\vgademo.b_cos[8] ),
    .B(_1345_),
    .Y(_1346_));
 sg13g2_mux2_1 _5280_ (.A0(_0070_),
    .A1(_0048_),
    .S(net956),
    .X(_1347_));
 sg13g2_nor2_1 _5281_ (.A(\vgademo.b_cos[7] ),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_xnor2_1 _5282_ (.Y(_1349_),
    .A(_3235_),
    .B(_1347_));
 sg13g2_nor2_1 _5283_ (.A(_3234_),
    .B(\vgademo.plane_du[2] ),
    .Y(_1350_));
 sg13g2_nand2_1 _5284_ (.Y(_1351_),
    .A(\vgademo.b_cos[6] ),
    .B(_1350_));
 sg13g2_o21ai_1 _5285_ (.B1(_0049_),
    .Y(_1352_),
    .A1(\vgademo.b_cos[6] ),
    .A2(_1350_));
 sg13g2_nand2_1 _5286_ (.Y(_1353_),
    .A(_1351_),
    .B(_1352_));
 sg13g2_nor2_2 _5287_ (.A(\vgademo.bayer_j[0] ),
    .B(_3234_),
    .Y(_1354_));
 sg13g2_nor2_1 _5288_ (.A(\vgademo.b_cos[6] ),
    .B(_1354_),
    .Y(_1355_));
 sg13g2_nand2_1 _5289_ (.Y(_1356_),
    .A(net1056),
    .B(_1354_));
 sg13g2_a21oi_1 _5290_ (.A1(net1056),
    .A2(_1354_),
    .Y(_1357_),
    .B1(_0071_));
 sg13g2_o21ai_1 _5291_ (.B1(net953),
    .Y(_1358_),
    .A1(_1355_),
    .A2(_1357_));
 sg13g2_o21ai_1 _5292_ (.B1(_1358_),
    .Y(_1359_),
    .A1(net953),
    .A2(_1353_));
 sg13g2_a21oi_2 _5293_ (.B1(_1348_),
    .Y(_1360_),
    .A2(_1359_),
    .A1(_1349_));
 sg13g2_inv_1 _5294_ (.Y(_1361_),
    .A(_1360_));
 sg13g2_xnor2_1 _5295_ (.Y(_1362_),
    .A(_3237_),
    .B(_1345_));
 sg13g2_a21oi_2 _5296_ (.B1(_1346_),
    .Y(_1363_),
    .A2(_1362_),
    .A1(_1361_));
 sg13g2_inv_1 _5297_ (.Y(_1364_),
    .A(_1363_));
 sg13g2_xnor2_1 _5298_ (.Y(_1365_),
    .A(_3238_),
    .B(_1342_));
 sg13g2_a21oi_1 _5299_ (.A1(_1364_),
    .A2(_1365_),
    .Y(_1366_),
    .B1(_1343_));
 sg13g2_mux2_1 _5300_ (.A0(_0062_),
    .A1(_0052_),
    .S(net956),
    .X(_1367_));
 sg13g2_xnor2_1 _5301_ (.Y(_1368_),
    .A(net1054),
    .B(_1367_));
 sg13g2_nand2b_1 _5302_ (.Y(_1369_),
    .B(_1368_),
    .A_N(_1366_));
 sg13g2_xnor2_1 _5303_ (.Y(_1370_),
    .A(_1366_),
    .B(_1368_));
 sg13g2_xnor2_1 _5304_ (.Y(_1371_),
    .A(_1360_),
    .B(_1362_));
 sg13g2_xor2_1 _5305_ (.B(_1362_),
    .A(_1360_),
    .X(_1372_));
 sg13g2_o21ai_1 _5306_ (.B1(net1083),
    .Y(_1373_),
    .A1(net1090),
    .A2(net1085));
 sg13g2_nand2_1 _5307_ (.Y(_1374_),
    .A(net1074),
    .B(_3199_));
 sg13g2_nor2_1 _5308_ (.A(net1079),
    .B(_1374_),
    .Y(_1375_));
 sg13g2_a21oi_1 _5309_ (.A1(_1373_),
    .A2(_1375_),
    .Y(_1376_),
    .B1(_0079_));
 sg13g2_nand3_1 _5310_ (.B(_3199_),
    .C(_1204_),
    .A(net1074),
    .Y(_1377_));
 sg13g2_nand2_1 _5311_ (.Y(_1378_),
    .A(_3200_),
    .B(net1083));
 sg13g2_nor3_1 _5312_ (.A(_1046_),
    .B(_1377_),
    .C(_1378_),
    .Y(_1379_));
 sg13g2_o21ai_1 _5313_ (.B1(net1070),
    .Y(_1380_),
    .A1(_1376_),
    .A2(_1379_));
 sg13g2_and3_2 _5314_ (.X(_1381_),
    .A(_3197_),
    .B(_1050_),
    .C(_1380_));
 sg13g2_a21oi_2 _5315_ (.B1(net1069),
    .Y(_1382_),
    .A2(_1044_),
    .A1(net1070));
 sg13g2_nand2_1 _5316_ (.Y(_1383_),
    .A(\vgademo.a_scrolly[13] ),
    .B(net1067));
 sg13g2_nor2_1 _5317_ (.A(_1382_),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_nor2_1 _5318_ (.A(_1065_),
    .B(_1384_),
    .Y(_1385_));
 sg13g2_o21ai_1 _5319_ (.B1(_1064_),
    .Y(_1386_),
    .A1(_1382_),
    .A2(_1383_));
 sg13g2_a21o_2 _5320_ (.A2(_1386_),
    .A1(_1063_),
    .B1(_1381_),
    .X(_1387_));
 sg13g2_nor2_1 _5321_ (.A(_1055_),
    .B(_1374_),
    .Y(_1388_));
 sg13g2_a21oi_1 _5322_ (.A1(_1107_),
    .A2(_1388_),
    .Y(_1389_),
    .B1(_1060_));
 sg13g2_nor4_1 _5323_ (.A(_1039_),
    .B(_1055_),
    .C(_1201_),
    .D(_1374_),
    .Y(_1390_));
 sg13g2_nor4_2 _5324_ (.A(net1067),
    .B(_1049_),
    .C(_1389_),
    .Y(_1391_),
    .D(_1390_));
 sg13g2_xor2_1 _5325_ (.B(_1218_),
    .A(_0077_),
    .X(_1392_));
 sg13g2_nand3_1 _5326_ (.B(_1039_),
    .C(_1373_),
    .A(_0074_),
    .Y(_1393_));
 sg13g2_nand2_1 _5327_ (.Y(_1394_),
    .A(_1041_),
    .B(_1393_));
 sg13g2_nor2_1 _5328_ (.A(net1045),
    .B(_1393_),
    .Y(_1395_));
 sg13g2_xnor2_1 _5329_ (.Y(_1396_),
    .A(net1045),
    .B(_1394_));
 sg13g2_a221oi_1 _5330_ (.B2(_1386_),
    .C1(_1387_),
    .B1(_1396_),
    .A1(net993),
    .Y(_1397_),
    .A2(_1392_));
 sg13g2_nor2_1 _5331_ (.A(_0030_),
    .B(net954),
    .Y(_1398_));
 sg13g2_nor3_1 _5332_ (.A(net1096),
    .B(net1093),
    .C(net1095),
    .Y(_1399_));
 sg13g2_and2_1 _5333_ (.A(_3193_),
    .B(_1399_),
    .X(_1400_));
 sg13g2_nor2_1 _5334_ (.A(_3192_),
    .B(_1400_),
    .Y(_1401_));
 sg13g2_nand2_1 _5335_ (.Y(_1402_),
    .A(\vgademo.h_count[6] ),
    .B(_1401_));
 sg13g2_inv_1 _5336_ (.Y(_1403_),
    .A(_1402_));
 sg13g2_nand2_1 _5337_ (.Y(_1404_),
    .A(_0036_),
    .B(_1402_));
 sg13g2_xor2_1 _5338_ (.B(_1404_),
    .A(_0037_),
    .X(_1405_));
 sg13g2_a21oi_2 _5339_ (.B1(_1398_),
    .Y(_1406_),
    .A2(_1405_),
    .A1(net953));
 sg13g2_nand2b_1 _5340_ (.Y(_1407_),
    .B(_1397_),
    .A_N(_1406_));
 sg13g2_nand2b_1 _5341_ (.Y(_1408_),
    .B(_1406_),
    .A_N(_1397_));
 sg13g2_xnor2_1 _5342_ (.Y(_1409_),
    .A(_1397_),
    .B(_1406_));
 sg13g2_inv_1 _5343_ (.Y(_1410_),
    .A(_1409_));
 sg13g2_o21ai_1 _5344_ (.B1(net993),
    .Y(_1411_),
    .A1(_1037_),
    .A2(_1219_));
 sg13g2_xnor2_1 _5345_ (.Y(_1412_),
    .A(_0074_),
    .B(_1373_));
 sg13g2_o21ai_1 _5346_ (.B1(_1411_),
    .Y(_1413_),
    .A1(_1385_),
    .A2(_1412_));
 sg13g2_nor2_1 _5347_ (.A(_1387_),
    .B(_1413_),
    .Y(_1414_));
 sg13g2_xnor2_1 _5348_ (.Y(_1415_),
    .A(_3194_),
    .B(_1402_));
 sg13g2_nor2_1 _5349_ (.A(_0045_),
    .B(net953),
    .Y(_1416_));
 sg13g2_a21oi_2 _5350_ (.B1(_1416_),
    .Y(_1417_),
    .A2(_1415_),
    .A1(net952));
 sg13g2_inv_1 _5351_ (.Y(_1418_),
    .A(_1417_));
 sg13g2_nor2b_2 _5352_ (.A(_1414_),
    .B_N(_1417_),
    .Y(_1419_));
 sg13g2_inv_1 _5353_ (.Y(_1420_),
    .A(_1419_));
 sg13g2_nor3_1 _5354_ (.A(_1387_),
    .B(_1413_),
    .C(_1417_),
    .Y(_1421_));
 sg13g2_o21ai_1 _5355_ (.B1(_1373_),
    .Y(_1422_),
    .A1(net1090),
    .A2(_1039_));
 sg13g2_a221oi_1 _5356_ (.B2(_1386_),
    .C1(_1387_),
    .B1(_1422_),
    .A1(net1083),
    .Y(_1423_),
    .A2(net993));
 sg13g2_nor2_1 _5357_ (.A(_0029_),
    .B(net953),
    .Y(_1424_));
 sg13g2_xnor2_1 _5358_ (.Y(_1425_),
    .A(_0035_),
    .B(_1401_));
 sg13g2_a21oi_2 _5359_ (.B1(_1424_),
    .Y(_1426_),
    .A2(_1425_),
    .A1(net952));
 sg13g2_nor2b_1 _5360_ (.A(_1426_),
    .B_N(_1423_),
    .Y(_1427_));
 sg13g2_nor2_2 _5361_ (.A(_1063_),
    .B(_1385_),
    .Y(_1428_));
 sg13g2_a22oi_1 _5362_ (.Y(_1429_),
    .B1(_1428_),
    .B2(_1211_),
    .A2(net993),
    .A1(_3204_));
 sg13g2_nor2_1 _5363_ (.A(_1381_),
    .B(_1429_),
    .Y(_1430_));
 sg13g2_inv_1 _5364_ (.Y(_1431_),
    .A(_1430_));
 sg13g2_xnor2_1 _5365_ (.Y(_1432_),
    .A(_3192_),
    .B(_1400_));
 sg13g2_mux2_1 _5366_ (.A0(_1432_),
    .A1(_0046_),
    .S(net955),
    .X(_1433_));
 sg13g2_or2_1 _5367_ (.X(_1434_),
    .B(_1433_),
    .A(_1431_));
 sg13g2_a22oi_1 _5368_ (.Y(_1435_),
    .B1(_1391_),
    .B2(_0063_),
    .A2(_1386_),
    .A1(net1090));
 sg13g2_nand2b_1 _5369_ (.Y(_1436_),
    .B(_1435_),
    .A_N(_1387_));
 sg13g2_xor2_1 _5370_ (.B(_1399_),
    .A(_0043_),
    .X(_1437_));
 sg13g2_mux2_2 _5371_ (.A0(_1437_),
    .A1(_0028_),
    .S(net956),
    .X(_1438_));
 sg13g2_nor2_1 _5372_ (.A(_1436_),
    .B(_1438_),
    .Y(_1439_));
 sg13g2_xor2_1 _5373_ (.B(\vgademo.h_count[2] ),
    .A(net1097),
    .X(_1440_));
 sg13g2_mux2_1 _5374_ (.A0(_1440_),
    .A1(_0027_),
    .S(net956),
    .X(_1441_));
 sg13g2_xor2_1 _5375_ (.B(_3324_),
    .A(_0033_),
    .X(_1442_));
 sg13g2_mux2_2 _5376_ (.A0(_1442_),
    .A1(_0047_),
    .S(_1341_),
    .X(_1443_));
 sg13g2_a21oi_2 _5377_ (.B1(_1387_),
    .Y(_1444_),
    .A2(_1443_),
    .A1(_1441_));
 sg13g2_nand2_1 _5378_ (.Y(_1445_),
    .A(_1436_),
    .B(_1438_));
 sg13g2_xnor2_1 _5379_ (.Y(_1446_),
    .A(_1436_),
    .B(_1438_));
 sg13g2_a21oi_2 _5380_ (.B1(_1439_),
    .Y(_1447_),
    .A2(_1445_),
    .A1(_1444_));
 sg13g2_xnor2_1 _5381_ (.Y(_1448_),
    .A(_1431_),
    .B(_1433_));
 sg13g2_o21ai_1 _5382_ (.B1(_1434_),
    .Y(_1449_),
    .A1(_1447_),
    .A2(_1448_));
 sg13g2_xnor2_1 _5383_ (.Y(_1450_),
    .A(_1423_),
    .B(_1426_));
 sg13g2_a21o_1 _5384_ (.A2(_1450_),
    .A1(_1449_),
    .B1(_1427_),
    .X(_1451_));
 sg13g2_a221oi_1 _5385_ (.B2(_1450_),
    .C1(_1427_),
    .B1(_1449_),
    .A1(_1414_),
    .Y(_1452_),
    .A2(_1418_));
 sg13g2_nor3_2 _5386_ (.A(_1410_),
    .B(_1419_),
    .C(_1452_),
    .Y(_1453_));
 sg13g2_nand3b_1 _5387_ (.B(_1409_),
    .C(_1420_),
    .Y(_1454_),
    .A_N(_1452_));
 sg13g2_nand2_2 _5388_ (.Y(_1455_),
    .A(_1407_),
    .B(_1454_));
 sg13g2_xnor2_1 _5389_ (.Y(_1456_),
    .A(_0079_),
    .B(_1042_));
 sg13g2_or2_1 _5390_ (.X(_1457_),
    .B(_1456_),
    .A(_1395_));
 sg13g2_inv_1 _5391_ (.Y(_1458_),
    .A(_1457_));
 sg13g2_xor2_1 _5392_ (.B(_1456_),
    .A(_1395_),
    .X(_1459_));
 sg13g2_o21ai_1 _5393_ (.B1(net1074),
    .Y(_1460_),
    .A1(net1077),
    .A2(_1038_));
 sg13g2_inv_1 _5394_ (.Y(_1461_),
    .A(_1460_));
 sg13g2_and3_1 _5395_ (.X(_1462_),
    .A(_0077_),
    .B(_1038_),
    .C(_1218_));
 sg13g2_a21oi_1 _5396_ (.A1(_1037_),
    .A2(net1041),
    .Y(_1463_),
    .B1(_1462_));
 sg13g2_a22oi_1 _5397_ (.Y(_1464_),
    .B1(_1463_),
    .B2(_1460_),
    .A2(_1462_),
    .A1(net1074));
 sg13g2_a22oi_1 _5398_ (.Y(_1465_),
    .B1(_1464_),
    .B2(net993),
    .A2(_1459_),
    .A1(_1428_));
 sg13g2_nor2_2 _5399_ (.A(_1381_),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_nor2_1 _5400_ (.A(_0044_),
    .B(net953),
    .Y(_1467_));
 sg13g2_nor3_2 _5401_ (.A(\vgademo.h_count[7] ),
    .B(\vgademo.h_count[8] ),
    .C(_1403_),
    .Y(_1468_));
 sg13g2_xnor2_1 _5402_ (.Y(_1469_),
    .A(\vgademo.h_count[9] ),
    .B(_1468_));
 sg13g2_a21oi_2 _5403_ (.B1(_1467_),
    .Y(_1470_),
    .A2(_1469_),
    .A1(net953));
 sg13g2_nor2b_1 _5404_ (.A(_1470_),
    .B_N(_1466_),
    .Y(_1471_));
 sg13g2_xnor2_1 _5405_ (.Y(_1472_),
    .A(_1466_),
    .B(_1470_));
 sg13g2_xor2_1 _5406_ (.B(_1472_),
    .A(_1455_),
    .X(_1473_));
 sg13g2_xnor2_1 _5407_ (.Y(_1474_),
    .A(_1455_),
    .B(_1472_));
 sg13g2_xor2_1 _5408_ (.B(_1450_),
    .A(_1449_),
    .X(_1475_));
 sg13g2_xnor2_1 _5409_ (.Y(_1476_),
    .A(_1449_),
    .B(_1450_));
 sg13g2_xor2_1 _5410_ (.B(_1448_),
    .A(_1447_),
    .X(_1477_));
 sg13g2_xnor2_1 _5411_ (.Y(_1478_),
    .A(_1447_),
    .B(_1448_));
 sg13g2_xnor2_1 _5412_ (.Y(_1479_),
    .A(_1444_),
    .B(_1446_));
 sg13g2_xor2_1 _5413_ (.B(_1446_),
    .A(_1444_),
    .X(_1480_));
 sg13g2_nor2b_1 _5414_ (.A(_1387_),
    .B_N(_1441_),
    .Y(_1481_));
 sg13g2_xnor2_1 _5415_ (.Y(_1482_),
    .A(_1443_),
    .B(_1481_));
 sg13g2_nor2_1 _5416_ (.A(_1479_),
    .B(_1482_),
    .Y(_1483_));
 sg13g2_or2_1 _5417_ (.X(_1484_),
    .B(_1482_),
    .A(net941));
 sg13g2_nand2_2 _5418_ (.Y(_1485_),
    .A(net940),
    .B(_1484_));
 sg13g2_nor2_1 _5419_ (.A(net932),
    .B(net938),
    .Y(_1486_));
 sg13g2_nand2b_2 _5420_ (.Y(_1487_),
    .B(net930),
    .A_N(_1485_));
 sg13g2_a221oi_1 _5421_ (.B2(_1451_),
    .C1(_1421_),
    .B1(_1420_),
    .A1(_1407_),
    .Y(_1488_),
    .A2(_1408_));
 sg13g2_o21ai_1 _5422_ (.B1(_1410_),
    .Y(_1489_),
    .A1(_1419_),
    .A2(_1452_));
 sg13g2_or3_1 _5423_ (.A(_1409_),
    .B(_1419_),
    .C(_1452_),
    .X(_1490_));
 sg13g2_o21ai_1 _5424_ (.B1(_1409_),
    .Y(_1491_),
    .A1(_1419_),
    .A2(_1452_));
 sg13g2_nor2_1 _5425_ (.A(_1453_),
    .B(_1488_),
    .Y(_1492_));
 sg13g2_nand2_1 _5426_ (.Y(_1493_),
    .A(_1454_),
    .B(_1489_));
 sg13g2_nor2_1 _5427_ (.A(net928),
    .B(net941),
    .Y(_1494_));
 sg13g2_nor2_2 _5428_ (.A(net939),
    .B(net941),
    .Y(_1495_));
 sg13g2_nand2_2 _5429_ (.Y(_1496_),
    .A(net938),
    .B(_1480_));
 sg13g2_nand2_1 _5430_ (.Y(_1497_),
    .A(net934),
    .B(_1495_));
 sg13g2_and3_1 _5431_ (.X(_1498_),
    .A(_1487_),
    .B(net908),
    .C(_1497_));
 sg13g2_nand3_1 _5432_ (.B(net907),
    .C(_1497_),
    .A(_1487_),
    .Y(_1499_));
 sg13g2_or2_1 _5433_ (.X(_1500_),
    .B(_1421_),
    .A(_1419_));
 sg13g2_xnor2_1 _5434_ (.Y(_1501_),
    .A(_1451_),
    .B(_1500_));
 sg13g2_xor2_1 _5435_ (.B(_1500_),
    .A(_1451_),
    .X(_1502_));
 sg13g2_nor2_2 _5436_ (.A(net928),
    .B(_1495_),
    .Y(_1503_));
 sg13g2_nand2_2 _5437_ (.Y(_1504_),
    .A(_1479_),
    .B(_1482_));
 sg13g2_nand2_2 _5438_ (.Y(_1505_),
    .A(net939),
    .B(net941));
 sg13g2_or2_2 _5439_ (.X(_1506_),
    .B(_1504_),
    .A(net938));
 sg13g2_a21oi_2 _5440_ (.B1(net924),
    .Y(_1507_),
    .A2(_1506_),
    .A1(_1503_));
 sg13g2_and2_1 _5441_ (.A(net930),
    .B(_1485_),
    .X(_1508_));
 sg13g2_o21ai_1 _5442_ (.B1(net910),
    .Y(_1509_),
    .A1(_1507_),
    .A2(_1508_));
 sg13g2_a21oi_1 _5443_ (.A1(_1499_),
    .A2(_1509_),
    .Y(_1510_),
    .B1(net906));
 sg13g2_xnor2_1 _5444_ (.Y(_1511_),
    .A(_1349_),
    .B(_1359_));
 sg13g2_inv_2 _5445_ (.Y(_1512_),
    .A(net937));
 sg13g2_nor3_2 _5446_ (.A(_1453_),
    .B(_1488_),
    .C(net937),
    .Y(_1513_));
 sg13g2_nand3_1 _5447_ (.B(_1489_),
    .C(_1512_),
    .A(_1454_),
    .Y(_1514_));
 sg13g2_nand2_1 _5448_ (.Y(_1515_),
    .A(net939),
    .B(_1480_));
 sg13g2_nand2_1 _5449_ (.Y(_1516_),
    .A(net932),
    .B(_1515_));
 sg13g2_nor2_1 _5450_ (.A(_1475_),
    .B(net940),
    .Y(_1517_));
 sg13g2_nand3_1 _5451_ (.B(net938),
    .C(_1504_),
    .A(net928),
    .Y(_1518_));
 sg13g2_nand3_1 _5452_ (.B(_1516_),
    .C(_1518_),
    .A(_1487_),
    .Y(_1519_));
 sg13g2_nor3_2 _5453_ (.A(_1453_),
    .B(_1488_),
    .C(_1512_),
    .Y(_1520_));
 sg13g2_nand3_1 _5454_ (.B(_1489_),
    .C(net937),
    .A(_1454_),
    .Y(_1521_));
 sg13g2_nand2_2 _5455_ (.Y(_1522_),
    .A(_1478_),
    .B(net941));
 sg13g2_o21ai_1 _5456_ (.B1(_1504_),
    .Y(_1523_),
    .A1(net940),
    .A2(_1480_));
 sg13g2_nor2_2 _5457_ (.A(net928),
    .B(_1478_),
    .Y(_1524_));
 sg13g2_nor2_1 _5458_ (.A(net928),
    .B(_1523_),
    .Y(_1525_));
 sg13g2_nor2_1 _5459_ (.A(net932),
    .B(_1495_),
    .Y(_1526_));
 sg13g2_nand2_1 _5460_ (.Y(_1527_),
    .A(net929),
    .B(_1496_));
 sg13g2_or2_1 _5461_ (.X(_1528_),
    .B(_1482_),
    .A(net940));
 sg13g2_a21oi_1 _5462_ (.A1(_1526_),
    .A2(_1528_),
    .Y(_1529_),
    .B1(_1525_));
 sg13g2_a22oi_1 _5463_ (.Y(_1530_),
    .B1(_1520_),
    .B2(_1529_),
    .A2(_1519_),
    .A1(_1513_));
 sg13g2_a21oi_2 _5464_ (.B1(net937),
    .Y(_1531_),
    .A2(_1489_),
    .A1(_1454_));
 sg13g2_nor2_1 _5465_ (.A(net930),
    .B(_1506_),
    .Y(_1532_));
 sg13g2_or2_1 _5466_ (.X(_1533_),
    .B(_1506_),
    .A(net930));
 sg13g2_nor2_1 _5467_ (.A(net924),
    .B(_1533_),
    .Y(_1534_));
 sg13g2_a21o_2 _5468_ (.A2(_1482_),
    .A1(_1480_),
    .B1(net940),
    .X(_1535_));
 sg13g2_and3_1 _5469_ (.X(_1536_),
    .A(net930),
    .B(_1485_),
    .C(_1535_));
 sg13g2_o21ai_1 _5470_ (.B1(net941),
    .Y(_1537_),
    .A1(net933),
    .A2(net938));
 sg13g2_nand2_1 _5471_ (.Y(_1538_),
    .A(net924),
    .B(_1537_));
 sg13g2_mux2_1 _5472_ (.A0(_1536_),
    .A1(_1537_),
    .S(net925),
    .X(_1539_));
 sg13g2_and2_1 _5473_ (.A(net908),
    .B(_1539_),
    .X(_1540_));
 sg13g2_nor2_2 _5474_ (.A(net933),
    .B(_1496_),
    .Y(_1541_));
 sg13g2_nand2_1 _5475_ (.Y(_1542_),
    .A(net931),
    .B(_1495_));
 sg13g2_xnor2_1 _5476_ (.Y(_1543_),
    .A(_1480_),
    .B(_1482_));
 sg13g2_xnor2_1 _5477_ (.Y(_1544_),
    .A(net941),
    .B(_1482_));
 sg13g2_a21oi_1 _5478_ (.A1(net932),
    .A2(_1496_),
    .Y(_1545_),
    .B1(_1543_));
 sg13g2_a21oi_1 _5479_ (.A1(_1542_),
    .A2(_1545_),
    .Y(_1546_),
    .B1(net922));
 sg13g2_a221oi_1 _5480_ (.B2(_1545_),
    .C1(net922),
    .B1(_1542_),
    .A1(_1490_),
    .Y(_1547_),
    .A2(_1491_));
 sg13g2_a221oi_1 _5481_ (.B2(net907),
    .C1(_1547_),
    .B1(_1539_),
    .A1(_1531_),
    .Y(_1548_),
    .A2(_1534_));
 sg13g2_o21ai_1 _5482_ (.B1(_1548_),
    .Y(_1549_),
    .A1(net919),
    .A2(_1530_));
 sg13g2_a21o_1 _5483_ (.A2(_1549_),
    .A1(net906),
    .B1(_1510_),
    .X(_1550_));
 sg13g2_xnor2_1 _5484_ (.Y(_1551_),
    .A(_1363_),
    .B(_1365_));
 sg13g2_xor2_1 _5485_ (.B(_1365_),
    .A(_1363_),
    .X(_1552_));
 sg13g2_nand2_2 _5486_ (.Y(_1553_),
    .A(net939),
    .B(_1504_));
 sg13g2_nand2_2 _5487_ (.Y(_1554_),
    .A(net939),
    .B(_1543_));
 sg13g2_nand3_1 _5488_ (.B(_1496_),
    .C(_1554_),
    .A(net934),
    .Y(_1555_));
 sg13g2_nand2_1 _5489_ (.Y(_1556_),
    .A(_1518_),
    .B(_1555_));
 sg13g2_nand2_1 _5490_ (.Y(_1557_),
    .A(net933),
    .B(_1553_));
 sg13g2_nand3_1 _5491_ (.B(_1518_),
    .C(_1557_),
    .A(_1487_),
    .Y(_1558_));
 sg13g2_a22oi_1 _5492_ (.Y(_1559_),
    .B1(_1558_),
    .B2(_1520_),
    .A2(_1556_),
    .A1(_1513_));
 sg13g2_nand2b_1 _5493_ (.Y(_1560_),
    .B(net926),
    .A_N(_1559_));
 sg13g2_nor2_2 _5494_ (.A(net938),
    .B(_1484_),
    .Y(_1561_));
 sg13g2_nand2_1 _5495_ (.Y(_1562_),
    .A(net939),
    .B(_1544_));
 sg13g2_nand3_1 _5496_ (.B(_1496_),
    .C(_1562_),
    .A(net929),
    .Y(_1563_));
 sg13g2_nand2_1 _5497_ (.Y(_1564_),
    .A(net919),
    .B(_1563_));
 sg13g2_a21oi_1 _5498_ (.A1(_1538_),
    .A2(_1564_),
    .Y(_1565_),
    .B1(net911));
 sg13g2_nor3_1 _5499_ (.A(_1474_),
    .B(_1547_),
    .C(_1565_),
    .Y(_1566_));
 sg13g2_nand2b_2 _5500_ (.Y(_1567_),
    .B(net931),
    .A_N(_1554_));
 sg13g2_and3_1 _5501_ (.X(_1568_),
    .A(net908),
    .B(_1497_),
    .C(_1567_));
 sg13g2_a21o_1 _5502_ (.A2(_1567_),
    .A1(net926),
    .B1(_1507_),
    .X(_1569_));
 sg13g2_and2_1 _5503_ (.A(net920),
    .B(_1561_),
    .X(_1570_));
 sg13g2_nand3_1 _5504_ (.B(_1496_),
    .C(_1562_),
    .A(net932),
    .Y(_1571_));
 sg13g2_and2_1 _5505_ (.A(net917),
    .B(_1571_),
    .X(_1572_));
 sg13g2_mux2_1 _5506_ (.A0(_1567_),
    .A1(_1571_),
    .S(net919),
    .X(_1573_));
 sg13g2_a21oi_1 _5507_ (.A1(net910),
    .A2(_1573_),
    .Y(_1574_),
    .B1(_1568_));
 sg13g2_a221oi_1 _5508_ (.B2(_1569_),
    .C1(net906),
    .B1(_1520_),
    .A1(_1498_),
    .Y(_1575_),
    .A2(_1511_));
 sg13g2_o21ai_1 _5509_ (.B1(_1575_),
    .Y(_1576_),
    .A1(_1511_),
    .A2(_1574_));
 sg13g2_a21oi_1 _5510_ (.A1(_1560_),
    .A2(_1566_),
    .Y(_1577_),
    .B1(net935));
 sg13g2_a221oi_1 _5511_ (.B2(_1577_),
    .C1(_1552_),
    .B1(_1576_),
    .A1(net935),
    .Y(_1578_),
    .A2(_1550_));
 sg13g2_nand3_1 _5512_ (.B(_1503_),
    .C(_1506_),
    .A(net924),
    .Y(_1579_));
 sg13g2_o21ai_1 _5513_ (.B1(_1508_),
    .Y(_1580_),
    .A1(net940),
    .A2(net919));
 sg13g2_a21oi_1 _5514_ (.A1(_1579_),
    .A2(_1580_),
    .Y(_1581_),
    .B1(net907));
 sg13g2_nor2_1 _5515_ (.A(net910),
    .B(_1533_),
    .Y(_1582_));
 sg13g2_o21ai_1 _5516_ (.B1(_1474_),
    .Y(_1583_),
    .A1(_1581_),
    .A2(_1582_));
 sg13g2_nand2_1 _5517_ (.Y(_1584_),
    .A(net938),
    .B(_1483_));
 sg13g2_nand2_1 _5518_ (.Y(_1585_),
    .A(net934),
    .B(_1584_));
 sg13g2_a21o_1 _5519_ (.A2(_1585_),
    .A1(_1554_),
    .B1(net925),
    .X(_1586_));
 sg13g2_nor2_1 _5520_ (.A(net907),
    .B(_1586_),
    .Y(_1587_));
 sg13g2_nand3_1 _5521_ (.B(_1503_),
    .C(_1544_),
    .A(net922),
    .Y(_1588_));
 sg13g2_a21oi_1 _5522_ (.A1(_1586_),
    .A2(_1588_),
    .Y(_1589_),
    .B1(net907));
 sg13g2_o21ai_1 _5523_ (.B1(net906),
    .Y(_1590_),
    .A1(_1540_),
    .A2(_1589_));
 sg13g2_a21oi_1 _5524_ (.A1(_1583_),
    .A2(_1590_),
    .Y(_1591_),
    .B1(_1371_));
 sg13g2_nor2_2 _5525_ (.A(net935),
    .B(net937),
    .Y(_1592_));
 sg13g2_nand2_1 _5526_ (.Y(_1593_),
    .A(_1371_),
    .B(_1512_));
 sg13g2_or2_1 _5527_ (.X(_1594_),
    .B(_1518_),
    .A(net919));
 sg13g2_a21oi_1 _5528_ (.A1(_1588_),
    .A2(_1594_),
    .Y(_1595_),
    .B1(net907));
 sg13g2_nor3_1 _5529_ (.A(_1540_),
    .B(_1547_),
    .C(_1595_),
    .Y(_1596_));
 sg13g2_nor2_1 _5530_ (.A(_1474_),
    .B(_1596_),
    .Y(_1597_));
 sg13g2_o21ai_1 _5531_ (.B1(_1592_),
    .Y(_1598_),
    .A1(_1510_),
    .A2(_1597_));
 sg13g2_nand2_2 _5532_ (.Y(_1599_),
    .A(_1371_),
    .B(_1511_));
 sg13g2_o21ai_1 _5533_ (.B1(net906),
    .Y(_1600_),
    .A1(_1587_),
    .A2(_1595_));
 sg13g2_nor3_2 _5534_ (.A(_1453_),
    .B(_1488_),
    .C(net919),
    .Y(_1601_));
 sg13g2_nand2_1 _5535_ (.Y(_1602_),
    .A(_1532_),
    .B(_1601_));
 sg13g2_o21ai_1 _5536_ (.B1(net920),
    .Y(_1603_),
    .A1(net934),
    .A2(_1535_));
 sg13g2_nor2_1 _5537_ (.A(net931),
    .B(_1505_),
    .Y(_1604_));
 sg13g2_o21ai_1 _5538_ (.B1(_1538_),
    .Y(_1605_),
    .A1(_1603_),
    .A2(_1604_));
 sg13g2_a22oi_1 _5539_ (.Y(_1606_),
    .B1(_1605_),
    .B2(net907),
    .A2(_1602_),
    .A1(_1474_));
 sg13g2_a21oi_1 _5540_ (.A1(_1600_),
    .A2(_1606_),
    .Y(_1607_),
    .B1(_1599_));
 sg13g2_nor3_1 _5541_ (.A(_1551_),
    .B(_1591_),
    .C(_1607_),
    .Y(_1608_));
 sg13g2_a21o_1 _5542_ (.A2(_1608_),
    .A1(_1598_),
    .B1(_1578_),
    .X(_1609_));
 sg13g2_o21ai_1 _5543_ (.B1(_1369_),
    .Y(_1610_),
    .A1(_3239_),
    .A2(_1367_));
 sg13g2_nand2b_2 _5544_ (.Y(_1611_),
    .B(\vgademo.b_cos[10] ),
    .A_N(\vgademo.b_cos[11] ));
 sg13g2_xnor2_1 _5545_ (.Y(_1612_),
    .A(\vgademo.b_cos[10] ),
    .B(\vgademo.b_cos[11] ));
 sg13g2_xor2_1 _5546_ (.B(\vgademo.b_cos[11] ),
    .A(\vgademo.b_cos[10] ),
    .X(_1613_));
 sg13g2_nand2_1 _5547_ (.Y(_1614_),
    .A(\vgademo.plane_du[8] ),
    .B(net956));
 sg13g2_o21ai_1 _5548_ (.B1(_1614_),
    .Y(_1615_),
    .A1(_3186_),
    .A2(net956));
 sg13g2_xnor2_1 _5549_ (.Y(_1616_),
    .A(_1612_),
    .B(_1615_));
 sg13g2_xor2_1 _5550_ (.B(_1616_),
    .A(_1610_),
    .X(_1617_));
 sg13g2_nor2_2 _5551_ (.A(_1371_),
    .B(_1512_),
    .Y(_1618_));
 sg13g2_nand2_1 _5552_ (.Y(_1619_),
    .A(net935),
    .B(net937));
 sg13g2_or4_1 _5553_ (.A(net912),
    .B(net920),
    .C(_1524_),
    .D(_1541_),
    .X(_1620_));
 sg13g2_nand2_1 _5554_ (.Y(_1621_),
    .A(net930),
    .B(_1506_));
 sg13g2_nor2_1 _5555_ (.A(net930),
    .B(_1485_),
    .Y(_1622_));
 sg13g2_nand2b_1 _5556_ (.Y(_1623_),
    .B(net924),
    .A_N(_1622_));
 sg13g2_nand3_1 _5557_ (.B(_1621_),
    .C(_1623_),
    .A(net911),
    .Y(_1624_));
 sg13g2_a21oi_1 _5558_ (.A1(_1620_),
    .A2(_1624_),
    .Y(_1625_),
    .B1(_1619_));
 sg13g2_a21oi_1 _5559_ (.A1(net924),
    .A2(_1505_),
    .Y(_1626_),
    .B1(net930));
 sg13g2_nand3_1 _5560_ (.B(_1619_),
    .C(_1626_),
    .A(net911),
    .Y(_1627_));
 sg13g2_and3_1 _5561_ (.X(_1628_),
    .A(net933),
    .B(_1496_),
    .C(_1528_));
 sg13g2_nand2b_1 _5562_ (.Y(_1629_),
    .B(net923),
    .A_N(_1628_));
 sg13g2_nand2b_1 _5563_ (.Y(_1630_),
    .B(net935),
    .A_N(_1504_));
 sg13g2_a21oi_1 _5564_ (.A1(_1517_),
    .A2(_1630_),
    .Y(_1631_),
    .B1(_1629_));
 sg13g2_a22oi_1 _5565_ (.Y(_1632_),
    .B1(net916),
    .B2(_1631_),
    .A2(_1570_),
    .A1(net931));
 sg13g2_o21ai_1 _5566_ (.B1(_1627_),
    .Y(_1633_),
    .A1(net911),
    .A2(_1632_));
 sg13g2_o21ai_1 _5567_ (.B1(net906),
    .Y(_1634_),
    .A1(_1625_),
    .A2(_1633_));
 sg13g2_a21o_1 _5568_ (.A2(_1634_),
    .A1(_1583_),
    .B1(_1551_),
    .X(_1635_));
 sg13g2_nand3_1 _5569_ (.B(_1522_),
    .C(_1533_),
    .A(net924),
    .Y(_1636_));
 sg13g2_o21ai_1 _5570_ (.B1(net919),
    .Y(_1637_),
    .A1(_1532_),
    .A2(_1536_));
 sg13g2_nand3_1 _5571_ (.B(_1636_),
    .C(_1637_),
    .A(_1531_),
    .Y(_1638_));
 sg13g2_nor2_1 _5572_ (.A(net917),
    .B(_1555_),
    .Y(_1639_));
 sg13g2_a21oi_1 _5573_ (.A1(_1553_),
    .A2(_1585_),
    .Y(_1640_),
    .B1(net923));
 sg13g2_or3_1 _5574_ (.A(_1514_),
    .B(_1639_),
    .C(_1640_),
    .X(_1641_));
 sg13g2_a21oi_1 _5575_ (.A1(_1638_),
    .A2(_1641_),
    .Y(_1642_),
    .B1(net936));
 sg13g2_o21ai_1 _5576_ (.B1(_1506_),
    .Y(_1643_),
    .A1(_1541_),
    .A2(_1628_));
 sg13g2_mux2_1 _5577_ (.A0(_1487_),
    .A1(_1643_),
    .S(net923),
    .X(_1644_));
 sg13g2_nor3_1 _5578_ (.A(net909),
    .B(net916),
    .C(_1644_),
    .Y(_1645_));
 sg13g2_nand2_1 _5579_ (.Y(_1646_),
    .A(net919),
    .B(_1567_));
 sg13g2_and2_1 _5580_ (.A(_1535_),
    .B(_1554_),
    .X(_1647_));
 sg13g2_nand2_1 _5581_ (.Y(_1648_),
    .A(_1535_),
    .B(_1554_));
 sg13g2_o21ai_1 _5582_ (.B1(net917),
    .Y(_1649_),
    .A1(net933),
    .A2(_1647_));
 sg13g2_a21oi_1 _5583_ (.A1(_1503_),
    .A2(_1505_),
    .Y(_1650_),
    .B1(net918));
 sg13g2_nand2_1 _5584_ (.Y(_1651_),
    .A(_1484_),
    .B(_1517_));
 sg13g2_nand3_1 _5585_ (.B(_1618_),
    .C(_1649_),
    .A(net909),
    .Y(_1652_));
 sg13g2_a21oi_1 _5586_ (.A1(_1650_),
    .A2(_1651_),
    .Y(_1653_),
    .B1(_1652_));
 sg13g2_nand2_1 _5587_ (.Y(_1654_),
    .A(_1475_),
    .B(_1561_));
 sg13g2_nand3_1 _5588_ (.B(_1522_),
    .C(_1654_),
    .A(net923),
    .Y(_1655_));
 sg13g2_a21oi_1 _5589_ (.A1(_1649_),
    .A2(_1655_),
    .Y(_1656_),
    .B1(net912));
 sg13g2_a21o_1 _5590_ (.A2(_1557_),
    .A1(_1527_),
    .B1(net918),
    .X(_1657_));
 sg13g2_nor2_1 _5591_ (.A(net934),
    .B(_1505_),
    .Y(_1658_));
 sg13g2_nand2b_1 _5592_ (.Y(_1659_),
    .B(net929),
    .A_N(_1505_));
 sg13g2_nand2_1 _5593_ (.Y(_1660_),
    .A(net918),
    .B(_1659_));
 sg13g2_a21oi_1 _5594_ (.A1(net923),
    .A2(_1553_),
    .Y(_1661_),
    .B1(net929));
 sg13g2_nor2_1 _5595_ (.A(_1584_),
    .B(_1599_),
    .Y(_1662_));
 sg13g2_a221oi_1 _5596_ (.B2(_1662_),
    .C1(net909),
    .B1(_1661_),
    .A1(_1657_),
    .Y(_1663_),
    .A2(_1660_));
 sg13g2_nor4_1 _5597_ (.A(_1592_),
    .B(_1618_),
    .C(_1656_),
    .D(_1663_),
    .Y(_1664_));
 sg13g2_or4_1 _5598_ (.A(_1642_),
    .B(_1645_),
    .C(_1653_),
    .D(_1664_),
    .X(_1665_));
 sg13g2_nand3_1 _5599_ (.B(_1522_),
    .C(_1553_),
    .A(net934),
    .Y(_1666_));
 sg13g2_nand3_1 _5600_ (.B(_1563_),
    .C(_1666_),
    .A(net924),
    .Y(_1667_));
 sg13g2_a21oi_1 _5601_ (.A1(_1646_),
    .A2(_1667_),
    .Y(_1668_),
    .B1(net907));
 sg13g2_a221oi_1 _5602_ (.B2(_1543_),
    .C1(_1541_),
    .B1(_1524_),
    .A1(_1454_),
    .Y(_1669_),
    .A2(_1489_));
 sg13g2_o21ai_1 _5603_ (.B1(net935),
    .Y(_1670_),
    .A1(_1668_),
    .A2(_1669_));
 sg13g2_nand3_1 _5604_ (.B(_1508_),
    .C(_1522_),
    .A(net926),
    .Y(_1671_));
 sg13g2_nand3_1 _5605_ (.B(_1646_),
    .C(_1671_),
    .A(_1579_),
    .Y(_1672_));
 sg13g2_a21oi_1 _5606_ (.A1(net910),
    .A2(_1672_),
    .Y(_1673_),
    .B1(_1669_));
 sg13g2_or2_1 _5607_ (.X(_1674_),
    .B(_1673_),
    .A(_1599_));
 sg13g2_o21ai_1 _5608_ (.B1(_1592_),
    .Y(_1675_),
    .A1(_1581_),
    .A2(_1582_));
 sg13g2_nand4_1 _5609_ (.B(_1670_),
    .C(_1674_),
    .A(_1474_),
    .Y(_1676_),
    .D(_1675_));
 sg13g2_a21oi_1 _5610_ (.A1(_1473_),
    .A2(_1665_),
    .Y(_1677_),
    .B1(_1552_));
 sg13g2_a21oi_1 _5611_ (.A1(_1676_),
    .A2(_1677_),
    .Y(_1678_),
    .B1(_1370_));
 sg13g2_a221oi_1 _5612_ (.B2(_1678_),
    .C1(_1617_),
    .B1(_1635_),
    .A1(_1370_),
    .Y(_1679_),
    .A2(_1609_));
 sg13g2_a221oi_1 _5613_ (.B2(net928),
    .C1(net922),
    .B1(_1648_),
    .A1(net938),
    .Y(_1680_),
    .A2(_1494_));
 sg13g2_a21oi_1 _5614_ (.A1(_1485_),
    .A2(_1503_),
    .Y(_1681_),
    .B1(net918));
 sg13g2_o21ai_1 _5615_ (.B1(net909),
    .Y(_1682_),
    .A1(_1680_),
    .A2(_1681_));
 sg13g2_nand3_1 _5616_ (.B(_1571_),
    .C(_1659_),
    .A(net918),
    .Y(_1683_));
 sg13g2_a21o_1 _5617_ (.A2(_1683_),
    .A1(_1657_),
    .B1(net909),
    .X(_1684_));
 sg13g2_nand3_1 _5618_ (.B(_1682_),
    .C(_1684_),
    .A(net937),
    .Y(_1685_));
 sg13g2_nor2_1 _5619_ (.A(_1650_),
    .B(_1680_),
    .Y(_1686_));
 sg13g2_o21ai_1 _5620_ (.B1(_1505_),
    .Y(_1687_),
    .A1(_1541_),
    .A2(_1628_));
 sg13g2_a22oi_1 _5621_ (.Y(_1688_),
    .B1(_1687_),
    .B2(net922),
    .A2(_1572_),
    .A1(_1487_));
 sg13g2_a221oi_1 _5622_ (.B2(_1513_),
    .C1(net935),
    .B1(_1688_),
    .A1(_1531_),
    .Y(_1689_),
    .A2(_1686_));
 sg13g2_a221oi_1 _5623_ (.B2(_1648_),
    .C1(net909),
    .B1(_1661_),
    .A1(_1657_),
    .Y(_1690_),
    .A2(_1660_));
 sg13g2_nand3b_1 _5624_ (.B(_1512_),
    .C(_1682_),
    .Y(_1691_),
    .A_N(_1690_));
 sg13g2_nand4_1 _5625_ (.B(_1482_),
    .C(_1515_),
    .A(net932),
    .Y(_1692_),
    .D(_1522_));
 sg13g2_nand2b_1 _5626_ (.Y(_1693_),
    .B(net929),
    .A_N(_1553_));
 sg13g2_a21oi_1 _5627_ (.A1(_1692_),
    .A2(_1693_),
    .Y(_1694_),
    .B1(net922));
 sg13g2_o21ai_1 _5628_ (.B1(net912),
    .Y(_1695_),
    .A1(_1639_),
    .A2(_1694_));
 sg13g2_nor3_1 _5629_ (.A(net932),
    .B(net922),
    .C(_1648_),
    .Y(_1696_));
 sg13g2_nand3_1 _5630_ (.B(net917),
    .C(_1647_),
    .A(net928),
    .Y(_1697_));
 sg13g2_mux2_1 _5631_ (.A0(_1495_),
    .A1(_1523_),
    .S(net932),
    .X(_1698_));
 sg13g2_o21ai_1 _5632_ (.B1(net937),
    .Y(_1699_),
    .A1(net917),
    .A2(_1698_));
 sg13g2_o21ai_1 _5633_ (.B1(_1521_),
    .Y(_1700_),
    .A1(_1696_),
    .A2(_1699_));
 sg13g2_a21oi_1 _5634_ (.A1(_1695_),
    .A2(_1700_),
    .Y(_1701_),
    .B1(_1371_));
 sg13g2_a221oi_1 _5635_ (.B2(_1701_),
    .C1(_1552_),
    .B1(_1691_),
    .A1(_1685_),
    .Y(_1702_),
    .A2(_1689_));
 sg13g2_nand3_1 _5636_ (.B(_1528_),
    .C(_1592_),
    .A(_1526_),
    .Y(_1703_));
 sg13g2_a21oi_1 _5637_ (.A1(_1486_),
    .A2(_1593_),
    .Y(_1704_),
    .B1(_1494_));
 sg13g2_a21oi_1 _5638_ (.A1(_1703_),
    .A2(_1704_),
    .Y(_1705_),
    .B1(net917));
 sg13g2_a21oi_1 _5639_ (.A1(_1483_),
    .A2(net923),
    .Y(_1706_),
    .B1(net916));
 sg13g2_a22oi_1 _5640_ (.Y(_1707_),
    .B1(_1706_),
    .B2(_1564_),
    .A2(_1697_),
    .A1(net916));
 sg13g2_o21ai_1 _5641_ (.B1(net909),
    .Y(_1708_),
    .A1(_1705_),
    .A2(_1707_));
 sg13g2_o21ai_1 _5642_ (.B1(_1588_),
    .Y(_1709_),
    .A1(net922),
    .A2(_1618_));
 sg13g2_nand4_1 _5643_ (.B(_1567_),
    .C(net916),
    .A(net917),
    .Y(_1710_),
    .D(_1692_));
 sg13g2_and2_1 _5644_ (.A(net912),
    .B(_1710_),
    .X(_1711_));
 sg13g2_o21ai_1 _5645_ (.B1(_1711_),
    .Y(_1712_),
    .A1(_1546_),
    .A2(_1709_));
 sg13g2_nand3b_1 _5646_ (.B(net936),
    .C(net910),
    .Y(_1713_),
    .A_N(_1594_));
 sg13g2_and4_1 _5647_ (.A(_1552_),
    .B(_1708_),
    .C(_1712_),
    .D(_1713_),
    .X(_1714_));
 sg13g2_o21ai_1 _5648_ (.B1(net906),
    .Y(_1715_),
    .A1(_1702_),
    .A2(_1714_));
 sg13g2_a21o_1 _5649_ (.A2(_1544_),
    .A1(_1486_),
    .B1(net917),
    .X(_1716_));
 sg13g2_or3_1 _5650_ (.A(net923),
    .B(_1517_),
    .C(_1561_),
    .X(_1717_));
 sg13g2_nand2_1 _5651_ (.Y(_1718_),
    .A(_1716_),
    .B(_1717_));
 sg13g2_nand4_1 _5652_ (.B(net916),
    .C(_1716_),
    .A(net912),
    .Y(_1719_),
    .D(_1717_));
 sg13g2_nand3_1 _5653_ (.B(_1573_),
    .C(_1618_),
    .A(net912),
    .Y(_1720_));
 sg13g2_a21oi_1 _5654_ (.A1(_1719_),
    .A2(_1720_),
    .Y(_1721_),
    .B1(_1551_));
 sg13g2_a221oi_1 _5655_ (.B2(_1718_),
    .C1(net916),
    .B1(_1579_),
    .A1(_1490_),
    .Y(_1722_),
    .A2(_1491_));
 sg13g2_and2_1 _5656_ (.A(net916),
    .B(_1668_),
    .X(_1723_));
 sg13g2_o21ai_1 _5657_ (.B1(_1551_),
    .Y(_1724_),
    .A1(_1722_),
    .A2(_1723_));
 sg13g2_nor3_1 _5658_ (.A(net906),
    .B(_1568_),
    .C(_1721_),
    .Y(_1725_));
 sg13g2_a21oi_1 _5659_ (.A1(_1724_),
    .A2(_1725_),
    .Y(_1726_),
    .B1(_1370_));
 sg13g2_o21ai_1 _5660_ (.B1(net920),
    .Y(_1727_),
    .A1(_1503_),
    .A2(_1561_));
 sg13g2_a21oi_1 _5661_ (.A1(_1629_),
    .A2(_1727_),
    .Y(_1728_),
    .B1(net910));
 sg13g2_nor2_1 _5662_ (.A(net925),
    .B(_1666_),
    .Y(_1729_));
 sg13g2_a22oi_1 _5663_ (.Y(_1730_),
    .B1(_1729_),
    .B2(net910),
    .A2(_1604_),
    .A1(_1601_));
 sg13g2_nand3_1 _5664_ (.B(_1507_),
    .C(_1621_),
    .A(net910),
    .Y(_1731_));
 sg13g2_a21oi_1 _5665_ (.A1(_1601_),
    .A2(_1622_),
    .Y(_1732_),
    .B1(_1599_));
 sg13g2_a22oi_1 _5666_ (.Y(_1733_),
    .B1(_1731_),
    .B2(_1732_),
    .A2(_1730_),
    .A1(net936));
 sg13g2_nand3_1 _5667_ (.B(_1623_),
    .C(_1727_),
    .A(_1531_),
    .Y(_1734_));
 sg13g2_mux2_1 _5668_ (.A0(_1524_),
    .A1(_1658_),
    .S(net920),
    .X(_1735_));
 sg13g2_or3_1 _5669_ (.A(_1514_),
    .B(_1729_),
    .C(_1735_),
    .X(_1736_));
 sg13g2_a21o_1 _5670_ (.A2(_1736_),
    .A1(_1734_),
    .B1(net936),
    .X(_1737_));
 sg13g2_o21ai_1 _5671_ (.B1(_1737_),
    .Y(_1738_),
    .A1(_1728_),
    .A2(_1733_));
 sg13g2_nand2_1 _5672_ (.Y(_1739_),
    .A(_1474_),
    .B(_1499_));
 sg13g2_o21ai_1 _5673_ (.B1(_1370_),
    .Y(_1740_),
    .A1(_1581_),
    .A2(_1739_));
 sg13g2_a21oi_1 _5674_ (.A1(_1473_),
    .A2(_1738_),
    .Y(_1741_),
    .B1(_1740_));
 sg13g2_a21o_1 _5675_ (.A2(_1726_),
    .A1(_1715_),
    .B1(_1741_),
    .X(_1742_));
 sg13g2_a21oi_1 _5676_ (.A1(_1455_),
    .A2(_1472_),
    .Y(_1743_),
    .B1(_1471_));
 sg13g2_xnor2_1 _5677_ (.Y(_1744_),
    .A(net1070),
    .B(_1043_));
 sg13g2_nor2_1 _5678_ (.A(_1458_),
    .B(_1744_),
    .Y(_1745_));
 sg13g2_a21oi_1 _5679_ (.A1(_1035_),
    .A2(_1044_),
    .Y(_1746_),
    .B1(_1382_));
 sg13g2_xor2_1 _5680_ (.B(_1746_),
    .A(_1745_),
    .X(_1747_));
 sg13g2_a21oi_1 _5681_ (.A1(_1428_),
    .A2(_1747_),
    .Y(_1748_),
    .B1(net993));
 sg13g2_nor2_1 _5682_ (.A(_1461_),
    .B(_1463_),
    .Y(_1749_));
 sg13g2_nor3_1 _5683_ (.A(_1035_),
    .B(_1200_),
    .C(_1749_),
    .Y(_1750_));
 sg13g2_a21oi_1 _5684_ (.A1(net1069),
    .A2(_1460_),
    .Y(_1751_),
    .B1(_1750_));
 sg13g2_nor2b_1 _5685_ (.A(_1751_),
    .B_N(net993),
    .Y(_1752_));
 sg13g2_nor3_2 _5686_ (.A(_1381_),
    .B(_1748_),
    .C(_1752_),
    .Y(_1753_));
 sg13g2_or3_1 _5687_ (.A(\vgademo.h_count[10] ),
    .B(_3195_),
    .C(_1468_),
    .X(_1754_));
 sg13g2_nand3_1 _5688_ (.B(net952),
    .C(_1754_),
    .A(_0060_),
    .Y(_1755_));
 sg13g2_o21ai_1 _5689_ (.B1(_1755_),
    .Y(_1756_),
    .A1(_3267_),
    .A2(net952));
 sg13g2_xor2_1 _5690_ (.B(_1756_),
    .A(_1753_),
    .X(_1757_));
 sg13g2_inv_1 _5691_ (.Y(_1758_),
    .A(_1757_));
 sg13g2_xor2_1 _5692_ (.B(_1749_),
    .A(net1070),
    .X(_1759_));
 sg13g2_xnor2_1 _5693_ (.Y(_1760_),
    .A(_1457_),
    .B(_1744_));
 sg13g2_a221oi_1 _5694_ (.B2(_1386_),
    .C1(_1387_),
    .B1(_1760_),
    .A1(net993),
    .Y(_1761_),
    .A2(_1759_));
 sg13g2_o21ai_1 _5695_ (.B1(\vgademo.h_count[10] ),
    .Y(_1762_),
    .A1(_3195_),
    .A2(_1468_));
 sg13g2_nand3_1 _5696_ (.B(_1754_),
    .C(_1762_),
    .A(net952),
    .Y(_1763_));
 sg13g2_o21ai_1 _5697_ (.B1(_1763_),
    .Y(_1764_),
    .A1(_0031_),
    .A2(net952));
 sg13g2_nand2_1 _5698_ (.Y(_1765_),
    .A(_1761_),
    .B(_1764_));
 sg13g2_o21ai_1 _5699_ (.B1(_1765_),
    .Y(_1766_),
    .A1(_1743_),
    .A2(_1757_));
 sg13g2_o21ai_1 _5700_ (.B1(_1758_),
    .Y(_1767_),
    .A1(_1761_),
    .A2(_1764_));
 sg13g2_nand2b_1 _5701_ (.Y(_1768_),
    .B(_1767_),
    .A_N(_1743_));
 sg13g2_mux2_1 _5702_ (.A0(_1767_),
    .A1(_1768_),
    .S(_1766_),
    .X(_1769_));
 sg13g2_a21o_1 _5703_ (.A2(_1742_),
    .A1(_1617_),
    .B1(_1769_),
    .X(_1770_));
 sg13g2_xnor2_1 _5704_ (.Y(_1771_),
    .A(net1055),
    .B(net1054));
 sg13g2_nand2_1 _5705_ (.Y(_1772_),
    .A(\vgademo.v_count[5] ),
    .B(_1771_));
 sg13g2_nand2_1 _5706_ (.Y(_1773_),
    .A(net1064),
    .B(_3237_));
 sg13g2_nand2b_1 _5707_ (.Y(_1774_),
    .B(\vgademo.b_cos[8] ),
    .A_N(net1064));
 sg13g2_o21ai_1 _5708_ (.B1(_3183_),
    .Y(_1775_),
    .A1(net1056),
    .A2(_1354_));
 sg13g2_a22oi_1 _5709_ (.Y(_1776_),
    .B1(_1356_),
    .B2(_1775_),
    .A2(_3235_),
    .A1(net1065));
 sg13g2_o21ai_1 _5710_ (.B1(_1774_),
    .Y(_1777_),
    .A1(\vgademo.v_count[2] ),
    .A2(_3235_));
 sg13g2_o21ai_1 _5711_ (.B1(_1773_),
    .Y(_1778_),
    .A1(_1776_),
    .A2(_1777_));
 sg13g2_a21oi_1 _5712_ (.A1(net1062),
    .A2(_1778_),
    .Y(_1779_),
    .B1(net1055));
 sg13g2_xnor2_1 _5713_ (.Y(_1780_),
    .A(_0062_),
    .B(_1771_));
 sg13g2_o21ai_1 _5714_ (.B1(_1780_),
    .Y(_1781_),
    .A1(net1062),
    .A2(_1778_));
 sg13g2_o21ai_1 _5715_ (.B1(_1772_),
    .Y(_1782_),
    .A1(_1779_),
    .A2(_1781_));
 sg13g2_nor2_1 _5716_ (.A(net1055),
    .B(\vgademo.b_cos[11] ),
    .Y(_1783_));
 sg13g2_a21oi_2 _5717_ (.B1(_1783_),
    .Y(_1784_),
    .A2(_1612_),
    .A1(net1055));
 sg13g2_xnor2_1 _5718_ (.Y(_1785_),
    .A(_0016_),
    .B(_1784_));
 sg13g2_and2_1 _5719_ (.A(net1061),
    .B(_1784_),
    .X(_1786_));
 sg13g2_a221oi_1 _5720_ (.B2(_1785_),
    .C1(_1786_),
    .B1(_1782_),
    .A1(net1060),
    .Y(_1787_),
    .A2(_3213_));
 sg13g2_or2_2 _5721_ (.X(_1788_),
    .B(_1611_),
    .A(_3238_));
 sg13g2_nand3_1 _5722_ (.B(_0018_),
    .C(_1788_),
    .A(net1060),
    .Y(_1789_));
 sg13g2_o21ai_1 _5723_ (.B1(_1789_),
    .Y(_1790_),
    .A1(_0018_),
    .A2(_1788_));
 sg13g2_nand2b_1 _5724_ (.Y(_1791_),
    .B(_1790_),
    .A_N(_1787_));
 sg13g2_o21ai_1 _5725_ (.B1(_3238_),
    .Y(_1792_),
    .A1(net1062),
    .A2(_1778_));
 sg13g2_a22oi_1 _5726_ (.Y(_1793_),
    .B1(_1778_),
    .B2(net1062),
    .A2(net1054),
    .A1(\vgademo.v_count[5] ));
 sg13g2_xnor2_1 _5727_ (.Y(_1794_),
    .A(_0016_),
    .B(_1612_));
 sg13g2_a221oi_1 _5728_ (.B2(_1793_),
    .C1(_1794_),
    .B1(_1792_),
    .A1(_3185_),
    .Y(_1795_),
    .A2(_3239_));
 sg13g2_a221oi_1 _5729_ (.B2(net1061),
    .C1(_1795_),
    .B1(_1613_),
    .A1(net1060),
    .Y(_1796_),
    .A2(_1611_));
 sg13g2_o21ai_1 _5730_ (.B1(_0018_),
    .Y(_1797_),
    .A1(net1060),
    .A2(_1611_));
 sg13g2_o21ai_1 _5731_ (.B1(_0021_),
    .Y(_1798_),
    .A1(_1796_),
    .A2(_1797_));
 sg13g2_nand2_1 _5732_ (.Y(_1799_),
    .A(_3312_),
    .B(_1798_));
 sg13g2_o21ai_1 _5733_ (.B1(_1799_),
    .Y(_1800_),
    .A1(_3315_),
    .A2(_1788_));
 sg13g2_nand2_2 _5734_ (.Y(_1801_),
    .A(_1791_),
    .B(_1800_));
 sg13g2_nor3_2 _5735_ (.A(net903),
    .B(net900),
    .C(_1801_),
    .Y(_1802_));
 sg13g2_or3_1 _5736_ (.A(net903),
    .B(net900),
    .C(_1801_),
    .X(_1803_));
 sg13g2_nand2_1 _5737_ (.Y(_1804_),
    .A(\vgademo.plane_du[8] ),
    .B(_1784_));
 sg13g2_xnor2_1 _5738_ (.Y(_1805_),
    .A(_0052_),
    .B(_1771_));
 sg13g2_o21ai_1 _5739_ (.B1(_3247_),
    .Y(_1806_),
    .A1(net1056),
    .A2(_1350_));
 sg13g2_a22oi_1 _5740_ (.Y(_1807_),
    .B1(_1351_),
    .B2(_1806_),
    .A2(\vgademo.plane_du[4] ),
    .A1(_3235_));
 sg13g2_a221oi_1 _5741_ (.B2(\vgademo.b_cos[8] ),
    .C1(_1807_),
    .B1(_3250_),
    .A1(\vgademo.b_cos[7] ),
    .Y(_1808_),
    .A2(_3248_));
 sg13g2_a21oi_1 _5742_ (.A1(_3237_),
    .A2(\vgademo.plane_du[5] ),
    .Y(_1809_),
    .B1(_1808_));
 sg13g2_nor2b_1 _5743_ (.A(_1809_),
    .B_N(\vgademo.plane_du[6] ),
    .Y(_1810_));
 sg13g2_nand2b_1 _5744_ (.Y(_1811_),
    .B(_1809_),
    .A_N(\vgademo.plane_du[6] ));
 sg13g2_a21o_1 _5745_ (.A2(_1811_),
    .A1(net1055),
    .B1(_1810_),
    .X(_1812_));
 sg13g2_a22oi_1 _5746_ (.Y(_1813_),
    .B1(_1805_),
    .B2(_1812_),
    .A2(_1771_),
    .A1(\vgademo.plane_du[7] ));
 sg13g2_xor2_1 _5747_ (.B(_1784_),
    .A(_0053_),
    .X(_1814_));
 sg13g2_o21ai_1 _5748_ (.B1(_1804_),
    .Y(_1815_),
    .A1(_1813_),
    .A2(_1814_));
 sg13g2_nand3_1 _5749_ (.B(_1788_),
    .C(_1815_),
    .A(\vgademo.plane_du[9] ),
    .Y(_1816_));
 sg13g2_a221oi_1 _5750_ (.B2(_3238_),
    .C1(_1810_),
    .B1(_1811_),
    .A1(net1054),
    .Y(_1817_),
    .A2(\vgademo.plane_du[7] ));
 sg13g2_xnor2_1 _5751_ (.Y(_1818_),
    .A(_0053_),
    .B(_1613_));
 sg13g2_o21ai_1 _5752_ (.B1(_1818_),
    .Y(_1819_),
    .A1(net1054),
    .A2(\vgademo.plane_du[7] ));
 sg13g2_a22oi_1 _5753_ (.Y(_1820_),
    .B1(_1613_),
    .B2(\vgademo.plane_du[8] ),
    .A2(_1611_),
    .A1(\vgademo.plane_du[9] ));
 sg13g2_o21ai_1 _5754_ (.B1(_1820_),
    .Y(_1821_),
    .A1(_1817_),
    .A2(_1819_));
 sg13g2_o21ai_1 _5755_ (.B1(_1821_),
    .Y(_1822_),
    .A1(\vgademo.plane_du[9] ),
    .A2(_1611_));
 sg13g2_nand2b_2 _5756_ (.Y(_1823_),
    .B(_1816_),
    .A_N(_1822_));
 sg13g2_nor3_2 _5757_ (.A(net902),
    .B(net899),
    .C(net947),
    .Y(_1824_));
 sg13g2_or3_1 _5758_ (.A(net904),
    .B(net901),
    .C(net948),
    .X(_1825_));
 sg13g2_nand2_1 _5759_ (.Y(_1826_),
    .A(net1087),
    .B(\vgademo.plane_du[5] ));
 sg13g2_and2_1 _5760_ (.A(net1091),
    .B(\vgademo.plane_du[4] ),
    .X(_1827_));
 sg13g2_nand2_1 _5761_ (.Y(_1828_),
    .A(_3201_),
    .B(_3250_));
 sg13g2_nand3_1 _5762_ (.B(_1827_),
    .C(_1828_),
    .A(_1826_),
    .Y(_1829_));
 sg13g2_xnor2_1 _5763_ (.Y(_1830_),
    .A(net1084),
    .B(\vgademo.plane_du[6] ));
 sg13g2_a21oi_1 _5764_ (.A1(_1826_),
    .A2(_1829_),
    .Y(_1831_),
    .B1(_1830_));
 sg13g2_a21oi_1 _5765_ (.A1(net1084),
    .A2(\vgademo.plane_du[6] ),
    .Y(_1832_),
    .B1(_1831_));
 sg13g2_xor2_1 _5766_ (.B(\vgademo.plane_du[7] ),
    .A(net1081),
    .X(_1833_));
 sg13g2_nand2b_1 _5767_ (.Y(_1834_),
    .B(_1833_),
    .A_N(_1832_));
 sg13g2_xnor2_1 _5768_ (.Y(_1835_),
    .A(_1832_),
    .B(_1833_));
 sg13g2_nand2_1 _5769_ (.Y(_1836_),
    .A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ));
 sg13g2_nor2_1 _5770_ (.A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ),
    .Y(_1837_));
 sg13g2_xor2_1 _5771_ (.B(\vgademo.plane_u[15] ),
    .A(\vgademo.a_cos[10] ),
    .X(_1838_));
 sg13g2_nand2_1 _5772_ (.Y(_1839_),
    .A(\vgademo.a_cos[8] ),
    .B(\vgademo.plane_u[13] ));
 sg13g2_and2_1 _5773_ (.A(\vgademo.a_cos[7] ),
    .B(\vgademo.plane_u[12] ),
    .X(_1840_));
 sg13g2_xor2_1 _5774_ (.B(\vgademo.plane_u[12] ),
    .A(\vgademo.a_cos[7] ),
    .X(_1841_));
 sg13g2_or2_1 _5775_ (.X(_1842_),
    .B(\vgademo.plane_u[10] ),
    .A(\vgademo.a_cos[5] ));
 sg13g2_nand3_1 _5776_ (.B(\vgademo.plane_u[9] ),
    .C(_1842_),
    .A(\vgademo.a_cos[4] ),
    .Y(_1843_));
 sg13g2_a22oi_1 _5777_ (.Y(_1844_),
    .B1(\vgademo.plane_u[11] ),
    .B2(\vgademo.a_cos[6] ),
    .A2(\vgademo.plane_u[10] ),
    .A1(\vgademo.a_cos[5] ));
 sg13g2_a22oi_1 _5778_ (.Y(_1845_),
    .B1(_1843_),
    .B2(_1844_),
    .A2(_3261_),
    .A1(_3231_));
 sg13g2_a21oi_1 _5779_ (.A1(_1841_),
    .A2(_1845_),
    .Y(_1846_),
    .B1(_1840_));
 sg13g2_nor2_1 _5780_ (.A(\vgademo.a_cos[8] ),
    .B(\vgademo.plane_u[13] ),
    .Y(_1847_));
 sg13g2_xor2_1 _5781_ (.B(\vgademo.plane_u[13] ),
    .A(\vgademo.a_cos[8] ),
    .X(_1848_));
 sg13g2_o21ai_1 _5782_ (.B1(_1839_),
    .Y(_1849_),
    .A1(_1846_),
    .A2(_1847_));
 sg13g2_a21o_1 _5783_ (.A2(\vgademo.plane_u[14] ),
    .A1(\vgademo.a_cos[9] ),
    .B1(_1849_),
    .X(_1850_));
 sg13g2_o21ai_1 _5784_ (.B1(_1850_),
    .Y(_1851_),
    .A1(\vgademo.a_cos[9] ),
    .A2(\vgademo.plane_u[14] ));
 sg13g2_o21ai_1 _5785_ (.B1(_1836_),
    .Y(_1852_),
    .A1(_1837_),
    .A2(_1851_));
 sg13g2_and2_1 _5786_ (.A(\vgademo.a_cos[11] ),
    .B(\vgademo.plane_u[16] ),
    .X(_1853_));
 sg13g2_xor2_1 _5787_ (.B(\vgademo.plane_u[16] ),
    .A(\vgademo.a_cos[11] ),
    .X(_1854_));
 sg13g2_xnor2_1 _5788_ (.Y(_1855_),
    .A(_1852_),
    .B(_1854_));
 sg13g2_inv_1 _5789_ (.Y(_1856_),
    .A(_1855_));
 sg13g2_nor2_1 _5790_ (.A(_1835_),
    .B(_1855_),
    .Y(_1857_));
 sg13g2_xor2_1 _5791_ (.B(_1855_),
    .A(_1835_),
    .X(_1858_));
 sg13g2_o21ai_1 _5792_ (.B1(_1834_),
    .Y(_1859_),
    .A1(_3200_),
    .A2(_3254_));
 sg13g2_xor2_1 _5793_ (.B(\vgademo.plane_du[8] ),
    .A(net1078),
    .X(_1860_));
 sg13g2_nand2_1 _5794_ (.Y(_1861_),
    .A(_1859_),
    .B(_1860_));
 sg13g2_xnor2_1 _5795_ (.Y(_1862_),
    .A(_1859_),
    .B(_1860_));
 sg13g2_nor2_1 _5796_ (.A(_1858_),
    .B(_1862_),
    .Y(_1863_));
 sg13g2_o21ai_1 _5797_ (.B1(_0074_),
    .Y(_1864_),
    .A1(_1204_),
    .A2(_1378_));
 sg13g2_a21oi_1 _5798_ (.A1(_1066_),
    .A2(_1864_),
    .Y(_1865_),
    .B1(_1068_));
 sg13g2_nor2_1 _5799_ (.A(_1064_),
    .B(_1865_),
    .Y(_1866_));
 sg13g2_o21ai_1 _5800_ (.B1(_1861_),
    .Y(_1867_),
    .A1(net1045),
    .A2(_3256_));
 sg13g2_nor2_1 _5801_ (.A(_3198_),
    .B(_3259_),
    .Y(_1868_));
 sg13g2_xor2_1 _5802_ (.B(\vgademo.plane_du[9] ),
    .A(net1076),
    .X(_1869_));
 sg13g2_xnor2_1 _5803_ (.Y(_1870_),
    .A(_1867_),
    .B(_1869_));
 sg13g2_and2_1 _5804_ (.A(\vgademo.a_cos[12] ),
    .B(\vgademo.plane_u[17] ),
    .X(_1871_));
 sg13g2_a21o_1 _5805_ (.A2(_1854_),
    .A1(_1852_),
    .B1(_1853_),
    .X(_1872_));
 sg13g2_xor2_1 _5806_ (.B(\vgademo.plane_u[17] ),
    .A(\vgademo.a_cos[12] ),
    .X(_1873_));
 sg13g2_a21o_1 _5807_ (.A2(_1873_),
    .A1(_1872_),
    .B1(_1871_),
    .X(_1874_));
 sg13g2_xor2_1 _5808_ (.B(\vgademo.plane_u[18] ),
    .A(\vgademo.a_cos[13] ),
    .X(_1875_));
 sg13g2_xnor2_1 _5809_ (.Y(_1876_),
    .A(_1874_),
    .B(_1875_));
 sg13g2_nor2_1 _5810_ (.A(_1870_),
    .B(_1876_),
    .Y(_1877_));
 sg13g2_nand2_1 _5811_ (.Y(_1878_),
    .A(_1870_),
    .B(_1876_));
 sg13g2_nand2b_1 _5812_ (.Y(_1879_),
    .B(_1878_),
    .A_N(_1877_));
 sg13g2_xnor2_1 _5813_ (.Y(_1880_),
    .A(_1872_),
    .B(_1873_));
 sg13g2_xor2_1 _5814_ (.B(_1880_),
    .A(_1862_),
    .X(_1881_));
 sg13g2_nand3_1 _5815_ (.B(_1856_),
    .C(_1881_),
    .A(_1835_),
    .Y(_1882_));
 sg13g2_o21ai_1 _5816_ (.B1(_1882_),
    .Y(_1883_),
    .A1(_1862_),
    .A2(_1880_));
 sg13g2_a21oi_1 _5817_ (.A1(_1878_),
    .A2(_1883_),
    .Y(_1884_),
    .B1(_1877_));
 sg13g2_a21o_1 _5818_ (.A2(\vgademo.plane_u[18] ),
    .A1(\vgademo.a_cos[13] ),
    .B1(_1874_),
    .X(_1885_));
 sg13g2_o21ai_1 _5819_ (.B1(_1885_),
    .Y(_1886_),
    .A1(\vgademo.a_cos[13] ),
    .A2(\vgademo.plane_u[18] ));
 sg13g2_a21oi_1 _5820_ (.A1(_1867_),
    .A2(_1869_),
    .Y(_1887_),
    .B1(_1868_));
 sg13g2_xor2_1 _5821_ (.B(\vgademo.a_cos[14] ),
    .A(net1073),
    .X(_1888_));
 sg13g2_xor2_1 _5822_ (.B(\vgademo.plane_u[19] ),
    .A(\vgademo.plane_du[10] ),
    .X(_1889_));
 sg13g2_xnor2_1 _5823_ (.Y(_1890_),
    .A(_1888_),
    .B(_1889_));
 sg13g2_xnor2_1 _5824_ (.Y(_1891_),
    .A(_1887_),
    .B(_1890_));
 sg13g2_xnor2_1 _5825_ (.Y(_1892_),
    .A(_1886_),
    .B(_1891_));
 sg13g2_xnor2_1 _5826_ (.Y(_1893_),
    .A(_1884_),
    .B(_1892_));
 sg13g2_xor2_1 _5827_ (.B(_1883_),
    .A(_1879_),
    .X(_1894_));
 sg13g2_nor2_1 _5828_ (.A(net1146),
    .B(_1858_),
    .Y(_1895_));
 sg13g2_nand2b_1 _5829_ (.Y(_1896_),
    .B(net1143),
    .A_N(_1881_));
 sg13g2_a21o_1 _5830_ (.A2(_1856_),
    .A1(_1835_),
    .B1(_1881_),
    .X(_1897_));
 sg13g2_and2_1 _5831_ (.A(net1049),
    .B(_1882_),
    .X(_1898_));
 sg13g2_a22oi_1 _5832_ (.Y(_1899_),
    .B1(_1897_),
    .B2(_1898_),
    .A2(_1896_),
    .A1(_1895_));
 sg13g2_o21ai_1 _5833_ (.B1(_1899_),
    .Y(_1900_),
    .A1(\vgademo.audio_songpos[4] ),
    .A2(_1894_));
 sg13g2_inv_1 _5834_ (.Y(_1901_),
    .A(_1900_));
 sg13g2_a221oi_1 _5835_ (.B2(\vgademo.audio_songpos[4] ),
    .C1(_1901_),
    .B1(_1894_),
    .A1(net1136),
    .Y(_1902_),
    .A2(_1893_));
 sg13g2_nor2_1 _5836_ (.A(net1136),
    .B(_1893_),
    .Y(_1903_));
 sg13g2_nor3_2 _5837_ (.A(_3383_),
    .B(_1902_),
    .C(_1903_),
    .Y(_1904_));
 sg13g2_or2_2 _5838_ (.X(_1905_),
    .B(_1904_),
    .A(_1866_));
 sg13g2_xnor2_1 _5839_ (.Y(_1906_),
    .A(_3170_),
    .B(_1879_));
 sg13g2_and2_1 _5840_ (.A(net1049),
    .B(_1835_),
    .X(_1907_));
 sg13g2_o21ai_1 _5841_ (.B1(net1131),
    .Y(_1908_),
    .A1(net1049),
    .A2(_1835_));
 sg13g2_xnor2_1 _5842_ (.Y(_1909_),
    .A(net1149),
    .B(_1855_));
 sg13g2_nor3_1 _5843_ (.A(_1907_),
    .B(_1908_),
    .C(_1909_),
    .Y(_1910_));
 sg13g2_xnor2_1 _5844_ (.Y(_1911_),
    .A(net1146),
    .B(_1881_));
 sg13g2_nand3_1 _5845_ (.B(_1910_),
    .C(_1911_),
    .A(_1906_),
    .Y(_1912_));
 sg13g2_nand2b_2 _5846_ (.Y(_1913_),
    .B(_1912_),
    .A_N(_1905_));
 sg13g2_inv_1 _5847_ (.Y(_1914_),
    .A(net905));
 sg13g2_or2_1 _5848_ (.X(_1915_),
    .B(_1913_),
    .A(_1863_));
 sg13g2_and2_1 _5849_ (.A(net955),
    .B(_1915_),
    .X(_1916_));
 sg13g2_nand2_1 _5850_ (.Y(_1917_),
    .A(net1156),
    .B(net1077));
 sg13g2_nand2_1 _5851_ (.Y(_1918_),
    .A(net1080),
    .B(net1153));
 sg13g2_nand2_1 _5852_ (.Y(_1919_),
    .A(net1077),
    .B(net1154));
 sg13g2_nand2_1 _5853_ (.Y(_1920_),
    .A(net1156),
    .B(net1080));
 sg13g2_xor2_1 _5854_ (.B(_1920_),
    .A(_1919_),
    .X(_1921_));
 sg13g2_nand2_1 _5855_ (.Y(_1922_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1921_));
 sg13g2_o21ai_1 _5856_ (.B1(_1922_),
    .Y(_1923_),
    .A1(_1919_),
    .A2(_1920_));
 sg13g2_nand2_1 _5857_ (.Y(_1924_),
    .A(net1156),
    .B(net1075));
 sg13g2_nand2_1 _5858_ (.Y(_1925_),
    .A(net1075),
    .B(net1154));
 sg13g2_xor2_1 _5859_ (.B(_1925_),
    .A(_1917_),
    .X(_1926_));
 sg13g2_nand2_1 _5860_ (.Y(_1927_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1926_));
 sg13g2_xnor2_1 _5861_ (.Y(_1928_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1926_));
 sg13g2_nor2b_1 _5862_ (.A(_1928_),
    .B_N(_1923_),
    .Y(_1929_));
 sg13g2_nand2b_1 _5863_ (.Y(_1930_),
    .B(_1928_),
    .A_N(_1923_));
 sg13g2_nand2b_1 _5864_ (.Y(_1931_),
    .B(_1930_),
    .A_N(_1929_));
 sg13g2_a21o_1 _5865_ (.A2(_1930_),
    .A1(net1072),
    .B1(_1929_),
    .X(_1932_));
 sg13g2_o21ai_1 _5866_ (.B1(_1927_),
    .Y(_1933_),
    .A1(_1917_),
    .A2(_1925_));
 sg13g2_nand2_1 _5867_ (.Y(_1934_),
    .A(net1072),
    .B(net1154));
 sg13g2_xor2_1 _5868_ (.B(_1934_),
    .A(_1924_),
    .X(_1935_));
 sg13g2_nand2_1 _5869_ (.Y(_1936_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1935_));
 sg13g2_xnor2_1 _5870_ (.Y(_1937_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1935_));
 sg13g2_nand2b_1 _5871_ (.Y(_1938_),
    .B(_1933_),
    .A_N(_1937_));
 sg13g2_xor2_1 _5872_ (.B(_1937_),
    .A(_1933_),
    .X(_1939_));
 sg13g2_xnor2_1 _5873_ (.Y(_1940_),
    .A(_3197_),
    .B(_1939_));
 sg13g2_inv_1 _5874_ (.Y(_1941_),
    .A(_1940_));
 sg13g2_xor2_1 _5875_ (.B(_1940_),
    .A(_1932_),
    .X(_1942_));
 sg13g2_nand2_1 _5876_ (.Y(_1943_),
    .A(net1155),
    .B(net1082));
 sg13g2_xor2_1 _5877_ (.B(_1943_),
    .A(_1918_),
    .X(_1944_));
 sg13g2_nand2_1 _5878_ (.Y(_1945_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1944_));
 sg13g2_o21ai_1 _5879_ (.B1(_1945_),
    .Y(_1946_),
    .A1(_1918_),
    .A2(_1943_));
 sg13g2_xnor2_1 _5880_ (.Y(_1947_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1921_));
 sg13g2_nand2b_1 _5881_ (.Y(_1948_),
    .B(_1946_),
    .A_N(_1947_));
 sg13g2_xor2_1 _5882_ (.B(_1947_),
    .A(_1946_),
    .X(_1949_));
 sg13g2_o21ai_1 _5883_ (.B1(_1948_),
    .Y(_1950_),
    .A1(_3198_),
    .A2(_1949_));
 sg13g2_xor2_1 _5884_ (.B(_1931_),
    .A(net1073),
    .X(_1951_));
 sg13g2_nor2b_1 _5885_ (.A(_1950_),
    .B_N(_1951_),
    .Y(_1952_));
 sg13g2_nand2b_1 _5886_ (.Y(_1953_),
    .B(_1950_),
    .A_N(_1951_));
 sg13g2_and4_1 _5887_ (.A(net1155),
    .B(net1082),
    .C(net1085),
    .D(net1152),
    .X(_1954_));
 sg13g2_nand4_1 _5888_ (.B(net1082),
    .C(net1085),
    .A(net1155),
    .Y(_1955_),
    .D(net1152));
 sg13g2_a22oi_1 _5889_ (.Y(_1956_),
    .B1(net1152),
    .B2(net1082),
    .A2(net1085),
    .A1(net1155));
 sg13g2_nand3b_1 _5890_ (.B(\vgademo.linelfsr[6] ),
    .C(_1955_),
    .Y(_1957_),
    .A_N(_1956_));
 sg13g2_nand2_1 _5891_ (.Y(_1958_),
    .A(_1955_),
    .B(_1957_));
 sg13g2_xnor2_1 _5892_ (.Y(_1959_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1944_));
 sg13g2_nand2b_1 _5893_ (.Y(_1960_),
    .B(_1958_),
    .A_N(_1959_));
 sg13g2_xor2_1 _5894_ (.B(_1959_),
    .A(_1958_),
    .X(_1961_));
 sg13g2_o21ai_1 _5895_ (.B1(_1960_),
    .Y(_1962_),
    .A1(net1045),
    .A2(_1961_));
 sg13g2_xnor2_1 _5896_ (.Y(_1963_),
    .A(_3198_),
    .B(_1949_));
 sg13g2_nor2b_1 _5897_ (.A(_1963_),
    .B_N(_1962_),
    .Y(_1964_));
 sg13g2_xor2_1 _5898_ (.B(_1963_),
    .A(_1962_),
    .X(_1965_));
 sg13g2_inv_1 _5899_ (.Y(_1966_),
    .A(_1965_));
 sg13g2_and4_1 _5900_ (.A(net1155),
    .B(net1088),
    .C(net1085),
    .D(net1152),
    .X(_1967_));
 sg13g2_nand4_1 _5901_ (.B(net1088),
    .C(net1085),
    .A(net1155),
    .Y(_1968_),
    .D(net1152));
 sg13g2_a22oi_1 _5902_ (.Y(_1969_),
    .B1(net1085),
    .B2(net1152),
    .A2(net1088),
    .A1(net1155));
 sg13g2_nand3b_1 _5903_ (.B(\vgademo.linelfsr[5] ),
    .C(_1968_),
    .Y(_1970_),
    .A_N(_1969_));
 sg13g2_nand2_1 _5904_ (.Y(_1971_),
    .A(_1968_),
    .B(_1970_));
 sg13g2_o21ai_1 _5905_ (.B1(_3168_),
    .Y(_1972_),
    .A1(_1954_),
    .A2(_1956_));
 sg13g2_nand2_1 _5906_ (.Y(_1973_),
    .A(_1957_),
    .B(_1972_));
 sg13g2_nand2b_1 _5907_ (.Y(_1974_),
    .B(_1971_),
    .A_N(_1973_));
 sg13g2_xor2_1 _5908_ (.B(_1973_),
    .A(_1971_),
    .X(_1975_));
 sg13g2_o21ai_1 _5909_ (.B1(_1974_),
    .Y(_1976_),
    .A1(_3200_),
    .A2(_1975_));
 sg13g2_xnor2_1 _5910_ (.Y(_1977_),
    .A(net1045),
    .B(_1961_));
 sg13g2_nor2b_1 _5911_ (.A(_1976_),
    .B_N(_1977_),
    .Y(_1978_));
 sg13g2_nand2b_1 _5912_ (.Y(_1979_),
    .B(_1976_),
    .A_N(_1977_));
 sg13g2_and3_1 _5913_ (.X(_1980_),
    .A(net1088),
    .B(net1153),
    .C(\vgademo.linelfsr[4] ));
 sg13g2_nand3_1 _5914_ (.B(net1152),
    .C(\vgademo.linelfsr[4] ),
    .A(net1088),
    .Y(_1981_));
 sg13g2_a21oi_1 _5915_ (.A1(net1088),
    .A2(net1152),
    .Y(_1982_),
    .B1(\vgademo.linelfsr[4] ));
 sg13g2_nor2_1 _5916_ (.A(_1980_),
    .B(_1982_),
    .Y(_1983_));
 sg13g2_o21ai_1 _5917_ (.B1(_1981_),
    .Y(_1984_),
    .A1(_3201_),
    .A2(_1982_));
 sg13g2_o21ai_1 _5918_ (.B1(_3268_),
    .Y(_1985_),
    .A1(_1967_),
    .A2(_1969_));
 sg13g2_and3_1 _5919_ (.X(_1986_),
    .A(_1970_),
    .B(_1984_),
    .C(_1985_));
 sg13g2_a21oi_1 _5920_ (.A1(_1970_),
    .A2(_1985_),
    .Y(_1987_),
    .B1(_1984_));
 sg13g2_nor2_1 _5921_ (.A(_1986_),
    .B(_1987_),
    .Y(_1988_));
 sg13g2_a21o_1 _5922_ (.A2(_1988_),
    .A1(\vgademo.a_scrolly[5] ),
    .B1(_1986_),
    .X(_1989_));
 sg13g2_xnor2_1 _5923_ (.Y(_1990_),
    .A(net1081),
    .B(_1975_));
 sg13g2_and2_1 _5924_ (.A(_1989_),
    .B(_1990_),
    .X(_1991_));
 sg13g2_xnor2_1 _5925_ (.Y(_1992_),
    .A(net1082),
    .B(_1988_));
 sg13g2_xnor2_1 _5926_ (.Y(_1993_),
    .A(net1087),
    .B(_1983_));
 sg13g2_nand2_1 _5927_ (.Y(_1994_),
    .A(\vgademo.linelfsr[3] ),
    .B(net1089));
 sg13g2_nor2_1 _5928_ (.A(_1993_),
    .B(_1994_),
    .Y(_1995_));
 sg13g2_nor2b_1 _5929_ (.A(_1992_),
    .B_N(_1995_),
    .Y(_1996_));
 sg13g2_or2_1 _5930_ (.X(_1997_),
    .B(_1990_),
    .A(_1989_));
 sg13g2_nand2b_1 _5931_ (.Y(_1998_),
    .B(_1997_),
    .A_N(_1991_));
 sg13g2_a21oi_1 _5932_ (.A1(_1996_),
    .A2(_1997_),
    .Y(_1999_),
    .B1(_1991_));
 sg13g2_o21ai_1 _5933_ (.B1(_1979_),
    .Y(_2000_),
    .A1(_1978_),
    .A2(_1999_));
 sg13g2_a21oi_1 _5934_ (.A1(_1966_),
    .A2(_2000_),
    .Y(_2001_),
    .B1(_1964_));
 sg13g2_o21ai_1 _5935_ (.B1(_1953_),
    .Y(_2002_),
    .A1(_1952_),
    .A2(_2001_));
 sg13g2_nor2b_1 _5936_ (.A(_1942_),
    .B_N(_2002_),
    .Y(_2003_));
 sg13g2_a21oi_1 _5937_ (.A1(_1932_),
    .A2(_1941_),
    .Y(_2004_),
    .B1(_2003_));
 sg13g2_o21ai_1 _5938_ (.B1(_1938_),
    .Y(_2005_),
    .A1(_3197_),
    .A2(_1939_));
 sg13g2_o21ai_1 _5939_ (.B1(_1936_),
    .Y(_2006_),
    .A1(_1924_),
    .A2(_1934_));
 sg13g2_nand2_1 _5940_ (.Y(_2007_),
    .A(net1156),
    .B(net1068));
 sg13g2_nor2_1 _5941_ (.A(_1934_),
    .B(_2007_),
    .Y(_2008_));
 sg13g2_a22oi_1 _5942_ (.Y(_2009_),
    .B1(net1154),
    .B2(net1068),
    .A2(net1072),
    .A1(net1156));
 sg13g2_nor2_1 _5943_ (.A(_2008_),
    .B(_2009_),
    .Y(_2010_));
 sg13g2_xnor2_1 _5944_ (.Y(_2011_),
    .A(\vgademo.linelfsr[11] ),
    .B(_2010_));
 sg13g2_nand2b_1 _5945_ (.Y(_2012_),
    .B(_2006_),
    .A_N(_2011_));
 sg13g2_xor2_1 _5946_ (.B(_2011_),
    .A(_2006_),
    .X(_2013_));
 sg13g2_xnor2_1 _5947_ (.Y(_2014_),
    .A(_3196_),
    .B(_2013_));
 sg13g2_nand2b_1 _5948_ (.Y(_2015_),
    .B(_2005_),
    .A_N(_2014_));
 sg13g2_xor2_1 _5949_ (.B(_2014_),
    .A(_2005_),
    .X(_2016_));
 sg13g2_xor2_1 _5950_ (.B(_2016_),
    .A(_2004_),
    .X(_2017_));
 sg13g2_xnor2_1 _5951_ (.Y(_2018_),
    .A(\vgademo.linelfsr[3] ),
    .B(net1089));
 sg13g2_inv_1 _5952_ (.Y(_2019_),
    .A(_2018_));
 sg13g2_nand2b_1 _5953_ (.Y(_2020_),
    .B(_2019_),
    .A_N(_1993_));
 sg13g2_nor2_1 _5954_ (.A(_1992_),
    .B(_2020_),
    .Y(_2021_));
 sg13g2_xor2_1 _5955_ (.B(_1995_),
    .A(_1992_),
    .X(_2022_));
 sg13g2_a21oi_1 _5956_ (.A1(_2020_),
    .A2(_2022_),
    .Y(_2023_),
    .B1(_2021_));
 sg13g2_xor2_1 _5957_ (.B(_1994_),
    .A(_1993_),
    .X(_2024_));
 sg13g2_mux2_1 _5958_ (.A0(_1993_),
    .A1(_2024_),
    .S(_2018_),
    .X(_2025_));
 sg13g2_and2_1 _5959_ (.A(_3225_),
    .B(_2025_),
    .X(_2026_));
 sg13g2_xnor2_1 _5960_ (.Y(_2027_),
    .A(net1107),
    .B(_2025_));
 sg13g2_xnor2_1 _5961_ (.Y(_2028_),
    .A(_3226_),
    .B(_2018_));
 sg13g2_nand2_1 _5962_ (.Y(_2029_),
    .A(\vgademo.linelfsr[2] ),
    .B(_3224_));
 sg13g2_or2_1 _5963_ (.X(_2030_),
    .B(_2029_),
    .A(_2028_));
 sg13g2_o21ai_1 _5964_ (.B1(_2030_),
    .Y(_2031_),
    .A1(net1111),
    .A2(_2019_));
 sg13g2_a21oi_1 _5965_ (.A1(_2027_),
    .A2(_2031_),
    .Y(_2032_),
    .B1(_2026_));
 sg13g2_nand2b_1 _5966_ (.Y(_2033_),
    .B(_2023_),
    .A_N(_2032_));
 sg13g2_nand2b_1 _5967_ (.Y(_2034_),
    .B(_1979_),
    .A_N(_1978_));
 sg13g2_nor3_2 _5968_ (.A(_1998_),
    .B(_2033_),
    .C(_2034_),
    .Y(_2035_));
 sg13g2_nor2b_1 _5969_ (.A(_1952_),
    .B_N(_1953_),
    .Y(_2036_));
 sg13g2_xnor2_1 _5970_ (.Y(_2037_),
    .A(_1966_),
    .B(_2000_));
 sg13g2_xor2_1 _5971_ (.B(_2034_),
    .A(_1999_),
    .X(_2038_));
 sg13g2_xnor2_1 _5972_ (.Y(_2039_),
    .A(_1996_),
    .B(_1998_));
 sg13g2_nand3_1 _5973_ (.B(_2038_),
    .C(_2039_),
    .A(_2021_),
    .Y(_2040_));
 sg13g2_nor2_1 _5974_ (.A(_2037_),
    .B(_2040_),
    .Y(_2041_));
 sg13g2_xor2_1 _5975_ (.B(_2040_),
    .A(_2037_),
    .X(_2042_));
 sg13g2_nand3_1 _5976_ (.B(_2035_),
    .C(_2036_),
    .A(_1966_),
    .Y(_2043_));
 sg13g2_nor2_1 _5977_ (.A(_1942_),
    .B(_2043_),
    .Y(_2044_));
 sg13g2_and2_1 _5978_ (.A(_2017_),
    .B(_2044_),
    .X(_2045_));
 sg13g2_o21ai_1 _5979_ (.B1(_2015_),
    .Y(_2046_),
    .A1(_2004_),
    .A2(_2016_));
 sg13g2_o21ai_1 _5980_ (.B1(_2012_),
    .Y(_2047_),
    .A1(_3196_),
    .A2(_2013_));
 sg13g2_a21oi_1 _5981_ (.A1(\vgademo.linelfsr[11] ),
    .A2(_2010_),
    .Y(_2048_),
    .B1(_2008_));
 sg13g2_xnor2_1 _5982_ (.Y(_2049_),
    .A(\vgademo.linelfsr[12] ),
    .B(_2007_));
 sg13g2_nand2_1 _5983_ (.Y(_2050_),
    .A(net1067),
    .B(net1154));
 sg13g2_xor2_1 _5984_ (.B(_2050_),
    .A(net1066),
    .X(_2051_));
 sg13g2_xnor2_1 _5985_ (.Y(_2052_),
    .A(_2049_),
    .B(_2051_));
 sg13g2_xnor2_1 _5986_ (.Y(_2053_),
    .A(_2048_),
    .B(_2052_));
 sg13g2_xnor2_1 _5987_ (.Y(_2054_),
    .A(_2047_),
    .B(_2053_));
 sg13g2_xnor2_1 _5988_ (.Y(_2055_),
    .A(_2046_),
    .B(_2054_));
 sg13g2_xor2_1 _5989_ (.B(_2002_),
    .A(_1942_),
    .X(_2056_));
 sg13g2_xnor2_1 _5990_ (.Y(_2057_),
    .A(_2001_),
    .B(_2036_));
 sg13g2_inv_1 _5991_ (.Y(_2058_),
    .A(_2057_));
 sg13g2_and2_1 _5992_ (.A(_2041_),
    .B(_2057_),
    .X(_2059_));
 sg13g2_nor2b_1 _5993_ (.A(_2056_),
    .B_N(_2059_),
    .Y(_2060_));
 sg13g2_nand3_1 _5994_ (.B(_2055_),
    .C(_2060_),
    .A(_2017_),
    .Y(_2061_));
 sg13g2_a21o_1 _5995_ (.A2(_2060_),
    .A1(_2017_),
    .B1(_2055_),
    .X(_2062_));
 sg13g2_a21oi_1 _5996_ (.A1(_2061_),
    .A2(_2062_),
    .Y(_2063_),
    .B1(_2045_));
 sg13g2_nand2_1 _5997_ (.Y(_2064_),
    .A(\vgademo.h_count[10] ),
    .B(_2063_));
 sg13g2_or2_1 _5998_ (.X(_2065_),
    .B(_2060_),
    .A(_2044_));
 sg13g2_xor2_1 _5999_ (.B(_2065_),
    .A(_2017_),
    .X(_2066_));
 sg13g2_nor2_1 _6000_ (.A(_3195_),
    .B(_2066_),
    .Y(_2067_));
 sg13g2_a21oi_1 _6001_ (.A1(_1966_),
    .A2(_2035_),
    .Y(_2068_),
    .B1(_2041_));
 sg13g2_xnor2_1 _6002_ (.Y(_2069_),
    .A(_2058_),
    .B(_2068_));
 sg13g2_nor2_1 _6003_ (.A(\vgademo.h_count[7] ),
    .B(_2069_),
    .Y(_2070_));
 sg13g2_xnor2_1 _6004_ (.Y(_2071_),
    .A(_2035_),
    .B(_2042_));
 sg13g2_nand2b_1 _6005_ (.Y(_2072_),
    .B(_2033_),
    .A_N(_2021_));
 sg13g2_nand2_1 _6006_ (.Y(_2073_),
    .A(_2039_),
    .B(_2072_));
 sg13g2_xor2_1 _6007_ (.B(_2038_),
    .A(_0034_),
    .X(_2074_));
 sg13g2_xor2_1 _6008_ (.B(_2072_),
    .A(_2039_),
    .X(_2075_));
 sg13g2_nor2_1 _6009_ (.A(_0043_),
    .B(_2075_),
    .Y(_2076_));
 sg13g2_xor2_1 _6010_ (.B(_2032_),
    .A(_2023_),
    .X(_2077_));
 sg13g2_nor2_1 _6011_ (.A(net1093),
    .B(_2077_),
    .Y(_2078_));
 sg13g2_xor2_1 _6012_ (.B(_2031_),
    .A(_2027_),
    .X(_2079_));
 sg13g2_nand2_1 _6013_ (.Y(_2080_),
    .A(net1098),
    .B(_2029_));
 sg13g2_o21ai_1 _6014_ (.B1(_2080_),
    .Y(_2081_),
    .A1(\vgademo.linelfsr[2] ),
    .A2(_3224_));
 sg13g2_o21ai_1 _6015_ (.B1(_2081_),
    .Y(_2082_),
    .A1(net1096),
    .A2(_2028_));
 sg13g2_nand2_1 _6016_ (.Y(_2083_),
    .A(net1096),
    .B(_2028_));
 sg13g2_nand3_1 _6017_ (.B(_2082_),
    .C(_2083_),
    .A(_2030_),
    .Y(_2084_));
 sg13g2_nor2b_1 _6018_ (.A(_0032_),
    .B_N(_2084_),
    .Y(_2085_));
 sg13g2_a21oi_1 _6019_ (.A1(_0032_),
    .A2(_2084_),
    .Y(_2086_),
    .B1(net1095));
 sg13g2_nor2_1 _6020_ (.A(_2079_),
    .B(_2086_),
    .Y(_2087_));
 sg13g2_a21oi_1 _6021_ (.A1(_2079_),
    .A2(_2085_),
    .Y(_2088_),
    .B1(_2087_));
 sg13g2_nand2_1 _6022_ (.Y(_2089_),
    .A(net1093),
    .B(_2077_));
 sg13g2_xnor2_1 _6023_ (.Y(_2090_),
    .A(_2073_),
    .B(_2074_));
 sg13g2_a221oi_1 _6024_ (.B2(_2089_),
    .C1(_2078_),
    .B1(_2088_),
    .A1(_0043_),
    .Y(_2091_),
    .A2(_2075_));
 sg13g2_o21ai_1 _6025_ (.B1(_2090_),
    .Y(_2092_),
    .A1(_2076_),
    .A2(_2091_));
 sg13g2_a21oi_1 _6026_ (.A1(_2038_),
    .A2(_2073_),
    .Y(_2093_),
    .B1(_3192_));
 sg13g2_or2_1 _6027_ (.X(_2094_),
    .B(_2038_),
    .A(_3192_));
 sg13g2_o21ai_1 _6028_ (.B1(_2093_),
    .Y(_2095_),
    .A1(_2038_),
    .A2(_2073_));
 sg13g2_nand2_1 _6029_ (.Y(_2096_),
    .A(_2092_),
    .B(_2095_));
 sg13g2_xnor2_1 _6030_ (.Y(_2097_),
    .A(_0035_),
    .B(_2071_));
 sg13g2_a22oi_1 _6031_ (.Y(_2098_),
    .B1(_2096_),
    .B2(_2097_),
    .A2(_2071_),
    .A1(\vgademo.h_count[6] ));
 sg13g2_nor2_1 _6032_ (.A(_2070_),
    .B(_2098_),
    .Y(_2099_));
 sg13g2_xor2_1 _6033_ (.B(_2059_),
    .A(_2056_),
    .X(_2100_));
 sg13g2_a21oi_1 _6034_ (.A1(_2043_),
    .A2(_2100_),
    .Y(_2101_),
    .B1(_2044_));
 sg13g2_or2_1 _6035_ (.X(_2102_),
    .B(_2101_),
    .A(_0037_));
 sg13g2_a21oi_1 _6036_ (.A1(\vgademo.h_count[7] ),
    .A2(_2069_),
    .Y(_2103_),
    .B1(_2099_));
 sg13g2_nand2_1 _6037_ (.Y(_2104_),
    .A(_0037_),
    .B(_2101_));
 sg13g2_o21ai_1 _6038_ (.B1(_2104_),
    .Y(_2105_),
    .A1(_0038_),
    .A2(_2066_));
 sg13g2_a221oi_1 _6039_ (.B2(_2103_),
    .C1(_2105_),
    .B1(_2102_),
    .A1(_0038_),
    .Y(_2106_),
    .A2(_2066_));
 sg13g2_xnor2_1 _6040_ (.Y(_2107_),
    .A(net1092),
    .B(_2063_));
 sg13g2_o21ai_1 _6041_ (.B1(_2107_),
    .Y(_2108_),
    .A1(_2067_),
    .A2(_2106_));
 sg13g2_nand2_1 _6042_ (.Y(_2109_),
    .A(_2064_),
    .B(_2108_));
 sg13g2_nand2_1 _6043_ (.Y(_2110_),
    .A(_2045_),
    .B(_2062_));
 sg13g2_nand3_1 _6044_ (.B(_2109_),
    .C(_2110_),
    .A(_2061_),
    .Y(_2111_));
 sg13g2_xnor2_1 _6045_ (.Y(_2112_),
    .A(_0037_),
    .B(_2056_));
 sg13g2_nor2_1 _6046_ (.A(_0043_),
    .B(_2039_),
    .Y(_2113_));
 sg13g2_a22oi_1 _6047_ (.Y(_2114_),
    .B1(_2019_),
    .B2(_3188_),
    .A2(_3189_),
    .A1(\vgademo.linelfsr[2] ));
 sg13g2_a21oi_1 _6048_ (.A1(net1096),
    .A2(_2018_),
    .Y(_2115_),
    .B1(_2114_));
 sg13g2_nand2b_1 _6049_ (.Y(_2116_),
    .B(net1095),
    .A_N(_2024_));
 sg13g2_xnor2_1 _6050_ (.Y(_2117_),
    .A(_0032_),
    .B(_2024_));
 sg13g2_o21ai_1 _6051_ (.B1(_2116_),
    .Y(_2118_),
    .A1(_2115_),
    .A2(_2117_));
 sg13g2_o21ai_1 _6052_ (.B1(_2118_),
    .Y(_2119_),
    .A1(net1093),
    .A2(_2022_));
 sg13g2_nand2_1 _6053_ (.Y(_2120_),
    .A(net1093),
    .B(_2022_));
 sg13g2_a22oi_1 _6054_ (.Y(_2121_),
    .B1(_2119_),
    .B2(_2120_),
    .A2(_2039_),
    .A1(_0043_));
 sg13g2_o21ai_1 _6055_ (.B1(_2074_),
    .Y(_2122_),
    .A1(_2113_),
    .A2(_2121_));
 sg13g2_xor2_1 _6056_ (.B(_2037_),
    .A(_0035_),
    .X(_2123_));
 sg13g2_a21oi_1 _6057_ (.A1(_2094_),
    .A2(_2122_),
    .Y(_2124_),
    .B1(_2123_));
 sg13g2_a221oi_1 _6058_ (.B2(\vgademo.h_count[7] ),
    .C1(_2124_),
    .B1(_2058_),
    .A1(\vgademo.h_count[6] ),
    .Y(_2125_),
    .A2(_2037_));
 sg13g2_a21oi_1 _6059_ (.A1(_3194_),
    .A2(_2057_),
    .Y(_2126_),
    .B1(_2125_));
 sg13g2_a22oi_1 _6060_ (.Y(_2127_),
    .B1(_2112_),
    .B2(_2126_),
    .A2(_2056_),
    .A1(\vgademo.h_count[8] ));
 sg13g2_a21oi_1 _6061_ (.A1(_3195_),
    .A2(_2017_),
    .Y(_2128_),
    .B1(_2127_));
 sg13g2_nor2_1 _6062_ (.A(_3195_),
    .B(_2017_),
    .Y(_2129_));
 sg13g2_nor2_1 _6063_ (.A(_2128_),
    .B(_2129_),
    .Y(_2130_));
 sg13g2_o21ai_1 _6064_ (.B1(_2130_),
    .Y(_2131_),
    .A1(net1092),
    .A2(_2055_));
 sg13g2_nor2_1 _6065_ (.A(\vgademo.v_count[8] ),
    .B(net1073),
    .Y(_2132_));
 sg13g2_nor2_1 _6066_ (.A(net1059),
    .B(net1069),
    .Y(_2133_));
 sg13g2_xor2_1 _6067_ (.B(net1069),
    .A(net1059),
    .X(_2134_));
 sg13g2_nand2_1 _6068_ (.Y(_2135_),
    .A(net1060),
    .B(net1076));
 sg13g2_xor2_1 _6069_ (.B(net1073),
    .A(\vgademo.v_count[8] ),
    .X(_2136_));
 sg13g2_or2_1 _6070_ (.X(_2137_),
    .B(_2136_),
    .A(_2135_));
 sg13g2_nor2_1 _6071_ (.A(net1061),
    .B(net1078),
    .Y(_2138_));
 sg13g2_xnor2_1 _6072_ (.Y(_2139_),
    .A(net1060),
    .B(net1076));
 sg13g2_nor2_1 _6073_ (.A(_2138_),
    .B(_2139_),
    .Y(_2140_));
 sg13g2_nor2_1 _6074_ (.A(\vgademo.v_count[5] ),
    .B(net1081),
    .Y(_2141_));
 sg13g2_xor2_1 _6075_ (.B(net1078),
    .A(net1061),
    .X(_2142_));
 sg13g2_nor2_1 _6076_ (.A(_2141_),
    .B(_2142_),
    .Y(_2143_));
 sg13g2_or2_1 _6077_ (.X(_2144_),
    .B(net1084),
    .A(net1063));
 sg13g2_xnor2_1 _6078_ (.Y(_2145_),
    .A(\vgademo.v_count[5] ),
    .B(net1081));
 sg13g2_or2_1 _6079_ (.X(_2146_),
    .B(_2145_),
    .A(_2144_));
 sg13g2_nor2_1 _6080_ (.A(net1065),
    .B(net1091),
    .Y(_2147_));
 sg13g2_xnor2_1 _6081_ (.Y(_2148_),
    .A(net1063),
    .B(net1084));
 sg13g2_o21ai_1 _6082_ (.B1(_2148_),
    .Y(_2149_),
    .A1(net1064),
    .A2(net1087));
 sg13g2_a21oi_1 _6083_ (.A1(net1064),
    .A2(net1087),
    .Y(_2150_),
    .B1(_2148_));
 sg13g2_or2_1 _6084_ (.X(_2151_),
    .B(_2150_),
    .A(_2147_));
 sg13g2_nand2_1 _6085_ (.Y(_2152_),
    .A(_2146_),
    .B(_2149_));
 sg13g2_nor2b_1 _6086_ (.A(_2149_),
    .B_N(_2146_),
    .Y(_2153_));
 sg13g2_a21oi_1 _6087_ (.A1(_2144_),
    .A2(_2145_),
    .Y(_2154_),
    .B1(_2153_));
 sg13g2_o21ai_1 _6088_ (.B1(_2154_),
    .Y(_2155_),
    .A1(_2151_),
    .A2(_2152_));
 sg13g2_xnor2_1 _6089_ (.Y(_2156_),
    .A(_2141_),
    .B(_2142_));
 sg13g2_inv_1 _6090_ (.Y(_2157_),
    .A(_2156_));
 sg13g2_a21oi_1 _6091_ (.A1(_2155_),
    .A2(_2157_),
    .Y(_2158_),
    .B1(_2143_));
 sg13g2_xnor2_1 _6092_ (.Y(_2159_),
    .A(_2138_),
    .B(_2139_));
 sg13g2_nor2_1 _6093_ (.A(_2158_),
    .B(_2159_),
    .Y(_2160_));
 sg13g2_nor2_1 _6094_ (.A(_2140_),
    .B(_2160_),
    .Y(_2161_));
 sg13g2_xnor2_1 _6095_ (.Y(_2162_),
    .A(_2135_),
    .B(_2136_));
 sg13g2_o21ai_1 _6096_ (.B1(_2137_),
    .Y(_2163_),
    .A1(_2161_),
    .A2(_2162_));
 sg13g2_xnor2_1 _6097_ (.Y(_2164_),
    .A(_2132_),
    .B(_2134_));
 sg13g2_nand2b_1 _6098_ (.Y(_2165_),
    .B(_2163_),
    .A_N(_2164_));
 sg13g2_o21ai_1 _6099_ (.B1(_2165_),
    .Y(_2166_),
    .A1(_2132_),
    .A2(_2134_));
 sg13g2_xnor2_1 _6100_ (.Y(_2167_),
    .A(_3196_),
    .B(_2133_));
 sg13g2_inv_1 _6101_ (.Y(_2168_),
    .A(_2167_));
 sg13g2_nor2_1 _6102_ (.A(_0019_),
    .B(_2133_),
    .Y(_2169_));
 sg13g2_a21oi_2 _6103_ (.B1(_2169_),
    .Y(_2170_),
    .A2(_2168_),
    .A1(_2166_));
 sg13g2_nand2b_1 _6104_ (.Y(_2171_),
    .B(_2170_),
    .A_N(net1066));
 sg13g2_nor2b_1 _6105_ (.A(\vgademo.a_scrolly[13] ),
    .B_N(_2171_),
    .Y(_2172_));
 sg13g2_xnor2_1 _6106_ (.Y(_2173_),
    .A(_0065_),
    .B(_2172_));
 sg13g2_a22oi_1 _6107_ (.Y(_2174_),
    .B1(_2171_),
    .B2(\vgademo.a_scrolly[13] ),
    .A2(_2170_),
    .A1(_1048_));
 sg13g2_xnor2_1 _6108_ (.Y(_2175_),
    .A(_2158_),
    .B(_2159_));
 sg13g2_xor2_1 _6109_ (.B(_2170_),
    .A(_0066_),
    .X(_2176_));
 sg13g2_nand2_1 _6110_ (.Y(_2177_),
    .A(_2174_),
    .B(_2176_));
 sg13g2_xor2_1 _6111_ (.B(_2162_),
    .A(_2161_),
    .X(_2178_));
 sg13g2_inv_1 _6112_ (.Y(_2179_),
    .A(_2178_));
 sg13g2_xnor2_1 _6113_ (.Y(_2180_),
    .A(_2155_),
    .B(_2156_));
 sg13g2_xnor2_1 _6114_ (.Y(_2181_),
    .A(_2166_),
    .B(_2168_));
 sg13g2_xor2_1 _6115_ (.B(_2164_),
    .A(_2163_),
    .X(_2182_));
 sg13g2_and2_1 _6116_ (.A(_2174_),
    .B(_2182_),
    .X(_2183_));
 sg13g2_inv_1 _6117_ (.Y(_2184_),
    .A(_2183_));
 sg13g2_nand3b_1 _6118_ (.B(_2178_),
    .C(_2180_),
    .Y(_2185_),
    .A_N(_2175_));
 sg13g2_o21ai_1 _6119_ (.B1(_2174_),
    .Y(_2186_),
    .A1(_2181_),
    .A2(_2185_));
 sg13g2_nand4_1 _6120_ (.B(_2177_),
    .C(_2184_),
    .A(_2173_),
    .Y(_2187_),
    .D(_2186_));
 sg13g2_nand3_1 _6121_ (.B(_2131_),
    .C(_2187_),
    .A(_2111_),
    .Y(_2188_));
 sg13g2_a21oi_2 _6122_ (.B1(_2188_),
    .Y(_2189_),
    .A2(_2055_),
    .A1(net1092));
 sg13g2_nor3_1 _6123_ (.A(_1038_),
    .B(_1046_),
    .C(_1377_),
    .Y(_2190_));
 sg13g2_o21ai_1 _6124_ (.B1(net1075),
    .Y(_2191_),
    .A1(_1038_),
    .A2(_1377_));
 sg13g2_nand3_1 _6125_ (.B(_1200_),
    .C(_2191_),
    .A(_1050_),
    .Y(_2192_));
 sg13g2_nor2_2 _6126_ (.A(_2190_),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_inv_1 _6127_ (.Y(_2194_),
    .A(_2193_));
 sg13g2_and2_1 _6128_ (.A(_0077_),
    .B(_2193_),
    .X(_2195_));
 sg13g2_o21ai_1 _6129_ (.B1(net951),
    .Y(_2196_),
    .A1(_2189_),
    .A2(_2195_));
 sg13g2_nand2_2 _6130_ (.Y(_2197_),
    .A(_2173_),
    .B(_2194_));
 sg13g2_inv_1 _6131_ (.Y(_2198_),
    .A(_2197_));
 sg13g2_nand2_1 _6132_ (.Y(_2199_),
    .A(net951),
    .B(_2198_));
 sg13g2_nand3_1 _6133_ (.B(_2177_),
    .C(_2198_),
    .A(net951),
    .Y(_2200_));
 sg13g2_nand2_1 _6134_ (.Y(_2201_),
    .A(_2196_),
    .B(_2200_));
 sg13g2_a21oi_1 _6135_ (.A1(net896),
    .A2(_1916_),
    .Y(_2202_),
    .B1(_2201_));
 sg13g2_nand2_1 _6136_ (.Y(_2203_),
    .A(net939),
    .B(_1551_));
 sg13g2_xnor2_1 _6137_ (.Y(_2204_),
    .A(net939),
    .B(_1551_));
 sg13g2_nand2_2 _6138_ (.Y(_2205_),
    .A(_1371_),
    .B(net941));
 sg13g2_o21ai_1 _6139_ (.B1(_2203_),
    .Y(_2206_),
    .A1(_2204_),
    .A2(_2205_));
 sg13g2_xnor2_1 _6140_ (.Y(_2207_),
    .A(_1370_),
    .B(net928));
 sg13g2_xnor2_1 _6141_ (.Y(_2208_),
    .A(_2206_),
    .B(_2207_));
 sg13g2_inv_1 _6142_ (.Y(_2209_),
    .A(_2208_));
 sg13g2_nor4_2 _6143_ (.A(net903),
    .B(net900),
    .C(_1801_),
    .Y(_2210_),
    .D(_2209_));
 sg13g2_nand2_1 _6144_ (.Y(_2211_),
    .A(net935),
    .B(_1480_));
 sg13g2_and2_1 _6145_ (.A(_2205_),
    .B(_2211_),
    .X(_2212_));
 sg13g2_nor2b_1 _6146_ (.A(_2204_),
    .B_N(_2212_),
    .Y(_2213_));
 sg13g2_nor2_1 _6147_ (.A(net963),
    .B(_2210_),
    .Y(_2214_));
 sg13g2_a21oi_2 _6148_ (.B1(_1295_),
    .Y(_2215_),
    .A2(_2213_),
    .A1(_2210_));
 sg13g2_o21ai_1 _6149_ (.B1(_2215_),
    .Y(_2216_),
    .A1(_1802_),
    .A2(_2202_));
 sg13g2_nand2_2 _6150_ (.Y(_2217_),
    .A(_1318_),
    .B(_2216_));
 sg13g2_a21oi_1 _6151_ (.A1(_0074_),
    .A2(_2193_),
    .Y(_2218_),
    .B1(_2189_));
 sg13g2_a21oi_1 _6152_ (.A1(_2174_),
    .A2(_2181_),
    .Y(_2219_),
    .B1(_2197_));
 sg13g2_nand2b_1 _6153_ (.Y(_2220_),
    .B(_2218_),
    .A_N(_2219_));
 sg13g2_and3_1 _6154_ (.X(_2221_),
    .A(_1835_),
    .B(_1855_),
    .C(_1912_));
 sg13g2_or2_1 _6155_ (.X(_2222_),
    .B(_1905_),
    .A(_0054_));
 sg13g2_a21oi_2 _6156_ (.B1(_2221_),
    .Y(_2223_),
    .A2(_2222_),
    .A1(_1913_));
 sg13g2_nor2_1 _6157_ (.A(net951),
    .B(_2223_),
    .Y(_2224_));
 sg13g2_a22oi_1 _6158_ (.Y(_2225_),
    .B1(_2224_),
    .B2(net896),
    .A2(_2220_),
    .A1(net951));
 sg13g2_o21ai_1 _6159_ (.B1(_2215_),
    .Y(_2226_),
    .A1(_1802_),
    .A2(_2225_));
 sg13g2_xnor2_1 _6160_ (.Y(_2227_),
    .A(net1098),
    .B(net1089));
 sg13g2_xnor2_1 _6161_ (.Y(_2228_),
    .A(_3184_),
    .B(net1040));
 sg13g2_xnor2_1 _6162_ (.Y(_2229_),
    .A(\vgademo.bayer_j[0] ),
    .B(net1040));
 sg13g2_nand2b_1 _6163_ (.Y(_2230_),
    .B(_2228_),
    .A_N(_2226_));
 sg13g2_nand2b_1 _6164_ (.Y(_2231_),
    .B(_2230_),
    .A_N(_2217_));
 sg13g2_nand2_1 _6165_ (.Y(_2232_),
    .A(_2226_),
    .B(_2229_));
 sg13g2_nand2_1 _6166_ (.Y(_2233_),
    .A(_2217_),
    .B(_2232_));
 sg13g2_and2_1 _6167_ (.A(_2231_),
    .B(_2233_),
    .X(_2234_));
 sg13g2_nand2_1 _6168_ (.Y(_2235_),
    .A(net962),
    .B(_2212_));
 sg13g2_xor2_1 _6169_ (.B(_2205_),
    .A(_2204_),
    .X(_2236_));
 sg13g2_nor4_1 _6170_ (.A(net903),
    .B(net900),
    .C(_1801_),
    .D(_2236_),
    .Y(_2237_));
 sg13g2_or3_1 _6171_ (.A(net963),
    .B(_2210_),
    .C(_2237_),
    .X(_2238_));
 sg13g2_nor2_1 _6172_ (.A(_2209_),
    .B(_2236_),
    .Y(_2239_));
 sg13g2_nand2_1 _6173_ (.Y(_2240_),
    .A(net962),
    .B(_2239_));
 sg13g2_nand2_1 _6174_ (.Y(_2241_),
    .A(_2238_),
    .B(_2240_));
 sg13g2_nand3_1 _6175_ (.B(_2238_),
    .C(_2240_),
    .A(_2235_),
    .Y(_2242_));
 sg13g2_nor2b_2 _6176_ (.A(_1858_),
    .B_N(_1912_),
    .Y(_2243_));
 sg13g2_inv_1 _6177_ (.Y(_2244_),
    .A(_2243_));
 sg13g2_nand3_1 _6178_ (.B(_1829_),
    .C(_1830_),
    .A(_1826_),
    .Y(_2245_));
 sg13g2_nor2b_1 _6179_ (.A(_1831_),
    .B_N(_2245_),
    .Y(_2246_));
 sg13g2_nand2_1 _6180_ (.Y(_2247_),
    .A(_2243_),
    .B(_2246_));
 sg13g2_or2_1 _6181_ (.X(_2248_),
    .B(_1905_),
    .A(_0056_));
 sg13g2_a22oi_1 _6182_ (.Y(_2249_),
    .B1(_2248_),
    .B2(_1913_),
    .A2(_2246_),
    .A1(_2243_));
 sg13g2_nor4_1 _6183_ (.A(net902),
    .B(net899),
    .C(net947),
    .D(_1915_),
    .Y(_2250_));
 sg13g2_a221oi_1 _6184_ (.B2(_2249_),
    .C1(_2250_),
    .B1(net896),
    .A1(net957),
    .Y(_2251_),
    .A2(net960));
 sg13g2_and2_1 _6185_ (.A(_0055_),
    .B(_2193_),
    .X(_2252_));
 sg13g2_o21ai_1 _6186_ (.B1(net951),
    .Y(_2253_),
    .A1(_2189_),
    .A2(_2252_));
 sg13g2_inv_1 _6187_ (.Y(_2254_),
    .A(_2253_));
 sg13g2_o21ai_1 _6188_ (.B1(_2253_),
    .Y(_2255_),
    .A1(_2183_),
    .A2(_2199_));
 sg13g2_o21ai_1 _6189_ (.B1(net898),
    .Y(_2256_),
    .A1(_2251_),
    .A2(_2255_));
 sg13g2_nand2_1 _6190_ (.Y(_2257_),
    .A(_2242_),
    .B(_2256_));
 sg13g2_a21o_1 _6191_ (.A2(_2256_),
    .A1(_2242_),
    .B1(net1040),
    .X(_2258_));
 sg13g2_nand3_1 _6192_ (.B(_2242_),
    .C(_2256_),
    .A(net1040),
    .Y(_2259_));
 sg13g2_and3_1 _6193_ (.X(_2260_),
    .A(_2226_),
    .B(_2258_),
    .C(_2259_));
 sg13g2_nand3_1 _6194_ (.B(_2258_),
    .C(_2259_),
    .A(_2226_),
    .Y(_2261_));
 sg13g2_nand2_1 _6195_ (.Y(_2262_),
    .A(_2258_),
    .B(_2261_));
 sg13g2_and2_1 _6196_ (.A(_2230_),
    .B(_2232_),
    .X(_2263_));
 sg13g2_xnor2_1 _6197_ (.Y(_2264_),
    .A(_2217_),
    .B(_2263_));
 sg13g2_nor2_1 _6198_ (.A(_2262_),
    .B(_2264_),
    .Y(_2265_));
 sg13g2_xor2_1 _6199_ (.B(net1091),
    .A(net1097),
    .X(_2266_));
 sg13g2_o21ai_1 _6200_ (.B1(net905),
    .Y(_2267_),
    .A1(_0057_),
    .A2(_1905_));
 sg13g2_o21ai_1 _6201_ (.B1(_2267_),
    .Y(_2268_),
    .A1(_3247_),
    .A2(_2244_));
 sg13g2_a21o_1 _6202_ (.A2(_1828_),
    .A1(_1826_),
    .B1(_1827_),
    .X(_2269_));
 sg13g2_nand3_1 _6203_ (.B(_2243_),
    .C(_2269_),
    .A(_1829_),
    .Y(_2270_));
 sg13g2_o21ai_1 _6204_ (.B1(net905),
    .Y(_2271_),
    .A1(_0061_),
    .A2(_1905_));
 sg13g2_nand2_1 _6205_ (.Y(_2272_),
    .A(_2270_),
    .B(_2271_));
 sg13g2_inv_1 _6206_ (.Y(_2273_),
    .A(_2272_));
 sg13g2_nor4_1 _6207_ (.A(net904),
    .B(net901),
    .C(net948),
    .D(_2273_),
    .Y(_2274_));
 sg13g2_a221oi_1 _6208_ (.B2(_2268_),
    .C1(_2274_),
    .B1(net897),
    .A1(net958),
    .Y(_2275_),
    .A2(_1339_));
 sg13g2_nor2_1 _6209_ (.A(net955),
    .B(_2189_),
    .Y(_2276_));
 sg13g2_inv_1 _6210_ (.Y(_2277_),
    .A(_2276_));
 sg13g2_nand2_1 _6211_ (.Y(_2278_),
    .A(_1803_),
    .B(_2277_));
 sg13g2_nor2b_1 _6212_ (.A(_2180_),
    .B_N(_2174_),
    .Y(_2279_));
 sg13g2_nor2_1 _6213_ (.A(_2197_),
    .B(_2279_),
    .Y(_2280_));
 sg13g2_o21ai_1 _6214_ (.B1(net898),
    .Y(_2281_),
    .A1(_2277_),
    .A2(_2280_));
 sg13g2_o21ai_1 _6215_ (.B1(net961),
    .Y(_2282_),
    .A1(_2275_),
    .A2(_2281_));
 sg13g2_nand2_1 _6216_ (.Y(_2283_),
    .A(_2266_),
    .B(_2282_));
 sg13g2_nand2_1 _6217_ (.Y(_2284_),
    .A(_0063_),
    .B(_2193_));
 sg13g2_a21o_1 _6218_ (.A2(_2284_),
    .A1(_2276_),
    .B1(_1802_),
    .X(_2285_));
 sg13g2_a21o_1 _6219_ (.A2(_2175_),
    .A1(_2174_),
    .B1(_2197_),
    .X(_2286_));
 sg13g2_o21ai_1 _6220_ (.B1(_2285_),
    .Y(_2287_),
    .A1(_1802_),
    .A2(_2286_));
 sg13g2_nor2_1 _6221_ (.A(net1091),
    .B(\vgademo.plane_du[4] ),
    .Y(_2288_));
 sg13g2_or3_1 _6222_ (.A(_1827_),
    .B(_2244_),
    .C(_2288_),
    .X(_2289_));
 sg13g2_o21ai_1 _6223_ (.B1(net905),
    .Y(_2290_),
    .A1(_0058_),
    .A2(_1905_));
 sg13g2_nand2_1 _6224_ (.Y(_2291_),
    .A(_2289_),
    .B(_2290_));
 sg13g2_a21oi_1 _6225_ (.A1(net897),
    .A2(_2291_),
    .Y(_2292_),
    .B1(net951));
 sg13g2_o21ai_1 _6226_ (.B1(_2292_),
    .Y(_2293_),
    .A1(net896),
    .A2(_2249_));
 sg13g2_a21oi_1 _6227_ (.A1(_2287_),
    .A2(_2293_),
    .Y(_2294_),
    .B1(net963));
 sg13g2_nor2_1 _6228_ (.A(_2266_),
    .B(_2282_),
    .Y(_2295_));
 sg13g2_xor2_1 _6229_ (.B(_2282_),
    .A(_2266_),
    .X(_2296_));
 sg13g2_o21ai_1 _6230_ (.B1(_2283_),
    .Y(_2297_),
    .A1(_2294_),
    .A2(_2295_));
 sg13g2_nor4_1 _6231_ (.A(net902),
    .B(net899),
    .C(net947),
    .D(_2223_),
    .Y(_2298_));
 sg13g2_a221oi_1 _6232_ (.B2(_2272_),
    .C1(_2298_),
    .B1(net896),
    .A1(net957),
    .Y(_2299_),
    .A2(net960));
 sg13g2_o21ai_1 _6233_ (.B1(_2276_),
    .Y(_2300_),
    .A1(_3204_),
    .A2(_2194_));
 sg13g2_nand2_1 _6234_ (.Y(_2301_),
    .A(net898),
    .B(_2300_));
 sg13g2_a21oi_1 _6235_ (.A1(_2174_),
    .A2(_2179_),
    .Y(_2302_),
    .B1(_2197_));
 sg13g2_o21ai_1 _6236_ (.B1(net898),
    .Y(_2303_),
    .A1(_2300_),
    .A2(_2302_));
 sg13g2_nor2_1 _6237_ (.A(_2299_),
    .B(_2303_),
    .Y(_2304_));
 sg13g2_nor2b_1 _6238_ (.A(_2304_),
    .B_N(_2214_),
    .Y(_2305_));
 sg13g2_o21ai_1 _6239_ (.B1(_2214_),
    .Y(_2306_),
    .A1(_2299_),
    .A2(_2303_));
 sg13g2_xnor2_1 _6240_ (.Y(_2307_),
    .A(_3183_),
    .B(_2266_));
 sg13g2_and2_1 _6241_ (.A(_2306_),
    .B(_2307_),
    .X(_2308_));
 sg13g2_xor2_1 _6242_ (.B(_2307_),
    .A(_2306_),
    .X(_2309_));
 sg13g2_xnor2_1 _6243_ (.Y(_2310_),
    .A(_2257_),
    .B(_2309_));
 sg13g2_nor2b_1 _6244_ (.A(_2310_),
    .B_N(_2297_),
    .Y(_2311_));
 sg13g2_xor2_1 _6245_ (.B(net1091),
    .A(\vgademo.h_count[2] ),
    .X(_2312_));
 sg13g2_inv_1 _6246_ (.Y(_2313_),
    .A(_2312_));
 sg13g2_a21oi_1 _6247_ (.A1(_1318_),
    .A2(_2216_),
    .Y(_2314_),
    .B1(_2312_));
 sg13g2_a221oi_1 _6248_ (.B2(_2216_),
    .C1(net963),
    .B1(_2312_),
    .A1(_2287_),
    .Y(_2315_),
    .A2(_2293_));
 sg13g2_o21ai_1 _6249_ (.B1(_2305_),
    .Y(_2316_),
    .A1(_2314_),
    .A2(_2315_));
 sg13g2_xnor2_1 _6250_ (.Y(_2317_),
    .A(_2294_),
    .B(_2296_));
 sg13g2_nor3_1 _6251_ (.A(_2305_),
    .B(_2314_),
    .C(_2315_),
    .Y(_2318_));
 sg13g2_a21oi_1 _6252_ (.A1(_2257_),
    .A2(_2309_),
    .Y(_2319_),
    .B1(_2308_));
 sg13g2_a21oi_1 _6253_ (.A1(_2258_),
    .A2(_2259_),
    .Y(_2320_),
    .B1(_2226_));
 sg13g2_a21o_1 _6254_ (.A2(_2259_),
    .A1(_2258_),
    .B1(_2226_),
    .X(_2321_));
 sg13g2_a221oi_1 _6255_ (.B2(_2261_),
    .C1(_2308_),
    .B1(_2321_),
    .A1(_2257_),
    .Y(_2322_),
    .A2(_2309_));
 sg13g2_o21ai_1 _6256_ (.B1(_2319_),
    .Y(_2323_),
    .A1(_2260_),
    .A2(_2320_));
 sg13g2_nor3_1 _6257_ (.A(_2260_),
    .B(_2319_),
    .C(_2320_),
    .Y(_2324_));
 sg13g2_xor2_1 _6258_ (.B(_2310_),
    .A(_2297_),
    .X(_2325_));
 sg13g2_o21ai_1 _6259_ (.B1(_2316_),
    .Y(_2326_),
    .A1(_2317_),
    .A2(_2318_));
 sg13g2_or4_1 _6260_ (.A(_2322_),
    .B(_2324_),
    .C(_2325_),
    .D(_2326_),
    .X(_2327_));
 sg13g2_a221oi_1 _6261_ (.B2(_2323_),
    .C1(_2324_),
    .B1(_2311_),
    .A1(_2262_),
    .Y(_2328_),
    .A2(_2264_));
 sg13g2_a21oi_1 _6262_ (.A1(_2327_),
    .A2(_2328_),
    .Y(_2329_),
    .B1(_2265_));
 sg13g2_nand2_1 _6263_ (.Y(_2330_),
    .A(_2234_),
    .B(_2329_));
 sg13g2_nor4_1 _6264_ (.A(net1094),
    .B(net1095),
    .C(\vgademo.h_count[5] ),
    .D(\vgademo.h_count[4] ),
    .Y(_2331_));
 sg13g2_o21ai_1 _6265_ (.B1(_3319_),
    .Y(_2332_),
    .A1(_3283_),
    .A2(_2331_));
 sg13g2_nor2b_2 _6266_ (.A(net1092),
    .B_N(_2332_),
    .Y(_2333_));
 sg13g2_nor4_2 _6267_ (.A(net1064),
    .B(net1065),
    .C(_3316_),
    .Y(_2334_),
    .D(_0587_));
 sg13g2_nor4_2 _6268_ (.A(net518),
    .B(_3314_),
    .C(_2333_),
    .Y(_2335_),
    .D(_2334_));
 sg13g2_or4_2 _6269_ (.A(net1059),
    .B(_3314_),
    .C(_2333_),
    .D(_2334_),
    .X(_2336_));
 sg13g2_o21ai_1 _6270_ (.B1(_2335_),
    .Y(_2337_),
    .A1(_2234_),
    .A2(_2329_));
 sg13g2_nor2b_1 _6271_ (.A(_2337_),
    .B_N(_2330_),
    .Y(_0255_));
 sg13g2_a21oi_1 _6272_ (.A1(_2231_),
    .A2(_2330_),
    .Y(_0256_),
    .B1(_2336_));
 sg13g2_nand2_1 _6273_ (.Y(_2338_),
    .A(\vgademo.a_sin[6] ),
    .B(net996));
 sg13g2_xnor2_1 _6274_ (.Y(_0257_),
    .A(net250),
    .B(_2338_));
 sg13g2_nor2_1 _6275_ (.A(net313),
    .B(net996),
    .Y(_2339_));
 sg13g2_nand2b_1 _6276_ (.Y(_2340_),
    .B(\vgademo.a_sin[6] ),
    .A_N(net250));
 sg13g2_nor2b_1 _6277_ (.A(\vgademo.a_sin[7] ),
    .B_N(\vgademo.a_cos[1] ),
    .Y(_2341_));
 sg13g2_xnor2_1 _6278_ (.Y(_2342_),
    .A(\vgademo.a_sin[7] ),
    .B(net313));
 sg13g2_xnor2_1 _6279_ (.Y(_2343_),
    .A(_2340_),
    .B(_2342_));
 sg13g2_a21oi_1 _6280_ (.A1(net996),
    .A2(_2343_),
    .Y(_0258_),
    .B1(_2339_));
 sg13g2_nor2_1 _6281_ (.A(net302),
    .B(net997),
    .Y(_2344_));
 sg13g2_a21o_1 _6282_ (.A2(_2342_),
    .A1(_2340_),
    .B1(_2341_),
    .X(_2345_));
 sg13g2_nor2b_1 _6283_ (.A(\vgademo.a_sin[8] ),
    .B_N(\vgademo.a_cos[2] ),
    .Y(_2346_));
 sg13g2_xnor2_1 _6284_ (.Y(_2347_),
    .A(\vgademo.a_sin[8] ),
    .B(net302));
 sg13g2_xnor2_1 _6285_ (.Y(_2348_),
    .A(_2345_),
    .B(_2347_));
 sg13g2_a21oi_1 _6286_ (.A1(net997),
    .A2(_2348_),
    .Y(_0259_),
    .B1(_2344_));
 sg13g2_nor2_1 _6287_ (.A(net394),
    .B(net996),
    .Y(_2349_));
 sg13g2_a21o_1 _6288_ (.A2(_2347_),
    .A1(_2345_),
    .B1(_2346_),
    .X(_2350_));
 sg13g2_nor2b_1 _6289_ (.A(\vgademo.a_sin[9] ),
    .B_N(\vgademo.a_cos[3] ),
    .Y(_2351_));
 sg13g2_xnor2_1 _6290_ (.Y(_2352_),
    .A(\vgademo.a_cos[3] ),
    .B(\vgademo.a_sin[9] ));
 sg13g2_xnor2_1 _6291_ (.Y(_2353_),
    .A(_2350_),
    .B(_2352_));
 sg13g2_a21oi_1 _6292_ (.A1(net996),
    .A2(_2353_),
    .Y(_0260_),
    .B1(_2349_));
 sg13g2_nand2_1 _6293_ (.Y(_2354_),
    .A(net444),
    .B(net1019));
 sg13g2_a21oi_1 _6294_ (.A1(_2350_),
    .A2(_2352_),
    .Y(_2355_),
    .B1(_2351_));
 sg13g2_nand2b_1 _6295_ (.Y(_2356_),
    .B(\vgademo.a_cos[4] ),
    .A_N(\vgademo.a_sin[10] ));
 sg13g2_xor2_1 _6296_ (.B(\vgademo.a_sin[10] ),
    .A(\vgademo.a_cos[4] ),
    .X(_2357_));
 sg13g2_xnor2_1 _6297_ (.Y(_2358_),
    .A(_2355_),
    .B(_2357_));
 sg13g2_o21ai_1 _6298_ (.B1(_2354_),
    .Y(_0261_),
    .A1(net1019),
    .A2(_2358_));
 sg13g2_nor2_1 _6299_ (.A(net443),
    .B(net1022),
    .Y(_2359_));
 sg13g2_o21ai_1 _6300_ (.B1(_2356_),
    .Y(_2360_),
    .A1(_2355_),
    .A2(_2357_));
 sg13g2_nor2b_1 _6301_ (.A(\vgademo.a_sin[11] ),
    .B_N(\vgademo.a_cos[5] ),
    .Y(_2361_));
 sg13g2_nand2b_1 _6302_ (.Y(_2362_),
    .B(\vgademo.a_sin[11] ),
    .A_N(\vgademo.a_cos[5] ));
 sg13g2_nor2b_1 _6303_ (.A(_2361_),
    .B_N(_2362_),
    .Y(_2363_));
 sg13g2_xnor2_1 _6304_ (.Y(_2364_),
    .A(_2360_),
    .B(_2363_));
 sg13g2_a21oi_1 _6305_ (.A1(net997),
    .A2(_2364_),
    .Y(_0262_),
    .B1(_2359_));
 sg13g2_nor2_1 _6306_ (.A(_3231_),
    .B(\vgademo.a_sin[12] ),
    .Y(_2365_));
 sg13g2_xor2_1 _6307_ (.B(\vgademo.a_sin[12] ),
    .A(\vgademo.a_cos[6] ),
    .X(_2366_));
 sg13g2_a21oi_1 _6308_ (.A1(_2360_),
    .A2(_2362_),
    .Y(_2367_),
    .B1(_2361_));
 sg13g2_nor2_1 _6309_ (.A(_2366_),
    .B(_2367_),
    .Y(_2368_));
 sg13g2_xor2_1 _6310_ (.B(_2367_),
    .A(_2366_),
    .X(_2369_));
 sg13g2_nand2_1 _6311_ (.Y(_2370_),
    .A(net1022),
    .B(_2369_));
 sg13g2_o21ai_1 _6312_ (.B1(_2370_),
    .Y(_0263_),
    .A1(_3231_),
    .A2(net997));
 sg13g2_xnor2_1 _6313_ (.Y(_2371_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.a_sin[13] ));
 sg13g2_o21ai_1 _6314_ (.B1(_2371_),
    .Y(_2372_),
    .A1(_2365_),
    .A2(_2368_));
 sg13g2_or3_1 _6315_ (.A(_2365_),
    .B(_2368_),
    .C(_2371_),
    .X(_2373_));
 sg13g2_and2_1 _6316_ (.A(_2372_),
    .B(_2373_),
    .X(_2374_));
 sg13g2_nand2_1 _6317_ (.Y(_2375_),
    .A(net997),
    .B(_2374_));
 sg13g2_o21ai_1 _6318_ (.B1(_2375_),
    .Y(_0264_),
    .A1(_3233_),
    .A2(net997));
 sg13g2_o21ai_1 _6319_ (.B1(_2372_),
    .Y(_2376_),
    .A1(_3233_),
    .A2(\vgademo.a_sin[13] ));
 sg13g2_xnor2_1 _6320_ (.Y(_2377_),
    .A(\vgademo.a_cos[8] ),
    .B(net1058));
 sg13g2_and2_1 _6321_ (.A(_2376_),
    .B(_2377_),
    .X(_2378_));
 sg13g2_xor2_1 _6322_ (.B(_2377_),
    .A(_2376_),
    .X(_2379_));
 sg13g2_mux2_1 _6323_ (.A0(net573),
    .A1(_2379_),
    .S(net996),
    .X(_0265_));
 sg13g2_nor2_1 _6324_ (.A(net522),
    .B(net1021),
    .Y(_2380_));
 sg13g2_xnor2_1 _6325_ (.Y(_2381_),
    .A(\vgademo.a_cos[9] ),
    .B(net1058));
 sg13g2_a21oi_1 _6326_ (.A1(\vgademo.a_cos[8] ),
    .A2(_3245_),
    .Y(_2382_),
    .B1(_2378_));
 sg13g2_xor2_1 _6327_ (.B(_2382_),
    .A(_2381_),
    .X(_2383_));
 sg13g2_a21oi_1 _6328_ (.A1(net1021),
    .A2(_2383_),
    .Y(_0266_),
    .B1(_2380_));
 sg13g2_xnor2_1 _6329_ (.Y(_2384_),
    .A(\vgademo.a_cos[10] ),
    .B(net1057));
 sg13g2_o21ai_1 _6330_ (.B1(_3245_),
    .Y(_2385_),
    .A1(\vgademo.a_cos[8] ),
    .A2(\vgademo.a_cos[9] ));
 sg13g2_inv_1 _6331_ (.Y(_2386_),
    .A(_2385_));
 sg13g2_a21oi_1 _6332_ (.A1(_2378_),
    .A2(_2381_),
    .Y(_2387_),
    .B1(_2386_));
 sg13g2_nand2b_1 _6333_ (.Y(_2388_),
    .B(_2384_),
    .A_N(_2387_));
 sg13g2_xnor2_1 _6334_ (.Y(_2389_),
    .A(_2384_),
    .B(_2387_));
 sg13g2_nand2_1 _6335_ (.Y(_2390_),
    .A(net998),
    .B(_2389_));
 sg13g2_o21ai_1 _6336_ (.B1(_2390_),
    .Y(_0267_),
    .A1(_3236_),
    .A2(net998));
 sg13g2_nor2_1 _6337_ (.A(net439),
    .B(net1023),
    .Y(_2391_));
 sg13g2_xnor2_1 _6338_ (.Y(_2392_),
    .A(\vgademo.a_cos[11] ),
    .B(net1057));
 sg13g2_o21ai_1 _6339_ (.B1(_2388_),
    .Y(_2393_),
    .A1(_3236_),
    .A2(net1057));
 sg13g2_xnor2_1 _6340_ (.Y(_2394_),
    .A(_2392_),
    .B(_2393_));
 sg13g2_a21oi_1 _6341_ (.A1(net1023),
    .A2(_2394_),
    .Y(_0268_),
    .B1(_2391_));
 sg13g2_nor2_1 _6342_ (.A(net437),
    .B(net1023),
    .Y(_2395_));
 sg13g2_nand4_1 _6343_ (.B(_2381_),
    .C(_2384_),
    .A(_2378_),
    .Y(_2396_),
    .D(_2392_));
 sg13g2_o21ai_1 _6344_ (.B1(_3245_),
    .Y(_2397_),
    .A1(\vgademo.a_cos[10] ),
    .A2(\vgademo.a_cos[11] ));
 sg13g2_nand3_1 _6345_ (.B(_2396_),
    .C(_2397_),
    .A(_2385_),
    .Y(_2398_));
 sg13g2_nor2b_1 _6346_ (.A(net1057),
    .B_N(\vgademo.a_cos[12] ),
    .Y(_2399_));
 sg13g2_xnor2_1 _6347_ (.Y(_2400_),
    .A(\vgademo.a_cos[12] ),
    .B(net1057));
 sg13g2_xnor2_1 _6348_ (.Y(_2401_),
    .A(_2398_),
    .B(_2400_));
 sg13g2_a21oi_1 _6349_ (.A1(net1023),
    .A2(_2401_),
    .Y(_0269_),
    .B1(_2395_));
 sg13g2_nor2_1 _6350_ (.A(net236),
    .B(net1023),
    .Y(_2402_));
 sg13g2_a21oi_1 _6351_ (.A1(_2398_),
    .A2(_2400_),
    .Y(_2403_),
    .B1(_2399_));
 sg13g2_nand2_1 _6352_ (.Y(_2404_),
    .A(\vgademo.a_cos[13] ),
    .B(_3245_));
 sg13g2_nor2_1 _6353_ (.A(\vgademo.a_cos[13] ),
    .B(_3245_),
    .Y(_2405_));
 sg13g2_xnor2_1 _6354_ (.Y(_2406_),
    .A(\vgademo.a_cos[13] ),
    .B(net1057));
 sg13g2_xnor2_1 _6355_ (.Y(_2407_),
    .A(_2403_),
    .B(_2406_));
 sg13g2_a21oi_1 _6356_ (.A1(net1023),
    .A2(_2407_),
    .Y(_0270_),
    .B1(_2402_));
 sg13g2_nor2_1 _6357_ (.A(net422),
    .B(net998),
    .Y(_2408_));
 sg13g2_o21ai_1 _6358_ (.B1(_2404_),
    .Y(_2409_),
    .A1(_2403_),
    .A2(_2405_));
 sg13g2_xnor2_1 _6359_ (.Y(_2410_),
    .A(\vgademo.a_cos[14] ),
    .B(net1057));
 sg13g2_xnor2_1 _6360_ (.Y(_2411_),
    .A(_2409_),
    .B(_2410_));
 sg13g2_inv_1 _6361_ (.Y(_2412_),
    .A(_2411_));
 sg13g2_a21oi_1 _6362_ (.A1(net998),
    .A2(net927),
    .Y(_0271_),
    .B1(_2408_));
 sg13g2_xnor2_1 _6363_ (.Y(_0272_),
    .A(net237),
    .B(_2370_));
 sg13g2_nor2_1 _6364_ (.A(net347),
    .B(net1022),
    .Y(_2413_));
 sg13g2_nand2_1 _6365_ (.Y(_2414_),
    .A(net237),
    .B(_2369_));
 sg13g2_xnor2_1 _6366_ (.Y(_2415_),
    .A(\vgademo.a_sin[1] ),
    .B(_2374_));
 sg13g2_nor2_1 _6367_ (.A(_2414_),
    .B(_2415_),
    .Y(_2416_));
 sg13g2_xnor2_1 _6368_ (.Y(_2417_),
    .A(_2414_),
    .B(_2415_));
 sg13g2_a21oi_1 _6369_ (.A1(net1022),
    .A2(_2417_),
    .Y(_0273_),
    .B1(_2413_));
 sg13g2_nor2_1 _6370_ (.A(net349),
    .B(net1021),
    .Y(_2418_));
 sg13g2_a21oi_2 _6371_ (.B1(_2416_),
    .Y(_2419_),
    .A2(_2374_),
    .A1(net347));
 sg13g2_and2_1 _6372_ (.A(\vgademo.a_sin[2] ),
    .B(_2379_),
    .X(_2420_));
 sg13g2_xnor2_1 _6373_ (.Y(_2421_),
    .A(net349),
    .B(_2379_));
 sg13g2_nor2_1 _6374_ (.A(_2419_),
    .B(_2421_),
    .Y(_2422_));
 sg13g2_xnor2_1 _6375_ (.Y(_2423_),
    .A(_2419_),
    .B(_2421_));
 sg13g2_a21oi_1 _6376_ (.A1(net1021),
    .A2(_2423_),
    .Y(_0274_),
    .B1(_2418_));
 sg13g2_or2_1 _6377_ (.X(_2424_),
    .B(_2383_),
    .A(_3240_));
 sg13g2_xnor2_1 _6378_ (.Y(_2425_),
    .A(\vgademo.a_sin[3] ),
    .B(_2383_));
 sg13g2_o21ai_1 _6379_ (.B1(_2425_),
    .Y(_2426_),
    .A1(_2420_),
    .A2(_2422_));
 sg13g2_or3_1 _6380_ (.A(_2420_),
    .B(_2422_),
    .C(_2425_),
    .X(_2427_));
 sg13g2_a21oi_1 _6381_ (.A1(_2426_),
    .A2(_2427_),
    .Y(_2428_),
    .B1(net1020));
 sg13g2_a21oi_1 _6382_ (.A1(_3240_),
    .A2(net1020),
    .Y(_0275_),
    .B1(_2428_));
 sg13g2_and2_1 _6383_ (.A(\vgademo.a_sin[4] ),
    .B(_2389_),
    .X(_2429_));
 sg13g2_xnor2_1 _6384_ (.Y(_2430_),
    .A(\vgademo.a_sin[4] ),
    .B(_2389_));
 sg13g2_a21oi_2 _6385_ (.B1(_2430_),
    .Y(_2431_),
    .A2(_2426_),
    .A1(_2424_));
 sg13g2_nand3_1 _6386_ (.B(_2426_),
    .C(_2430_),
    .A(_2424_),
    .Y(_2432_));
 sg13g2_o21ai_1 _6387_ (.B1(net355),
    .Y(_2433_),
    .A1(net1034),
    .A2(_0590_));
 sg13g2_nand2_1 _6388_ (.Y(_2434_),
    .A(net998),
    .B(_2432_));
 sg13g2_o21ai_1 _6389_ (.B1(_2433_),
    .Y(_0276_),
    .A1(_2431_),
    .A2(_2434_));
 sg13g2_nand2b_1 _6390_ (.Y(_2435_),
    .B(net311),
    .A_N(_2394_));
 sg13g2_xnor2_1 _6391_ (.Y(_2436_),
    .A(\vgademo.a_sin[5] ),
    .B(_2394_));
 sg13g2_o21ai_1 _6392_ (.B1(_2436_),
    .Y(_2437_),
    .A1(_2429_),
    .A2(_2431_));
 sg13g2_or3_1 _6393_ (.A(_2429_),
    .B(_2431_),
    .C(_2436_),
    .X(_2438_));
 sg13g2_a21oi_1 _6394_ (.A1(_2437_),
    .A2(_2438_),
    .Y(_2439_),
    .B1(net1019));
 sg13g2_a21oi_1 _6395_ (.A1(_3241_),
    .A2(net1019),
    .Y(_0277_),
    .B1(_2439_));
 sg13g2_nor2_1 _6396_ (.A(_3171_),
    .B(_2401_),
    .Y(_2440_));
 sg13g2_xnor2_1 _6397_ (.Y(_2441_),
    .A(_3171_),
    .B(_2401_));
 sg13g2_a21oi_1 _6398_ (.A1(_2435_),
    .A2(_2437_),
    .Y(_2442_),
    .B1(_2441_));
 sg13g2_nand3_1 _6399_ (.B(_2437_),
    .C(_2441_),
    .A(_2435_),
    .Y(_2443_));
 sg13g2_nand3b_1 _6400_ (.B(_2443_),
    .C(net998),
    .Y(_2444_),
    .A_N(_2442_));
 sg13g2_o21ai_1 _6401_ (.B1(_2444_),
    .Y(_0278_),
    .A1(_3171_),
    .A2(net998));
 sg13g2_nand2_1 _6402_ (.Y(_2445_),
    .A(\vgademo.a_sin[7] ),
    .B(_2407_));
 sg13g2_xnor2_1 _6403_ (.Y(_2446_),
    .A(_3242_),
    .B(_2407_));
 sg13g2_o21ai_1 _6404_ (.B1(_2446_),
    .Y(_2447_),
    .A1(_2440_),
    .A2(_2442_));
 sg13g2_or3_1 _6405_ (.A(_2440_),
    .B(_2442_),
    .C(_2446_),
    .X(_2448_));
 sg13g2_a21oi_1 _6406_ (.A1(_2447_),
    .A2(_2448_),
    .Y(_2449_),
    .B1(net1019));
 sg13g2_a21oi_1 _6407_ (.A1(_3242_),
    .A2(net1019),
    .Y(_0279_),
    .B1(_2449_));
 sg13g2_xor2_1 _6408_ (.B(net927),
    .A(\vgademo.a_sin[8] ),
    .X(_2450_));
 sg13g2_a21oi_2 _6409_ (.B1(_2450_),
    .Y(_2451_),
    .A2(_2447_),
    .A1(_2445_));
 sg13g2_nand3_1 _6410_ (.B(_2447_),
    .C(_2450_),
    .A(_2445_),
    .Y(_2452_));
 sg13g2_o21ai_1 _6411_ (.B1(net574),
    .Y(_2453_),
    .A1(net1034),
    .A2(_0590_));
 sg13g2_nand2_1 _6412_ (.Y(_2454_),
    .A(net998),
    .B(_2452_));
 sg13g2_o21ai_1 _6413_ (.B1(_2453_),
    .Y(_0280_),
    .A1(_2451_),
    .A2(_2454_));
 sg13g2_nor2_1 _6414_ (.A(net474),
    .B(net1021),
    .Y(_2455_));
 sg13g2_a21oi_1 _6415_ (.A1(\vgademo.a_sin[8] ),
    .A2(_2412_),
    .Y(_2456_),
    .B1(_2451_));
 sg13g2_xnor2_1 _6416_ (.Y(_2457_),
    .A(\vgademo.a_sin[9] ),
    .B(_2411_));
 sg13g2_xor2_1 _6417_ (.B(_2457_),
    .A(_2456_),
    .X(_2458_));
 sg13g2_a21oi_1 _6418_ (.A1(net996),
    .A2(_2458_),
    .Y(_0281_),
    .B1(_2455_));
 sg13g2_nor2_1 _6419_ (.A(net479),
    .B(net1021),
    .Y(_2459_));
 sg13g2_o21ai_1 _6420_ (.B1(_2412_),
    .Y(_2460_),
    .A1(\vgademo.a_sin[8] ),
    .A2(\vgademo.a_sin[9] ));
 sg13g2_and2_1 _6421_ (.A(_2451_),
    .B(_2457_),
    .X(_2461_));
 sg13g2_nor2b_1 _6422_ (.A(_2461_),
    .B_N(_2460_),
    .Y(_2462_));
 sg13g2_nand2_1 _6423_ (.Y(_2463_),
    .A(\vgademo.a_sin[10] ),
    .B(_2412_));
 sg13g2_xor2_1 _6424_ (.B(net927),
    .A(\vgademo.a_sin[10] ),
    .X(_2464_));
 sg13g2_xnor2_1 _6425_ (.Y(_2465_),
    .A(_2462_),
    .B(_2464_));
 sg13g2_a21oi_1 _6426_ (.A1(net1021),
    .A2(_2465_),
    .Y(_0282_),
    .B1(_2459_));
 sg13g2_nand2_1 _6427_ (.Y(_2466_),
    .A(net451),
    .B(net1019));
 sg13g2_o21ai_1 _6428_ (.B1(_2463_),
    .Y(_2467_),
    .A1(_2462_),
    .A2(_2464_));
 sg13g2_xnor2_1 _6429_ (.Y(_2468_),
    .A(\vgademo.a_sin[11] ),
    .B(net927));
 sg13g2_xnor2_1 _6430_ (.Y(_2469_),
    .A(_2467_),
    .B(_2468_));
 sg13g2_o21ai_1 _6431_ (.B1(_2466_),
    .Y(_0283_),
    .A1(net1019),
    .A2(_2469_));
 sg13g2_a21oi_1 _6432_ (.A1(_3243_),
    .A2(net927),
    .Y(_2470_),
    .B1(_2464_));
 sg13g2_o21ai_1 _6433_ (.B1(_2412_),
    .Y(_2471_),
    .A1(\vgademo.a_sin[10] ),
    .A2(\vgademo.a_sin[11] ));
 sg13g2_nand2_1 _6434_ (.Y(_2472_),
    .A(_2460_),
    .B(_2471_));
 sg13g2_a21oi_2 _6435_ (.B1(_2472_),
    .Y(_2473_),
    .A2(_2470_),
    .A1(_2461_));
 sg13g2_xnor2_1 _6436_ (.Y(_2474_),
    .A(\vgademo.a_sin[12] ),
    .B(net927));
 sg13g2_nand2b_1 _6437_ (.Y(_2475_),
    .B(_2474_),
    .A_N(_2473_));
 sg13g2_xnor2_1 _6438_ (.Y(_2476_),
    .A(_2473_),
    .B(_2474_));
 sg13g2_nand2_1 _6439_ (.Y(_2477_),
    .A(net1021),
    .B(_2476_));
 sg13g2_o21ai_1 _6440_ (.B1(_2477_),
    .Y(_0284_),
    .A1(_3244_),
    .A2(net996));
 sg13g2_nand2_1 _6441_ (.Y(_2478_),
    .A(net927),
    .B(_2475_));
 sg13g2_a21oi_1 _6442_ (.A1(_3244_),
    .A2(_2473_),
    .Y(_2479_),
    .B1(net927));
 sg13g2_nor2_1 _6443_ (.A(net1020),
    .B(_2479_),
    .Y(_2480_));
 sg13g2_nand2_1 _6444_ (.Y(_2481_),
    .A(_2478_),
    .B(_2480_));
 sg13g2_xnor2_1 _6445_ (.Y(_0285_),
    .A(net501),
    .B(_2481_));
 sg13g2_nor2_1 _6446_ (.A(net501),
    .B(_2412_),
    .Y(_2482_));
 sg13g2_a21oi_1 _6447_ (.A1(net501),
    .A2(_2475_),
    .Y(_2483_),
    .B1(_2482_));
 sg13g2_nand2_1 _6448_ (.Y(_2484_),
    .A(_2480_),
    .B(_2483_));
 sg13g2_xnor2_1 _6449_ (.Y(_0286_),
    .A(net1058),
    .B(_2484_));
 sg13g2_and4_1 _6450_ (.A(\vgademo.h_count[10] ),
    .B(net1181),
    .C(_3319_),
    .D(_0579_),
    .X(_2485_));
 sg13g2_nand2_1 _6451_ (.Y(_2486_),
    .A(_0498_),
    .B(net988));
 sg13g2_o21ai_1 _6452_ (.B1(_2486_),
    .Y(_0287_),
    .A1(_3282_),
    .A2(net992));
 sg13g2_mux2_1 _6453_ (.A0(net353),
    .A1(_0513_),
    .S(net988),
    .X(_0288_));
 sg13g2_mux2_1 _6454_ (.A0(net332),
    .A1(_0527_),
    .S(net992),
    .X(_0289_));
 sg13g2_nand2_1 _6455_ (.Y(_2487_),
    .A(_0543_),
    .B(net988));
 sg13g2_o21ai_1 _6456_ (.B1(_2487_),
    .Y(_0290_),
    .A1(_3281_),
    .A2(net988));
 sg13g2_mux2_1 _6457_ (.A0(net425),
    .A1(_0557_),
    .S(net988),
    .X(_0291_));
 sg13g2_nand2_1 _6458_ (.Y(_2488_),
    .A(_0563_),
    .B(net988));
 sg13g2_o21ai_1 _6459_ (.B1(_2488_),
    .Y(_0292_),
    .A1(_3280_),
    .A2(net988));
 sg13g2_mux2_1 _6460_ (.A0(net447),
    .A1(_0562_),
    .S(net988),
    .X(_0293_));
 sg13g2_o21ai_1 _6461_ (.B1(net325),
    .Y(_2489_),
    .A1(_3227_),
    .A2(net1026));
 sg13g2_nor2_2 _6462_ (.A(net325),
    .B(_3227_),
    .Y(_2490_));
 sg13g2_nor2_1 _6463_ (.A(net1008),
    .B(net1025),
    .Y(_2491_));
 sg13g2_nand2_2 _6464_ (.Y(_2492_),
    .A(net1006),
    .B(_0582_));
 sg13g2_a22oi_1 _6465_ (.Y(_2493_),
    .B1(_2490_),
    .B2(_2491_),
    .A2(net985),
    .A1(\vgademo.a_cos[3] ));
 sg13g2_o21ai_1 _6466_ (.B1(_2493_),
    .Y(_0294_),
    .A1(net985),
    .A2(_2489_));
 sg13g2_xnor2_1 _6467_ (.Y(_2494_),
    .A(net441),
    .B(\vgademo.b_sin[8] ));
 sg13g2_nor2b_1 _6468_ (.A(_2490_),
    .B_N(_2494_),
    .Y(_2495_));
 sg13g2_xor2_1 _6469_ (.B(_2494_),
    .A(_2490_),
    .X(_2496_));
 sg13g2_nand2b_1 _6470_ (.Y(_2497_),
    .B(net985),
    .A_N(\vgademo.a_cos[4] ));
 sg13g2_o21ai_1 _6471_ (.B1(_2497_),
    .Y(_2498_),
    .A1(net441),
    .A2(_0582_));
 sg13g2_a21oi_1 _6472_ (.A1(net984),
    .A2(_2496_),
    .Y(_0295_),
    .B1(net442));
 sg13g2_nand2b_1 _6473_ (.Y(_2499_),
    .B(net985),
    .A_N(net443));
 sg13g2_a21oi_1 _6474_ (.A1(\vgademo.b_cos[1] ),
    .A2(_3228_),
    .Y(_2500_),
    .B1(_2495_));
 sg13g2_xnor2_1 _6475_ (.Y(_2501_),
    .A(net449),
    .B(\vgademo.b_sin[9] ));
 sg13g2_nor2b_1 _6476_ (.A(_2500_),
    .B_N(_2501_),
    .Y(_2502_));
 sg13g2_xor2_1 _6477_ (.B(_2501_),
    .A(_2500_),
    .X(_2503_));
 sg13g2_o21ai_1 _6478_ (.B1(_2499_),
    .Y(_2504_),
    .A1(net449),
    .A2(_0582_));
 sg13g2_a21oi_1 _6479_ (.A1(net984),
    .A2(_2503_),
    .Y(_0296_),
    .B1(_2504_));
 sg13g2_a21oi_1 _6480_ (.A1(\vgademo.b_cos[2] ),
    .A2(_3229_),
    .Y(_2505_),
    .B1(_2502_));
 sg13g2_xnor2_1 _6481_ (.Y(_2506_),
    .A(\vgademo.b_cos[3] ),
    .B(\vgademo.b_sin[10] ));
 sg13g2_nor2b_1 _6482_ (.A(_2505_),
    .B_N(_2506_),
    .Y(_2507_));
 sg13g2_xor2_1 _6483_ (.B(_2506_),
    .A(_2505_),
    .X(_2508_));
 sg13g2_nor2_1 _6484_ (.A(net357),
    .B(net1027),
    .Y(_2509_));
 sg13g2_a221oi_1 _6485_ (.B2(_2508_),
    .C1(_2509_),
    .B1(net984),
    .A1(_3231_),
    .Y(_0297_),
    .A2(net985));
 sg13g2_a21oi_2 _6486_ (.B1(_2507_),
    .Y(_2510_),
    .A2(_3230_),
    .A1(\vgademo.b_cos[3] ));
 sg13g2_xnor2_1 _6487_ (.Y(_2511_),
    .A(\vgademo.b_cos[4] ),
    .B(net1051));
 sg13g2_nor2b_1 _6488_ (.A(_2510_),
    .B_N(_2511_),
    .Y(_2512_));
 sg13g2_xor2_1 _6489_ (.B(_2511_),
    .A(_2510_),
    .X(_2513_));
 sg13g2_nor2_1 _6490_ (.A(net392),
    .B(net1027),
    .Y(_2514_));
 sg13g2_a221oi_1 _6491_ (.B2(_2513_),
    .C1(_2514_),
    .B1(net984),
    .A1(_3233_),
    .Y(_0298_),
    .A2(net987));
 sg13g2_xnor2_1 _6492_ (.Y(_2515_),
    .A(net1051),
    .B(\vgademo.b_cos[5] ));
 sg13g2_a21oi_1 _6493_ (.A1(\vgademo.b_cos[4] ),
    .A2(_3232_),
    .Y(_2516_),
    .B1(_2512_));
 sg13g2_a21o_1 _6494_ (.A2(net1027),
    .A1(\vgademo.a_cos[8] ),
    .B1(net983),
    .X(_2517_));
 sg13g2_xnor2_1 _6495_ (.Y(_2518_),
    .A(_2515_),
    .B(_2516_));
 sg13g2_o21ai_1 _6496_ (.B1(_2517_),
    .Y(_2519_),
    .A1(net1008),
    .A2(_2518_));
 sg13g2_o21ai_1 _6497_ (.B1(_2519_),
    .Y(_0299_),
    .A1(_3234_),
    .A2(net1027));
 sg13g2_o21ai_1 _6498_ (.B1(_3232_),
    .Y(_2520_),
    .A1(\vgademo.b_cos[4] ),
    .A2(\vgademo.b_cos[5] ));
 sg13g2_nand2_1 _6499_ (.Y(_2521_),
    .A(_2512_),
    .B(_2515_));
 sg13g2_xor2_1 _6500_ (.B(net1056),
    .A(net1050),
    .X(_2522_));
 sg13g2_a21oi_1 _6501_ (.A1(_2520_),
    .A2(_2521_),
    .Y(_2523_),
    .B1(_2522_));
 sg13g2_nand3_1 _6502_ (.B(_2521_),
    .C(_2522_),
    .A(_2520_),
    .Y(_2524_));
 sg13g2_nand2_1 _6503_ (.Y(_2525_),
    .A(net983),
    .B(_2524_));
 sg13g2_a22oi_1 _6504_ (.Y(_2526_),
    .B1(net986),
    .B2(net522),
    .A2(net1026),
    .A1(net1056));
 sg13g2_o21ai_1 _6505_ (.B1(_2526_),
    .Y(_0300_),
    .A1(_2523_),
    .A2(_2525_));
 sg13g2_xnor2_1 _6506_ (.Y(_2527_),
    .A(net1051),
    .B(\vgademo.b_cos[7] ));
 sg13g2_a21oi_1 _6507_ (.A1(_3232_),
    .A2(net1056),
    .Y(_2528_),
    .B1(_2523_));
 sg13g2_xnor2_1 _6508_ (.Y(_2529_),
    .A(_2527_),
    .B(_2528_));
 sg13g2_nand2_1 _6509_ (.Y(_2530_),
    .A(net461),
    .B(net986));
 sg13g2_a22oi_1 _6510_ (.Y(_2531_),
    .B1(net983),
    .B2(_2529_),
    .A2(net1024),
    .A1(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6511_ (.Y(_0301_),
    .A(_2530_),
    .B(_2531_));
 sg13g2_nand2b_1 _6512_ (.Y(_2532_),
    .B(_2527_),
    .A_N(_2522_));
 sg13g2_nor2_1 _6513_ (.A(_2521_),
    .B(_2532_),
    .Y(_2533_));
 sg13g2_o21ai_1 _6514_ (.B1(_3232_),
    .Y(_2534_),
    .A1(net1056),
    .A2(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6515_ (.Y(_2535_),
    .A(_2520_),
    .B(_2534_));
 sg13g2_nor2_1 _6516_ (.A(_2533_),
    .B(_2535_),
    .Y(_2536_));
 sg13g2_xnor2_1 _6517_ (.Y(_2537_),
    .A(net1050),
    .B(\vgademo.b_cos[8] ));
 sg13g2_o21ai_1 _6518_ (.B1(_2537_),
    .Y(_2538_),
    .A1(_2533_),
    .A2(_2535_));
 sg13g2_xnor2_1 _6519_ (.Y(_2539_),
    .A(_2536_),
    .B(_2537_));
 sg13g2_nand2_1 _6520_ (.Y(_2540_),
    .A(net439),
    .B(net986));
 sg13g2_a22oi_1 _6521_ (.Y(_2541_),
    .B1(net983),
    .B2(_2539_),
    .A2(net1024),
    .A1(\vgademo.b_cos[8] ));
 sg13g2_nand2_1 _6522_ (.Y(_0302_),
    .A(_2540_),
    .B(_2541_));
 sg13g2_o21ai_1 _6523_ (.B1(_2538_),
    .Y(_2542_),
    .A1(net1050),
    .A2(_3237_));
 sg13g2_nand2_1 _6524_ (.Y(_2543_),
    .A(net1050),
    .B(_3238_));
 sg13g2_nor2_1 _6525_ (.A(net1050),
    .B(_3238_),
    .Y(_2544_));
 sg13g2_xor2_1 _6526_ (.B(net1055),
    .A(net1050),
    .X(_2545_));
 sg13g2_xnor2_1 _6527_ (.Y(_2546_),
    .A(_2542_),
    .B(_2545_));
 sg13g2_nand2_1 _6528_ (.Y(_2547_),
    .A(net437),
    .B(net987));
 sg13g2_a22oi_1 _6529_ (.Y(_2548_),
    .B1(net983),
    .B2(_2546_),
    .A2(net1024),
    .A1(net1055));
 sg13g2_nand2_1 _6530_ (.Y(_0303_),
    .A(_2547_),
    .B(_2548_));
 sg13g2_nand2_1 _6531_ (.Y(_2549_),
    .A(_3232_),
    .B(net1054));
 sg13g2_xor2_1 _6532_ (.B(net1054),
    .A(net1050),
    .X(_2550_));
 sg13g2_a21oi_1 _6533_ (.A1(_2542_),
    .A2(_2543_),
    .Y(_2551_),
    .B1(_2544_));
 sg13g2_xor2_1 _6534_ (.B(_2551_),
    .A(_2550_),
    .X(_2552_));
 sg13g2_a22oi_1 _6535_ (.Y(_2553_),
    .B1(net983),
    .B2(_2552_),
    .A2(net987),
    .A1(net542));
 sg13g2_o21ai_1 _6536_ (.B1(_2553_),
    .Y(_0304_),
    .A1(_3239_),
    .A2(net1027));
 sg13g2_o21ai_1 _6537_ (.B1(_2549_),
    .Y(_2554_),
    .A1(_2550_),
    .A2(_2551_));
 sg13g2_xor2_1 _6538_ (.B(\vgademo.b_cos[11] ),
    .A(net1050),
    .X(_2555_));
 sg13g2_xnor2_1 _6539_ (.Y(_2556_),
    .A(_2554_),
    .B(_2555_));
 sg13g2_nand2_1 _6540_ (.Y(_2557_),
    .A(net422),
    .B(net987));
 sg13g2_a22oi_1 _6541_ (.Y(_2558_),
    .B1(net983),
    .B2(_2556_),
    .A2(net1024),
    .A1(\vgademo.b_cos[11] ));
 sg13g2_nand2_1 _6542_ (.Y(_0305_),
    .A(_2557_),
    .B(_2558_));
 sg13g2_mux2_1 _6543_ (.A0(net334),
    .A1(_0225_),
    .S(_0666_),
    .X(_0306_));
 sg13g2_nand2b_1 _6544_ (.Y(_2559_),
    .B(_1093_),
    .A_N(_1085_));
 sg13g2_a21oi_1 _6545_ (.A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ),
    .Y(_2560_),
    .B1(net1052));
 sg13g2_o21ai_1 _6546_ (.B1(_2560_),
    .Y(_2561_),
    .A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ));
 sg13g2_o21ai_1 _6547_ (.B1(_2561_),
    .Y(_2562_),
    .A1(_3172_),
    .A2(_0069_));
 sg13g2_nand2_1 _6548_ (.Y(_2563_),
    .A(net334),
    .B(_2562_));
 sg13g2_xnor2_1 _6549_ (.Y(_2564_),
    .A(net334),
    .B(_2562_));
 sg13g2_nand2_1 _6550_ (.Y(_2565_),
    .A(net1014),
    .B(_2564_));
 sg13g2_nand3_1 _6551_ (.B(_1094_),
    .C(_2565_),
    .A(_1085_),
    .Y(_2566_));
 sg13g2_a22oi_1 _6552_ (.Y(_0307_),
    .B1(_2559_),
    .B2(_2566_),
    .A2(net1012),
    .A1(_3206_));
 sg13g2_nand2_1 _6553_ (.Y(_2567_),
    .A(_1084_),
    .B(_1093_));
 sg13g2_nor2b_1 _6554_ (.A(_1105_),
    .B_N(_2567_),
    .Y(_2568_));
 sg13g2_xor2_1 _6555_ (.B(_2567_),
    .A(_1105_),
    .X(_2569_));
 sg13g2_nor2_1 _6556_ (.A(net338),
    .B(_0666_),
    .Y(_2570_));
 sg13g2_o21ai_1 _6557_ (.B1(\vgademo.plane_dx_div.d[18] ),
    .Y(_2571_),
    .A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ));
 sg13g2_or3_2 _6558_ (.A(\vgademo.plane_dx_div.d[16] ),
    .B(\vgademo.plane_dx_div.d[17] ),
    .C(\vgademo.plane_dx_div.d[18] ),
    .X(_2572_));
 sg13g2_a21oi_1 _6559_ (.A1(_2571_),
    .A2(_2572_),
    .Y(_2573_),
    .B1(net1052));
 sg13g2_a21oi_1 _6560_ (.A1(net1052),
    .A2(_0072_),
    .Y(_2574_),
    .B1(_2573_));
 sg13g2_nand2_1 _6561_ (.Y(_2575_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2574_));
 sg13g2_xnor2_1 _6562_ (.Y(_2576_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2574_));
 sg13g2_xnor2_1 _6563_ (.Y(_2577_),
    .A(_2563_),
    .B(_2576_));
 sg13g2_a221oi_1 _6564_ (.B2(net1015),
    .C1(_2570_),
    .B1(_2577_),
    .A1(net1031),
    .Y(_0308_),
    .A2(_2569_));
 sg13g2_nor2b_1 _6565_ (.A(_1119_),
    .B_N(_2568_),
    .Y(_2578_));
 sg13g2_xor2_1 _6566_ (.B(_2568_),
    .A(_1119_),
    .X(_2579_));
 sg13g2_nor2_1 _6567_ (.A(net344),
    .B(_0666_),
    .Y(_2580_));
 sg13g2_o21ai_1 _6568_ (.B1(_2575_),
    .Y(_2581_),
    .A1(_2563_),
    .A2(_2576_));
 sg13g2_a21oi_1 _6569_ (.A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2572_),
    .Y(_2582_),
    .B1(net1053));
 sg13g2_o21ai_1 _6570_ (.B1(_2582_),
    .Y(_2583_),
    .A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2572_));
 sg13g2_o21ai_1 _6571_ (.B1(_2583_),
    .Y(_2584_),
    .A1(_3172_),
    .A2(_0075_));
 sg13g2_and2_1 _6572_ (.A(\vgademo.plane_dx_div.r[18] ),
    .B(_2584_),
    .X(_2585_));
 sg13g2_xor2_1 _6573_ (.B(_2584_),
    .A(net338),
    .X(_2586_));
 sg13g2_xnor2_1 _6574_ (.Y(_2587_),
    .A(_2581_),
    .B(_2586_));
 sg13g2_a221oi_1 _6575_ (.B2(net1015),
    .C1(_2580_),
    .B1(_2587_),
    .A1(net1030),
    .Y(_0309_),
    .A2(_2579_));
 sg13g2_nand2_1 _6576_ (.Y(_2588_),
    .A(_1135_),
    .B(_2578_));
 sg13g2_xnor2_1 _6577_ (.Y(_2589_),
    .A(_1135_),
    .B(_2578_));
 sg13g2_nor2_1 _6578_ (.A(net262),
    .B(_0666_),
    .Y(_2590_));
 sg13g2_a21oi_2 _6579_ (.B1(_2585_),
    .Y(_2591_),
    .A2(_2586_),
    .A1(_2581_));
 sg13g2_o21ai_1 _6580_ (.B1(\vgademo.plane_dx_div.d[20] ),
    .Y(_2592_),
    .A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2572_));
 sg13g2_or3_2 _6581_ (.A(\vgademo.plane_dx_div.d[19] ),
    .B(\vgademo.plane_dx_div.d[20] ),
    .C(_2572_),
    .X(_2593_));
 sg13g2_a21oi_1 _6582_ (.A1(_2592_),
    .A2(_2593_),
    .Y(_2594_),
    .B1(net1053));
 sg13g2_a21oi_1 _6583_ (.A1(net1053),
    .A2(_0078_),
    .Y(_2595_),
    .B1(_2594_));
 sg13g2_nand2_1 _6584_ (.Y(_2596_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .B(_2595_));
 sg13g2_xnor2_1 _6585_ (.Y(_2597_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .B(_2595_));
 sg13g2_xnor2_1 _6586_ (.Y(_2598_),
    .A(_2591_),
    .B(_2597_));
 sg13g2_a221oi_1 _6587_ (.B2(net1014),
    .C1(_2590_),
    .B1(_2598_),
    .A1(net1030),
    .Y(_0310_),
    .A2(_2589_));
 sg13g2_nor2_1 _6588_ (.A(_1149_),
    .B(_2588_),
    .Y(_2599_));
 sg13g2_xnor2_1 _6589_ (.Y(_2600_),
    .A(_1149_),
    .B(_2588_));
 sg13g2_nor2_1 _6590_ (.A(net299),
    .B(_0666_),
    .Y(_2601_));
 sg13g2_o21ai_1 _6591_ (.B1(_2596_),
    .Y(_2602_),
    .A1(_2591_),
    .A2(_2597_));
 sg13g2_xor2_1 _6592_ (.B(_2593_),
    .A(\vgademo.plane_dx_div.d[21] ),
    .X(_2603_));
 sg13g2_nor2_1 _6593_ (.A(net1052),
    .B(_2603_),
    .Y(_2604_));
 sg13g2_and2_1 _6594_ (.A(net1052),
    .B(_0080_),
    .X(_2605_));
 sg13g2_nor3_1 _6595_ (.A(_3208_),
    .B(_2604_),
    .C(_2605_),
    .Y(_2606_));
 sg13g2_o21ai_1 _6596_ (.B1(_3208_),
    .Y(_2607_),
    .A1(_2604_),
    .A2(_2605_));
 sg13g2_nor2b_1 _6597_ (.A(_2606_),
    .B_N(_2607_),
    .Y(_2608_));
 sg13g2_xnor2_1 _6598_ (.Y(_2609_),
    .A(_2602_),
    .B(_2608_));
 sg13g2_a221oi_1 _6599_ (.B2(net1014),
    .C1(_2601_),
    .B1(_2609_),
    .A1(net1030),
    .Y(_0311_),
    .A2(_2600_));
 sg13g2_nand2_1 _6600_ (.Y(_2610_),
    .A(_1170_),
    .B(_2599_));
 sg13g2_xnor2_1 _6601_ (.Y(_2611_),
    .A(_1170_),
    .B(_2599_));
 sg13g2_a21oi_1 _6602_ (.A1(_2602_),
    .A2(_2607_),
    .Y(_2612_),
    .B1(_2606_));
 sg13g2_nand2b_1 _6603_ (.Y(_2613_),
    .B(net1052),
    .A_N(_0013_));
 sg13g2_o21ai_1 _6604_ (.B1(\vgademo.plane_dx_div.d[22] ),
    .Y(_2614_),
    .A1(\vgademo.plane_dx_div.d[21] ),
    .A2(_2593_));
 sg13g2_nor3_1 _6605_ (.A(\vgademo.plane_dx_div.d[21] ),
    .B(\vgademo.plane_dx_div.d[22] ),
    .C(_2593_),
    .Y(_2615_));
 sg13g2_nand2_1 _6606_ (.Y(_2616_),
    .A(_3172_),
    .B(_2614_));
 sg13g2_o21ai_1 _6607_ (.B1(_2613_),
    .Y(_2617_),
    .A1(_2615_),
    .A2(_2616_));
 sg13g2_nor2_1 _6608_ (.A(\vgademo.plane_dx_div.r[21] ),
    .B(_2617_),
    .Y(_2618_));
 sg13g2_and2_1 _6609_ (.A(\vgademo.plane_dx_div.r[21] ),
    .B(_2617_),
    .X(_2619_));
 sg13g2_nor2_1 _6610_ (.A(_2618_),
    .B(_2619_),
    .Y(_2620_));
 sg13g2_o21ai_1 _6611_ (.B1(net1014),
    .Y(_2621_),
    .A1(_2612_),
    .A2(_2620_));
 sg13g2_a21oi_1 _6612_ (.A1(_2612_),
    .A2(_2620_),
    .Y(_2622_),
    .B1(_2621_));
 sg13g2_a221oi_1 _6613_ (.B2(net1030),
    .C1(_2622_),
    .B1(_2611_),
    .A1(_3211_),
    .Y(_0312_),
    .A2(net1013));
 sg13g2_nand2_1 _6614_ (.Y(_2623_),
    .A(_1187_),
    .B(_2610_));
 sg13g2_nor2_1 _6615_ (.A(_1187_),
    .B(_2610_),
    .Y(_2624_));
 sg13g2_nand3b_1 _6616_ (.B(net1032),
    .C(_2623_),
    .Y(_2625_),
    .A_N(_2624_));
 sg13g2_nand2b_1 _6617_ (.Y(_2626_),
    .B(\vgademo.plane_dx_div.d[23] ),
    .A_N(_2615_));
 sg13g2_nand2b_1 _6618_ (.Y(_2627_),
    .B(_2615_),
    .A_N(\vgademo.plane_dx_div.d[23] ));
 sg13g2_nand3_1 _6619_ (.B(_2626_),
    .C(_2627_),
    .A(_3172_),
    .Y(_2628_));
 sg13g2_o21ai_1 _6620_ (.B1(_2628_),
    .Y(_2629_),
    .A1(_3172_),
    .A2(_0017_));
 sg13g2_and2_1 _6621_ (.A(\vgademo.plane_dx_div.r[22] ),
    .B(_2629_),
    .X(_2630_));
 sg13g2_xnor2_1 _6622_ (.Y(_2631_),
    .A(_3211_),
    .B(_2629_));
 sg13g2_nor2b_1 _6623_ (.A(_2619_),
    .B_N(_2612_),
    .Y(_2632_));
 sg13g2_nor2_1 _6624_ (.A(_2618_),
    .B(_2632_),
    .Y(_2633_));
 sg13g2_or2_1 _6625_ (.X(_2634_),
    .B(_2633_),
    .A(_2631_));
 sg13g2_and2_1 _6626_ (.A(_2631_),
    .B(_2633_),
    .X(_2635_));
 sg13g2_nor2_1 _6627_ (.A(net1032),
    .B(_2635_),
    .Y(_2636_));
 sg13g2_a21oi_1 _6628_ (.A1(_2634_),
    .A2(_2636_),
    .Y(_2637_),
    .B1(net1013));
 sg13g2_a22oi_1 _6629_ (.Y(_0313_),
    .B1(_2625_),
    .B2(_2637_),
    .A2(net1013),
    .A1(_3216_));
 sg13g2_o21ai_1 _6630_ (.B1(_1198_),
    .Y(_2638_),
    .A1(_1187_),
    .A2(_2610_));
 sg13g2_nand2_1 _6631_ (.Y(_2639_),
    .A(\vgademo.plane_dx_div.d[24] ),
    .B(_2627_));
 sg13g2_nor2_1 _6632_ (.A(\vgademo.plane_dx_div.d[24] ),
    .B(_2627_),
    .Y(_2640_));
 sg13g2_nor2_1 _6633_ (.A(net1052),
    .B(_2640_),
    .Y(_2641_));
 sg13g2_a22oi_1 _6634_ (.Y(_2642_),
    .B1(_2639_),
    .B2(_2641_),
    .A2(_3215_),
    .A1(net1052));
 sg13g2_xnor2_1 _6635_ (.Y(_2643_),
    .A(\vgademo.plane_dx_div.r[23] ),
    .B(_2642_));
 sg13g2_nor3_1 _6636_ (.A(_2630_),
    .B(_2635_),
    .C(_2643_),
    .Y(_2644_));
 sg13g2_o21ai_1 _6637_ (.B1(_2643_),
    .Y(_2645_),
    .A1(_2630_),
    .A2(_2635_));
 sg13g2_nor2b_1 _6638_ (.A(_2644_),
    .B_N(_2645_),
    .Y(_2646_));
 sg13g2_o21ai_1 _6639_ (.B1(_1199_),
    .Y(_2647_),
    .A1(_0663_),
    .A2(_2624_));
 sg13g2_a221oi_1 _6640_ (.B2(_2638_),
    .C1(net1012),
    .B1(_2647_),
    .A1(_0663_),
    .Y(_2648_),
    .A2(_2646_));
 sg13g2_a21oi_1 _6641_ (.A1(_3217_),
    .A2(net1012),
    .Y(_0314_),
    .B1(_2648_));
 sg13g2_o21ai_1 _6642_ (.B1(_2645_),
    .Y(_2649_),
    .A1(_3216_),
    .A2(_2642_));
 sg13g2_xnor2_1 _6643_ (.Y(_2650_),
    .A(_3217_),
    .B(_2641_));
 sg13g2_xnor2_1 _6644_ (.Y(_2651_),
    .A(_2649_),
    .B(_2650_));
 sg13g2_nor2_1 _6645_ (.A(net1032),
    .B(_2651_),
    .Y(_2652_));
 sg13g2_nor3_1 _6646_ (.A(net1012),
    .B(_2647_),
    .C(_2652_),
    .Y(_2653_));
 sg13g2_a21oi_1 _6647_ (.A1(_3172_),
    .A2(net1013),
    .Y(_0315_),
    .B1(_2653_));
 sg13g2_o21ai_1 _6648_ (.B1(_1914_),
    .Y(_2654_),
    .A1(_1858_),
    .A2(_1870_));
 sg13g2_nand3_1 _6649_ (.B(net896),
    .C(_2654_),
    .A(net955),
    .Y(_2655_));
 sg13g2_and2_1 _6650_ (.A(_1803_),
    .B(_2196_),
    .X(_2656_));
 sg13g2_nor2_1 _6651_ (.A(_2212_),
    .B(_2236_),
    .Y(_2657_));
 sg13g2_nor2_1 _6652_ (.A(_2208_),
    .B(_2657_),
    .Y(_2658_));
 sg13g2_a221oi_1 _6653_ (.B2(_1802_),
    .C1(net963),
    .B1(_2658_),
    .A1(_2655_),
    .Y(_2659_),
    .A2(_2656_));
 sg13g2_and2_1 _6654_ (.A(_1295_),
    .B(_1316_),
    .X(_2660_));
 sg13g2_nor2_2 _6655_ (.A(_2659_),
    .B(_2660_),
    .Y(_2661_));
 sg13g2_a22oi_1 _6656_ (.Y(_2662_),
    .B1(net905),
    .B2(_2222_),
    .A2(_1912_),
    .A1(_1863_));
 sg13g2_o21ai_1 _6657_ (.B1(net955),
    .Y(_2663_),
    .A1(_1824_),
    .A2(_2662_));
 sg13g2_a21oi_1 _6658_ (.A1(net951),
    .A2(_2218_),
    .Y(_2664_),
    .B1(_1802_));
 sg13g2_nand2_1 _6659_ (.Y(_2665_),
    .A(_2663_),
    .B(_2664_));
 sg13g2_nor2_1 _6660_ (.A(net898),
    .B(_2239_),
    .Y(_2666_));
 sg13g2_nand2b_1 _6661_ (.Y(_2667_),
    .B(_2666_),
    .A_N(_2657_));
 sg13g2_and3_1 _6662_ (.X(_2668_),
    .A(net962),
    .B(_2665_),
    .C(_2667_));
 sg13g2_nand3_1 _6663_ (.B(_2665_),
    .C(_2667_),
    .A(net961),
    .Y(_2669_));
 sg13g2_a21o_1 _6664_ (.A2(_2668_),
    .A1(_2228_),
    .B1(_2661_),
    .X(_2670_));
 sg13g2_o21ai_1 _6665_ (.B1(_2661_),
    .Y(_2671_),
    .A1(_2228_),
    .A2(_2668_));
 sg13g2_nand2_1 _6666_ (.Y(_2672_),
    .A(_2670_),
    .B(_2671_));
 sg13g2_a21oi_2 _6667_ (.B1(_2221_),
    .Y(_2673_),
    .A2(_2248_),
    .A1(net905));
 sg13g2_nor4_1 _6668_ (.A(net902),
    .B(net899),
    .C(net947),
    .D(_2654_),
    .Y(_2674_));
 sg13g2_a221oi_1 _6669_ (.B2(_2673_),
    .C1(_2674_),
    .B1(net897),
    .A1(net957),
    .Y(_2675_),
    .A2(net960));
 sg13g2_o21ai_1 _6670_ (.B1(net898),
    .Y(_2676_),
    .A1(_2254_),
    .A2(_2675_));
 sg13g2_nand2_1 _6671_ (.Y(_2677_),
    .A(_2241_),
    .B(_2676_));
 sg13g2_a21oi_1 _6672_ (.A1(_2241_),
    .A2(_2676_),
    .Y(_2678_),
    .B1(_2227_));
 sg13g2_a21o_1 _6673_ (.A2(_2676_),
    .A1(_2241_),
    .B1(_2227_),
    .X(_2679_));
 sg13g2_nand3_1 _6674_ (.B(_2241_),
    .C(_2676_),
    .A(net1040),
    .Y(_2680_));
 sg13g2_and3_1 _6675_ (.X(_2681_),
    .A(_2669_),
    .B(_2679_),
    .C(_2680_));
 sg13g2_or2_1 _6676_ (.X(_2682_),
    .B(_2681_),
    .A(_2678_));
 sg13g2_xnor2_1 _6677_ (.Y(_2683_),
    .A(_2229_),
    .B(_2668_));
 sg13g2_xnor2_1 _6678_ (.Y(_2684_),
    .A(_2661_),
    .B(_2683_));
 sg13g2_nor2_1 _6679_ (.A(_2682_),
    .B(_2684_),
    .Y(_2685_));
 sg13g2_nor4_1 _6680_ (.A(net902),
    .B(net899),
    .C(net947),
    .D(_2662_),
    .Y(_2686_));
 sg13g2_and2_1 _6681_ (.A(_2247_),
    .B(_2271_),
    .X(_2687_));
 sg13g2_nand2_1 _6682_ (.Y(_2688_),
    .A(_2247_),
    .B(_2271_));
 sg13g2_a221oi_1 _6683_ (.B2(_2688_),
    .C1(_2686_),
    .B1(net897),
    .A1(net957),
    .Y(_2689_),
    .A2(net960));
 sg13g2_nor3_1 _6684_ (.A(_2208_),
    .B(_2212_),
    .C(_2236_),
    .Y(_2690_));
 sg13g2_a221oi_1 _6685_ (.B2(_1802_),
    .C1(net963),
    .B1(_2690_),
    .A1(_2210_),
    .Y(_2691_),
    .A2(_2213_));
 sg13g2_nand3b_1 _6686_ (.B(_1802_),
    .C(_2209_),
    .Y(_2692_),
    .A_N(_2236_));
 sg13g2_o21ai_1 _6687_ (.B1(_2691_),
    .Y(_2693_),
    .A1(_2301_),
    .A2(_2689_));
 sg13g2_and2_1 _6688_ (.A(_2307_),
    .B(_2693_),
    .X(_2694_));
 sg13g2_xor2_1 _6689_ (.B(_2693_),
    .A(_2307_),
    .X(_2695_));
 sg13g2_a21oi_1 _6690_ (.A1(_2677_),
    .A2(_2695_),
    .Y(_2696_),
    .B1(_2694_));
 sg13g2_a21oi_1 _6691_ (.A1(_2679_),
    .A2(_2680_),
    .Y(_2697_),
    .B1(_2669_));
 sg13g2_nor3_1 _6692_ (.A(_2681_),
    .B(_2696_),
    .C(_2697_),
    .Y(_2698_));
 sg13g2_or3_1 _6693_ (.A(_2681_),
    .B(_2696_),
    .C(_2697_),
    .X(_2699_));
 sg13g2_o21ai_1 _6694_ (.B1(_2696_),
    .Y(_2700_),
    .A1(_2681_),
    .A2(_2697_));
 sg13g2_nand2_1 _6695_ (.Y(_2701_),
    .A(_2267_),
    .B(_2289_));
 sg13g2_nor4_1 _6696_ (.A(net904),
    .B(net901),
    .C(net948),
    .D(_2687_),
    .Y(_2702_));
 sg13g2_a221oi_1 _6697_ (.B2(_2701_),
    .C1(_2702_),
    .B1(net897),
    .A1(net958),
    .Y(_2703_),
    .A2(net960));
 sg13g2_o21ai_1 _6698_ (.B1(net962),
    .Y(_2704_),
    .A1(_2278_),
    .A2(_2703_));
 sg13g2_and2_1 _6699_ (.A(_2266_),
    .B(_2704_),
    .X(_2705_));
 sg13g2_nand2_1 _6700_ (.Y(_2706_),
    .A(_2270_),
    .B(_2290_));
 sg13g2_nor4_1 _6701_ (.A(net902),
    .B(net899),
    .C(net947),
    .D(_2673_),
    .Y(_2707_));
 sg13g2_a221oi_1 _6702_ (.B2(_2706_),
    .C1(_2707_),
    .B1(net897),
    .A1(net957),
    .Y(_2708_),
    .A2(_1339_));
 sg13g2_o21ai_1 _6703_ (.B1(net962),
    .Y(_2709_),
    .A1(_2285_),
    .A2(_2708_));
 sg13g2_xor2_1 _6704_ (.B(_2704_),
    .A(_2266_),
    .X(_2710_));
 sg13g2_a21o_1 _6705_ (.A2(_2710_),
    .A1(_2709_),
    .B1(_2705_),
    .X(_2711_));
 sg13g2_xnor2_1 _6706_ (.Y(_2712_),
    .A(_2677_),
    .B(_2695_));
 sg13g2_a21o_1 _6707_ (.A2(_2659_),
    .A1(_2312_),
    .B1(_2709_),
    .X(_2713_));
 sg13g2_or3_1 _6708_ (.A(_2312_),
    .B(_2659_),
    .C(_2660_),
    .X(_2714_));
 sg13g2_a21oi_1 _6709_ (.A1(_2713_),
    .A2(_2714_),
    .Y(_2715_),
    .B1(_2693_));
 sg13g2_nor2b_1 _6710_ (.A(_2712_),
    .B_N(_2711_),
    .Y(_2716_));
 sg13g2_xnor2_1 _6711_ (.Y(_2717_),
    .A(_2709_),
    .B(_2710_));
 sg13g2_nand3_1 _6712_ (.B(_2713_),
    .C(_2714_),
    .A(_2693_),
    .Y(_2718_));
 sg13g2_xnor2_1 _6713_ (.Y(_2719_),
    .A(_2711_),
    .B(_2712_));
 sg13g2_a21oi_1 _6714_ (.A1(_2717_),
    .A2(_2718_),
    .Y(_2720_),
    .B1(_2715_));
 sg13g2_nand4_1 _6715_ (.B(_2700_),
    .C(_2719_),
    .A(_2699_),
    .Y(_2721_),
    .D(_2720_));
 sg13g2_a221oi_1 _6716_ (.B2(_2716_),
    .C1(_2698_),
    .B1(_2700_),
    .A1(_2682_),
    .Y(_2722_),
    .A2(_2684_));
 sg13g2_a21o_1 _6717_ (.A2(_2722_),
    .A1(_2721_),
    .B1(_2685_),
    .X(_2723_));
 sg13g2_or2_1 _6718_ (.X(_2724_),
    .B(_2723_),
    .A(_2672_));
 sg13g2_a21oi_1 _6719_ (.A1(_2672_),
    .A2(_2723_),
    .Y(_2725_),
    .B1(_2336_));
 sg13g2_and2_1 _6720_ (.A(_2724_),
    .B(_2725_),
    .X(_0316_));
 sg13g2_a21oi_1 _6721_ (.A1(_2670_),
    .A2(_2724_),
    .Y(_0317_),
    .B1(_2336_));
 sg13g2_nand2_1 _6722_ (.Y(_2726_),
    .A(\vgademo.b_sin[0] ),
    .B(_2529_));
 sg13g2_xnor2_1 _6723_ (.Y(_2727_),
    .A(net411),
    .B(_2529_));
 sg13g2_a22oi_1 _6724_ (.Y(_2728_),
    .B1(net986),
    .B2(net324),
    .A2(net1026),
    .A1(net411));
 sg13g2_o21ai_1 _6725_ (.B1(_2728_),
    .Y(_0318_),
    .A1(_2492_),
    .A2(_2727_));
 sg13g2_xnor2_1 _6726_ (.Y(_2729_),
    .A(net363),
    .B(_2539_));
 sg13g2_nor2_1 _6727_ (.A(_2726_),
    .B(_2729_),
    .Y(_2730_));
 sg13g2_a21o_1 _6728_ (.A2(_2729_),
    .A1(_2726_),
    .B1(_2492_),
    .X(_2731_));
 sg13g2_a22oi_1 _6729_ (.Y(_2732_),
    .B1(net986),
    .B2(net355),
    .A2(net1024),
    .A1(net363));
 sg13g2_o21ai_1 _6730_ (.B1(_2732_),
    .Y(_0319_),
    .A1(_2730_),
    .A2(_2731_));
 sg13g2_a21oi_1 _6731_ (.A1(net363),
    .A2(_2539_),
    .Y(_2733_),
    .B1(_2730_));
 sg13g2_nand2_1 _6732_ (.Y(_2734_),
    .A(net382),
    .B(_2546_));
 sg13g2_xnor2_1 _6733_ (.Y(_2735_),
    .A(net382),
    .B(_2546_));
 sg13g2_or2_1 _6734_ (.X(_2736_),
    .B(_2735_),
    .A(_2733_));
 sg13g2_a21oi_1 _6735_ (.A1(_2733_),
    .A2(_2735_),
    .Y(_2737_),
    .B1(_2492_));
 sg13g2_nand2_1 _6736_ (.Y(_2738_),
    .A(_2736_),
    .B(_2737_));
 sg13g2_a22oi_1 _6737_ (.Y(_2739_),
    .B1(net986),
    .B2(net311),
    .A2(net1024),
    .A1(net382));
 sg13g2_nand2_1 _6738_ (.Y(_0320_),
    .A(_2738_),
    .B(_2739_));
 sg13g2_nand2_1 _6739_ (.Y(_2740_),
    .A(net389),
    .B(_2552_));
 sg13g2_xnor2_1 _6740_ (.Y(_2741_),
    .A(\vgademo.b_sin[3] ),
    .B(_2552_));
 sg13g2_nand3_1 _6741_ (.B(_2736_),
    .C(_2741_),
    .A(_2734_),
    .Y(_2742_));
 sg13g2_a21o_1 _6742_ (.A2(_2736_),
    .A1(_2734_),
    .B1(_2741_),
    .X(_2743_));
 sg13g2_nand3_1 _6743_ (.B(_2742_),
    .C(_2743_),
    .A(net984),
    .Y(_2744_));
 sg13g2_a22oi_1 _6744_ (.Y(_2745_),
    .B1(net986),
    .B2(\vgademo.a_sin[6] ),
    .A2(net1026),
    .A1(net389));
 sg13g2_nand2_1 _6745_ (.Y(_0321_),
    .A(_2744_),
    .B(net390));
 sg13g2_nand2_1 _6746_ (.Y(_2746_),
    .A(\vgademo.b_sin[4] ),
    .B(net915));
 sg13g2_xnor2_1 _6747_ (.Y(_2747_),
    .A(\vgademo.b_sin[4] ),
    .B(_2556_));
 sg13g2_a21o_2 _6748_ (.A2(_2743_),
    .A1(_2740_),
    .B1(_2747_),
    .X(_2748_));
 sg13g2_nand3_1 _6749_ (.B(_2743_),
    .C(_2747_),
    .A(_2740_),
    .Y(_2749_));
 sg13g2_nand3_1 _6750_ (.B(_2748_),
    .C(_2749_),
    .A(net983),
    .Y(_2750_));
 sg13g2_a22oi_1 _6751_ (.Y(_2751_),
    .B1(net986),
    .B2(\vgademo.a_sin[7] ),
    .A2(net1024),
    .A1(net493));
 sg13g2_nand2_1 _6752_ (.Y(_0322_),
    .A(_2750_),
    .B(net494));
 sg13g2_nand2_1 _6753_ (.Y(_2752_),
    .A(net283),
    .B(net1025));
 sg13g2_xnor2_1 _6754_ (.Y(_2753_),
    .A(\vgademo.b_sin[5] ),
    .B(net915));
 sg13g2_nand2_1 _6755_ (.Y(_2754_),
    .A(_2746_),
    .B(_2748_));
 sg13g2_o21ai_1 _6756_ (.B1(net1006),
    .Y(_2755_),
    .A1(_2753_),
    .A2(_2754_));
 sg13g2_a21oi_1 _6757_ (.A1(_2753_),
    .A2(_2754_),
    .Y(_2756_),
    .B1(_2755_));
 sg13g2_o21ai_1 _6758_ (.B1(net1027),
    .Y(_2757_),
    .A1(\vgademo.a_sin[8] ),
    .A2(net1006));
 sg13g2_o21ai_1 _6759_ (.B1(_2752_),
    .Y(_0323_),
    .A1(_2756_),
    .A2(_2757_));
 sg13g2_o21ai_1 _6760_ (.B1(net913),
    .Y(_2758_),
    .A1(\vgademo.b_sin[4] ),
    .A2(\vgademo.b_sin[5] ));
 sg13g2_o21ai_1 _6761_ (.B1(_2758_),
    .Y(_2759_),
    .A1(_2748_),
    .A2(_2753_));
 sg13g2_xnor2_1 _6762_ (.Y(_2760_),
    .A(\vgademo.b_sin[6] ),
    .B(net913));
 sg13g2_inv_1 _6763_ (.Y(_2761_),
    .A(_2760_));
 sg13g2_and2_1 _6764_ (.A(_2759_),
    .B(_2761_),
    .X(_2762_));
 sg13g2_o21ai_1 _6765_ (.B1(net984),
    .Y(_2763_),
    .A1(_2759_),
    .A2(_2761_));
 sg13g2_a22oi_1 _6766_ (.Y(_2764_),
    .B1(net985),
    .B2(\vgademo.a_sin[9] ),
    .A2(net1025),
    .A1(net426));
 sg13g2_o21ai_1 _6767_ (.B1(net427),
    .Y(_0324_),
    .A1(_2762_),
    .A2(_2763_));
 sg13g2_nand2_1 _6768_ (.Y(_2765_),
    .A(net307),
    .B(net1025));
 sg13g2_a21oi_1 _6769_ (.A1(\vgademo.b_sin[6] ),
    .A2(net913),
    .Y(_2766_),
    .B1(_2762_));
 sg13g2_xnor2_1 _6770_ (.Y(_2767_),
    .A(_3227_),
    .B(net913));
 sg13g2_o21ai_1 _6771_ (.B1(net1006),
    .Y(_2768_),
    .A1(_2766_),
    .A2(_2767_));
 sg13g2_a21oi_1 _6772_ (.A1(_2766_),
    .A2(_2767_),
    .Y(_2769_),
    .B1(_2768_));
 sg13g2_o21ai_1 _6773_ (.B1(net1027),
    .Y(_2770_),
    .A1(\vgademo.a_sin[10] ),
    .A2(net1006));
 sg13g2_o21ai_1 _6774_ (.B1(_2765_),
    .Y(_0325_),
    .A1(_2769_),
    .A2(_2770_));
 sg13g2_nor3_1 _6775_ (.A(_2748_),
    .B(_2753_),
    .C(_2760_),
    .Y(_2771_));
 sg13g2_o21ai_1 _6776_ (.B1(_2771_),
    .Y(_2772_),
    .A1(\vgademo.b_sin[7] ),
    .A2(net913));
 sg13g2_o21ai_1 _6777_ (.B1(net913),
    .Y(_2773_),
    .A1(\vgademo.b_sin[7] ),
    .A2(\vgademo.b_sin[6] ));
 sg13g2_and3_1 _6778_ (.X(_2774_),
    .A(_2758_),
    .B(_2772_),
    .C(_2773_));
 sg13g2_xnor2_1 _6779_ (.Y(_2775_),
    .A(\vgademo.b_sin[8] ),
    .B(net913));
 sg13g2_nor2_1 _6780_ (.A(_2774_),
    .B(_2775_),
    .Y(_2776_));
 sg13g2_a21o_1 _6781_ (.A2(_2775_),
    .A1(_2774_),
    .B1(_2492_),
    .X(_2777_));
 sg13g2_a22oi_1 _6782_ (.Y(_2778_),
    .B1(net985),
    .B2(net451),
    .A2(net1025),
    .A1(net486));
 sg13g2_o21ai_1 _6783_ (.B1(_2778_),
    .Y(_0326_),
    .A1(_2776_),
    .A2(_2777_));
 sg13g2_a21oi_1 _6784_ (.A1(\vgademo.b_sin[8] ),
    .A2(net913),
    .Y(_2779_),
    .B1(_2776_));
 sg13g2_nand2_1 _6785_ (.Y(_2780_),
    .A(\vgademo.b_sin[9] ),
    .B(net914));
 sg13g2_nor2_1 _6786_ (.A(\vgademo.b_sin[9] ),
    .B(net914),
    .Y(_2781_));
 sg13g2_xnor2_1 _6787_ (.Y(_2782_),
    .A(\vgademo.b_sin[9] ),
    .B(net914));
 sg13g2_xnor2_1 _6788_ (.Y(_2783_),
    .A(_2779_),
    .B(_2782_));
 sg13g2_a22oi_1 _6789_ (.Y(_2784_),
    .B1(net987),
    .B2(net497),
    .A2(net1025),
    .A1(\vgademo.b_sin[9] ));
 sg13g2_o21ai_1 _6790_ (.B1(net498),
    .Y(_0327_),
    .A1(_2492_),
    .A2(_2783_));
 sg13g2_xnor2_1 _6791_ (.Y(_2785_),
    .A(\vgademo.b_sin[10] ),
    .B(net914));
 sg13g2_or2_1 _6792_ (.X(_2786_),
    .B(_2781_),
    .A(_2779_));
 sg13g2_nand3_1 _6793_ (.B(_2785_),
    .C(_2786_),
    .A(_2780_),
    .Y(_2787_));
 sg13g2_a21oi_1 _6794_ (.A1(_2780_),
    .A2(_2786_),
    .Y(_2788_),
    .B1(_2785_));
 sg13g2_nand2_1 _6795_ (.Y(_2789_),
    .A(net984),
    .B(_2787_));
 sg13g2_a22oi_1 _6796_ (.Y(_2790_),
    .B1(net985),
    .B2(\vgademo.a_sin[13] ),
    .A2(net1025),
    .A1(net480));
 sg13g2_o21ai_1 _6797_ (.B1(net481),
    .Y(_0328_),
    .A1(_2788_),
    .A2(_2789_));
 sg13g2_nand2_1 _6798_ (.Y(_2791_),
    .A(net1051),
    .B(net1024));
 sg13g2_a21o_1 _6799_ (.A2(net914),
    .A1(\vgademo.b_sin[10] ),
    .B1(_2788_),
    .X(_2792_));
 sg13g2_xor2_1 _6800_ (.B(_2554_),
    .A(\vgademo.b_cos[11] ),
    .X(_2793_));
 sg13g2_o21ai_1 _6801_ (.B1(net1002),
    .Y(_2794_),
    .A1(_2792_),
    .A2(_2793_));
 sg13g2_a21oi_1 _6802_ (.A1(_2792_),
    .A2(_2793_),
    .Y(_2795_),
    .B1(_2794_));
 sg13g2_o21ai_1 _6803_ (.B1(net1027),
    .Y(_2796_),
    .A1(net1058),
    .A2(net1002));
 sg13g2_o21ai_1 _6804_ (.B1(_2791_),
    .Y(_0329_),
    .A1(_2795_),
    .A2(_2796_));
 sg13g2_nand2_1 _6805_ (.Y(_2797_),
    .A(net1007),
    .B(_2333_));
 sg13g2_nand2_2 _6806_ (.Y(_2798_),
    .A(net1182),
    .B(_2797_));
 sg13g2_inv_4 _6807_ (.A(net970),
    .Y(_2799_));
 sg13g2_nand2_1 _6808_ (.Y(_2800_),
    .A(net233),
    .B(\vgademo.plane_du[0] ));
 sg13g2_nand2_1 _6809_ (.Y(_2801_),
    .A(net290),
    .B(net305));
 sg13g2_xor2_1 _6810_ (.B(\vgademo.plane_du[1] ),
    .A(\vgademo.plane_u[1] ),
    .X(_2802_));
 sg13g2_nand2b_1 _6811_ (.Y(_2803_),
    .B(_2802_),
    .A_N(_2800_));
 sg13g2_xor2_1 _6812_ (.B(_2802_),
    .A(_2800_),
    .X(_2804_));
 sg13g2_nor2_1 _6813_ (.A(net1010),
    .B(_2804_),
    .Y(_2805_));
 sg13g2_a21oi_1 _6814_ (.A1(\vgademo.plane_dx[0] ),
    .A2(net1010),
    .Y(_2806_),
    .B1(_2805_));
 sg13g2_nand2_1 _6815_ (.Y(_2807_),
    .A(net290),
    .B(net973));
 sg13g2_o21ai_1 _6816_ (.B1(_2807_),
    .Y(_0330_),
    .A1(net972),
    .A2(_2806_));
 sg13g2_nand2_1 _6817_ (.Y(_2808_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_xnor2_1 _6818_ (.Y(_2809_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_nand3_1 _6819_ (.B(_2803_),
    .C(_2809_),
    .A(_2801_),
    .Y(_2810_));
 sg13g2_a21o_1 _6820_ (.A2(_2803_),
    .A1(_2801_),
    .B1(_2809_),
    .X(_2811_));
 sg13g2_nand3_1 _6821_ (.B(_2810_),
    .C(_2811_),
    .A(net1004),
    .Y(_2812_));
 sg13g2_nand2_1 _6822_ (.Y(_2813_),
    .A(_3165_),
    .B(net1053));
 sg13g2_xnor2_1 _6823_ (.Y(_2814_),
    .A(\vgademo.plane_dx[1] ),
    .B(net1053));
 sg13g2_a21oi_1 _6824_ (.A1(net1009),
    .A2(_2814_),
    .Y(_2815_),
    .B1(net972));
 sg13g2_a22oi_1 _6825_ (.Y(_0331_),
    .B1(_2812_),
    .B2(_2815_),
    .A2(net972),
    .A1(_3246_));
 sg13g2_nand2_1 _6826_ (.Y(_2816_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_xnor2_1 _6827_ (.Y(_2817_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_nand3_1 _6828_ (.B(_2811_),
    .C(_2817_),
    .A(_2808_),
    .Y(_2818_));
 sg13g2_a21o_1 _6829_ (.A2(_2811_),
    .A1(_2808_),
    .B1(_2817_),
    .X(_2819_));
 sg13g2_nor2_1 _6830_ (.A(\vgademo.plane_dx[2] ),
    .B(_2813_),
    .Y(_2820_));
 sg13g2_xnor2_1 _6831_ (.Y(_2821_),
    .A(\vgademo.plane_dx[2] ),
    .B(_2813_));
 sg13g2_a21oi_1 _6832_ (.A1(_2818_),
    .A2(_2819_),
    .Y(_2822_),
    .B1(net1009));
 sg13g2_a21oi_1 _6833_ (.A1(net1009),
    .A2(_2821_),
    .Y(_2823_),
    .B1(_2822_));
 sg13g2_mux2_1 _6834_ (.A0(_2823_),
    .A1(net388),
    .S(net972),
    .X(_0332_));
 sg13g2_xnor2_1 _6835_ (.Y(_2824_),
    .A(\vgademo.plane_u[4] ),
    .B(\vgademo.plane_du[4] ));
 sg13g2_a21oi_1 _6836_ (.A1(_2816_),
    .A2(_2819_),
    .Y(_2825_),
    .B1(_2824_));
 sg13g2_and3_1 _6837_ (.X(_2826_),
    .A(_2816_),
    .B(_2819_),
    .C(_2824_));
 sg13g2_o21ai_1 _6838_ (.B1(net1005),
    .Y(_2827_),
    .A1(_2825_),
    .A2(_2826_));
 sg13g2_nor2_1 _6839_ (.A(net1130),
    .B(_2820_),
    .Y(_2828_));
 sg13g2_xnor2_1 _6840_ (.Y(_2829_),
    .A(net1130),
    .B(_2820_));
 sg13g2_o21ai_1 _6841_ (.B1(_2827_),
    .Y(_2830_),
    .A1(net1005),
    .A2(_2829_));
 sg13g2_nand2_1 _6842_ (.Y(_2831_),
    .A(net289),
    .B(net972));
 sg13g2_o21ai_1 _6843_ (.B1(_2831_),
    .Y(_0333_),
    .A1(net972),
    .A2(_2830_));
 sg13g2_a21o_1 _6844_ (.A2(\vgademo.plane_du[4] ),
    .A1(\vgademo.plane_u[4] ),
    .B1(_2825_),
    .X(_2832_));
 sg13g2_xnor2_1 _6845_ (.Y(_2833_),
    .A(\vgademo.plane_u[5] ),
    .B(\vgademo.plane_du[5] ));
 sg13g2_xnor2_1 _6846_ (.Y(_2834_),
    .A(_2832_),
    .B(_2833_));
 sg13g2_nand2b_1 _6847_ (.Y(_2835_),
    .B(\vgademo.plane_dx[0] ),
    .A_N(_0023_));
 sg13g2_xnor2_1 _6848_ (.Y(_2836_),
    .A(\vgademo.plane_dx[0] ),
    .B(net1129));
 sg13g2_nand2_1 _6849_ (.Y(_2837_),
    .A(_0022_),
    .B(_2836_));
 sg13g2_xnor2_1 _6850_ (.Y(_2838_),
    .A(_0022_),
    .B(_2836_));
 sg13g2_xnor2_1 _6851_ (.Y(_2839_),
    .A(_2828_),
    .B(_2838_));
 sg13g2_a21oi_1 _6852_ (.A1(net1009),
    .A2(_2839_),
    .Y(_2840_),
    .B1(net972));
 sg13g2_o21ai_1 _6853_ (.B1(_2840_),
    .Y(_2841_),
    .A1(net1009),
    .A2(_2834_));
 sg13g2_o21ai_1 _6854_ (.B1(_2841_),
    .Y(_0334_),
    .A1(_3249_),
    .A2(_2799_));
 sg13g2_nand2_1 _6855_ (.Y(_2842_),
    .A(net297),
    .B(\vgademo.plane_du[6] ));
 sg13g2_xnor2_1 _6856_ (.Y(_2843_),
    .A(\vgademo.plane_u[6] ),
    .B(\vgademo.plane_du[6] ));
 sg13g2_a21oi_1 _6857_ (.A1(\vgademo.plane_u[5] ),
    .A2(\vgademo.plane_du[5] ),
    .Y(_2844_),
    .B1(_2832_));
 sg13g2_a21oi_2 _6858_ (.B1(_2844_),
    .Y(_2845_),
    .A2(_3250_),
    .A1(_3249_));
 sg13g2_nand2b_1 _6859_ (.Y(_2846_),
    .B(_2845_),
    .A_N(_2843_));
 sg13g2_xnor2_1 _6860_ (.Y(_2847_),
    .A(_2843_),
    .B(_2845_));
 sg13g2_o21ai_1 _6861_ (.B1(_2837_),
    .Y(_2848_),
    .A1(_2828_),
    .A2(_2838_));
 sg13g2_nand2_1 _6862_ (.Y(_2849_),
    .A(net1128),
    .B(\vgademo.plane_dx[1] ));
 sg13g2_xor2_1 _6863_ (.B(\vgademo.plane_dx[1] ),
    .A(net1127),
    .X(_2850_));
 sg13g2_nand2b_1 _6864_ (.Y(_2851_),
    .B(_2850_),
    .A_N(_2835_));
 sg13g2_xnor2_1 _6865_ (.Y(_2852_),
    .A(_2835_),
    .B(_2850_));
 sg13g2_xnor2_1 _6866_ (.Y(_2853_),
    .A(net1053),
    .B(_2852_));
 sg13g2_nor2b_1 _6867_ (.A(_2836_),
    .B_N(_2853_),
    .Y(_2854_));
 sg13g2_xnor2_1 _6868_ (.Y(_2855_),
    .A(_2836_),
    .B(_2853_));
 sg13g2_and2_1 _6869_ (.A(_2848_),
    .B(_2855_),
    .X(_2856_));
 sg13g2_o21ai_1 _6870_ (.B1(net1009),
    .Y(_2857_),
    .A1(_2848_),
    .A2(_2855_));
 sg13g2_o21ai_1 _6871_ (.B1(_2799_),
    .Y(_2858_),
    .A1(_2856_),
    .A2(_2857_));
 sg13g2_a21oi_1 _6872_ (.A1(net1004),
    .A2(_2847_),
    .Y(_2859_),
    .B1(_2858_));
 sg13g2_a21oi_1 _6873_ (.A1(_3252_),
    .A2(net973),
    .Y(_0335_),
    .B1(_2859_));
 sg13g2_nand2_1 _6874_ (.Y(_2860_),
    .A(net365),
    .B(\vgademo.plane_du[7] ));
 sg13g2_xnor2_1 _6875_ (.Y(_2861_),
    .A(\vgademo.plane_u[7] ),
    .B(\vgademo.plane_du[7] ));
 sg13g2_nand3_1 _6876_ (.B(_2846_),
    .C(_2861_),
    .A(_2842_),
    .Y(_2862_));
 sg13g2_a21o_1 _6877_ (.A2(_2846_),
    .A1(_2842_),
    .B1(_2861_),
    .X(_2863_));
 sg13g2_nand3_1 _6878_ (.B(_2862_),
    .C(_2863_),
    .A(net1003),
    .Y(_2864_));
 sg13g2_nor2_1 _6879_ (.A(_2854_),
    .B(_2856_),
    .Y(_2865_));
 sg13g2_nand2_1 _6880_ (.Y(_2866_),
    .A(\vgademo.plane_dx[0] ),
    .B(_2852_));
 sg13g2_xnor2_1 _6881_ (.Y(_2867_),
    .A(\vgademo.plane_dx_div.q[5] ),
    .B(\vgademo.plane_dx[2] ));
 sg13g2_a21oi_1 _6882_ (.A1(_2849_),
    .A2(_2851_),
    .Y(_2868_),
    .B1(_2867_));
 sg13g2_nand3_1 _6883_ (.B(_2851_),
    .C(_2867_),
    .A(_2849_),
    .Y(_2869_));
 sg13g2_nor2b_1 _6884_ (.A(_2868_),
    .B_N(_2869_),
    .Y(_2870_));
 sg13g2_xnor2_1 _6885_ (.Y(_2871_),
    .A(_0024_),
    .B(_2870_));
 sg13g2_nand2b_1 _6886_ (.Y(_2872_),
    .B(_2866_),
    .A_N(_2871_));
 sg13g2_xor2_1 _6887_ (.B(_2871_),
    .A(_2866_),
    .X(_2873_));
 sg13g2_xor2_1 _6888_ (.B(_2873_),
    .A(_2853_),
    .X(_2874_));
 sg13g2_nor2b_1 _6889_ (.A(_2874_),
    .B_N(_2865_),
    .Y(_2875_));
 sg13g2_nor2b_1 _6890_ (.A(_2865_),
    .B_N(_2874_),
    .Y(_2876_));
 sg13g2_inv_1 _6891_ (.Y(_2877_),
    .A(_2876_));
 sg13g2_nor3_1 _6892_ (.A(net1004),
    .B(_2875_),
    .C(_2876_),
    .Y(_2878_));
 sg13g2_nor2_1 _6893_ (.A(net971),
    .B(_2878_),
    .Y(_2879_));
 sg13g2_a22oi_1 _6894_ (.Y(_0336_),
    .B1(_2864_),
    .B2(_2879_),
    .A2(net971),
    .A1(_3253_));
 sg13g2_xnor2_1 _6895_ (.Y(_2880_),
    .A(\vgademo.plane_u[8] ),
    .B(\vgademo.plane_du[8] ));
 sg13g2_nand3_1 _6896_ (.B(_2863_),
    .C(_2880_),
    .A(_2860_),
    .Y(_2881_));
 sg13g2_a21o_1 _6897_ (.A2(_2863_),
    .A1(_2860_),
    .B1(_2880_),
    .X(_2882_));
 sg13g2_nand3_1 _6898_ (.B(_2881_),
    .C(_2882_),
    .A(net1003),
    .Y(_2883_));
 sg13g2_o21ai_1 _6899_ (.B1(_2877_),
    .Y(_2884_),
    .A1(_2853_),
    .A2(_2873_));
 sg13g2_nand2_1 _6900_ (.Y(_2885_),
    .A(\vgademo.plane_dx[1] ),
    .B(_2870_));
 sg13g2_a21oi_1 _6901_ (.A1(\vgademo.plane_dx_div.q[5] ),
    .A2(_3257_),
    .Y(_2886_),
    .B1(_2868_));
 sg13g2_xor2_1 _6902_ (.B(net1130),
    .A(net1125),
    .X(_2887_));
 sg13g2_nand2b_1 _6903_ (.Y(_2888_),
    .B(_2887_),
    .A_N(_2886_));
 sg13g2_xnor2_1 _6904_ (.Y(_2889_),
    .A(_2886_),
    .B(_2887_));
 sg13g2_xnor2_1 _6905_ (.Y(_2890_),
    .A(_0025_),
    .B(_2889_));
 sg13g2_nand2b_1 _6906_ (.Y(_2891_),
    .B(_2885_),
    .A_N(_2890_));
 sg13g2_xor2_1 _6907_ (.B(_2890_),
    .A(_2885_),
    .X(_2892_));
 sg13g2_xor2_1 _6908_ (.B(_2892_),
    .A(_2872_),
    .X(_2893_));
 sg13g2_nor2_1 _6909_ (.A(_2884_),
    .B(_2893_),
    .Y(_2894_));
 sg13g2_nand2_1 _6910_ (.Y(_2895_),
    .A(_2884_),
    .B(_2893_));
 sg13g2_nor2_1 _6911_ (.A(net1003),
    .B(_2894_),
    .Y(_2896_));
 sg13g2_a21oi_1 _6912_ (.A1(_2895_),
    .A2(_2896_),
    .Y(_2897_),
    .B1(net971));
 sg13g2_a22oi_1 _6913_ (.Y(_0337_),
    .B1(_2883_),
    .B2(_2897_),
    .A2(net970),
    .A1(_3255_));
 sg13g2_xnor2_1 _6914_ (.Y(_2898_),
    .A(\vgademo.plane_u[9] ),
    .B(\vgademo.plane_du[9] ));
 sg13g2_o21ai_1 _6915_ (.B1(_2882_),
    .Y(_2899_),
    .A1(_3255_),
    .A2(_3256_));
 sg13g2_xnor2_1 _6916_ (.Y(_2900_),
    .A(_2898_),
    .B(_2899_));
 sg13g2_o21ai_1 _6917_ (.B1(_2895_),
    .Y(_2901_),
    .A1(_2872_),
    .A2(_2892_));
 sg13g2_nand2_1 _6918_ (.Y(_2902_),
    .A(\vgademo.plane_dx[2] ),
    .B(_2889_));
 sg13g2_o21ai_1 _6919_ (.B1(_2888_),
    .Y(_2903_),
    .A1(_3164_),
    .A2(_0022_));
 sg13g2_nor2b_1 _6920_ (.A(net1129),
    .B_N(net1123),
    .Y(_2904_));
 sg13g2_xnor2_1 _6921_ (.Y(_2905_),
    .A(net1124),
    .B(net1129));
 sg13g2_xnor2_1 _6922_ (.Y(_2906_),
    .A(_2903_),
    .B(_2905_));
 sg13g2_nor2_1 _6923_ (.A(net1130),
    .B(_3172_),
    .Y(_2907_));
 sg13g2_xnor2_1 _6924_ (.Y(_2908_),
    .A(net1130),
    .B(net1053));
 sg13g2_xnor2_1 _6925_ (.Y(_2909_),
    .A(_2906_),
    .B(_2908_));
 sg13g2_nand2b_1 _6926_ (.Y(_2910_),
    .B(_2902_),
    .A_N(_2909_));
 sg13g2_xor2_1 _6927_ (.B(_2909_),
    .A(_2902_),
    .X(_2911_));
 sg13g2_xor2_1 _6928_ (.B(_2911_),
    .A(_2891_),
    .X(_2912_));
 sg13g2_nor2_1 _6929_ (.A(_2901_),
    .B(_2912_),
    .Y(_2913_));
 sg13g2_nand2_1 _6930_ (.Y(_2914_),
    .A(_2901_),
    .B(_2912_));
 sg13g2_nor2_1 _6931_ (.A(net1003),
    .B(_2913_),
    .Y(_2915_));
 sg13g2_a221oi_1 _6932_ (.B2(_2915_),
    .C1(net970),
    .B1(_2914_),
    .A1(net1003),
    .Y(_2916_),
    .A2(_2900_));
 sg13g2_a21oi_1 _6933_ (.A1(_3258_),
    .A2(net970),
    .Y(_0338_),
    .B1(_2916_));
 sg13g2_nand2_1 _6934_ (.Y(_2917_),
    .A(\vgademo.plane_u[10] ),
    .B(\vgademo.plane_du[10] ));
 sg13g2_xnor2_1 _6935_ (.Y(_2918_),
    .A(\vgademo.plane_u[10] ),
    .B(\vgademo.plane_du[10] ));
 sg13g2_o21ai_1 _6936_ (.B1(_2899_),
    .Y(_2919_),
    .A1(\vgademo.plane_u[9] ),
    .A2(\vgademo.plane_du[9] ));
 sg13g2_o21ai_1 _6937_ (.B1(_2919_),
    .Y(_2920_),
    .A1(_3258_),
    .A2(_3259_));
 sg13g2_nand2b_1 _6938_ (.Y(_2921_),
    .B(_2920_),
    .A_N(_2918_));
 sg13g2_xnor2_1 _6939_ (.Y(_2922_),
    .A(_2918_),
    .B(_2920_));
 sg13g2_o21ai_1 _6940_ (.B1(_2914_),
    .Y(_2923_),
    .A1(_2891_),
    .A2(_2911_));
 sg13g2_a21oi_2 _6941_ (.B1(_2907_),
    .Y(_2924_),
    .A2(_2908_),
    .A1(_2906_));
 sg13g2_xor2_1 _6942_ (.B(net1129),
    .A(\vgademo.plane_dx[1] ),
    .X(_2925_));
 sg13g2_a21oi_1 _6943_ (.A1(_2903_),
    .A2(_2905_),
    .Y(_2926_),
    .B1(_2904_));
 sg13g2_nand2_1 _6944_ (.Y(_2927_),
    .A(net1122),
    .B(net1127));
 sg13g2_nor2_1 _6945_ (.A(net1122),
    .B(net1127),
    .Y(_2928_));
 sg13g2_xor2_1 _6946_ (.B(net1127),
    .A(net1122),
    .X(_2929_));
 sg13g2_xnor2_1 _6947_ (.Y(_2930_),
    .A(_2926_),
    .B(_2929_));
 sg13g2_nor2_1 _6948_ (.A(_2925_),
    .B(_2930_),
    .Y(_2931_));
 sg13g2_xnor2_1 _6949_ (.Y(_2932_),
    .A(_2925_),
    .B(_2930_));
 sg13g2_nor2_1 _6950_ (.A(_2924_),
    .B(_2932_),
    .Y(_2933_));
 sg13g2_xor2_1 _6951_ (.B(_2932_),
    .A(_2924_),
    .X(_2934_));
 sg13g2_nor2b_1 _6952_ (.A(_2910_),
    .B_N(_2934_),
    .Y(_2935_));
 sg13g2_xnor2_1 _6953_ (.Y(_2936_),
    .A(_2910_),
    .B(_2934_));
 sg13g2_nor2_1 _6954_ (.A(_2923_),
    .B(_2936_),
    .Y(_2937_));
 sg13g2_nand2_1 _6955_ (.Y(_2938_),
    .A(_2923_),
    .B(_2936_));
 sg13g2_nor2_1 _6956_ (.A(net1003),
    .B(_2937_),
    .Y(_2939_));
 sg13g2_a221oi_1 _6957_ (.B2(_2939_),
    .C1(net970),
    .B1(_2938_),
    .A1(net1003),
    .Y(_2940_),
    .A2(_2922_));
 sg13g2_a21oi_1 _6958_ (.A1(_3260_),
    .A2(net970),
    .Y(_0339_),
    .B1(_2940_));
 sg13g2_a21oi_2 _6959_ (.B1(_0026_),
    .Y(_2941_),
    .A2(_2921_),
    .A1(_2917_));
 sg13g2_nand3_1 _6960_ (.B(_2917_),
    .C(_2921_),
    .A(_0026_),
    .Y(_2942_));
 sg13g2_nor2_1 _6961_ (.A(net1008),
    .B(_2941_),
    .Y(_2943_));
 sg13g2_nand2_1 _6962_ (.Y(_2944_),
    .A(_2942_),
    .B(_2943_));
 sg13g2_a21oi_1 _6963_ (.A1(_2923_),
    .A2(_2936_),
    .Y(_2945_),
    .B1(_2935_));
 sg13g2_a21oi_1 _6964_ (.A1(net1129),
    .A2(_0024_),
    .Y(_2946_),
    .B1(_2931_));
 sg13g2_xnor2_1 _6965_ (.Y(_2947_),
    .A(net1120),
    .B(net1126));
 sg13g2_o21ai_1 _6966_ (.B1(_2927_),
    .Y(_2948_),
    .A1(_2926_),
    .A2(_2928_));
 sg13g2_nor2b_1 _6967_ (.A(_2947_),
    .B_N(_2948_),
    .Y(_2949_));
 sg13g2_xor2_1 _6968_ (.B(_2948_),
    .A(_2947_),
    .X(_2950_));
 sg13g2_xor2_1 _6969_ (.B(\vgademo.plane_dx[2] ),
    .A(net1128),
    .X(_2951_));
 sg13g2_nand2_1 _6970_ (.Y(_2952_),
    .A(_2950_),
    .B(_2951_));
 sg13g2_xor2_1 _6971_ (.B(_2951_),
    .A(_2950_),
    .X(_2953_));
 sg13g2_nor2b_1 _6972_ (.A(_2946_),
    .B_N(_2953_),
    .Y(_2954_));
 sg13g2_xor2_1 _6973_ (.B(_2953_),
    .A(_2946_),
    .X(_2955_));
 sg13g2_or3_1 _6974_ (.A(_2924_),
    .B(_2932_),
    .C(_2955_),
    .X(_2956_));
 sg13g2_xor2_1 _6975_ (.B(_2955_),
    .A(_2933_),
    .X(_2957_));
 sg13g2_or2_1 _6976_ (.X(_2958_),
    .B(_2957_),
    .A(_2945_));
 sg13g2_a21oi_1 _6977_ (.A1(_2945_),
    .A2(_2957_),
    .Y(_2959_),
    .B1(net1003));
 sg13g2_a21oi_1 _6978_ (.A1(_2958_),
    .A2(_2959_),
    .Y(_2960_),
    .B1(net970));
 sg13g2_a22oi_1 _6979_ (.Y(_0340_),
    .B1(_2944_),
    .B2(_2960_),
    .A2(net970),
    .A1(_3261_));
 sg13g2_a21oi_1 _6980_ (.A1(_0027_),
    .A2(_2941_),
    .Y(_2961_),
    .B1(net1009));
 sg13g2_o21ai_1 _6981_ (.B1(_2961_),
    .Y(_2962_),
    .A1(_0027_),
    .A2(_2941_));
 sg13g2_nand2_1 _6982_ (.Y(_2963_),
    .A(_2956_),
    .B(_2958_));
 sg13g2_o21ai_1 _6983_ (.B1(_2952_),
    .Y(_2964_),
    .A1(net1128),
    .A2(_3257_));
 sg13g2_a21oi_1 _6984_ (.A1(net1120),
    .A2(net1126),
    .Y(_2965_),
    .B1(_2949_));
 sg13g2_nor2_1 _6985_ (.A(_3164_),
    .B(_2965_),
    .Y(_2966_));
 sg13g2_xnor2_1 _6986_ (.Y(_2967_),
    .A(net1125),
    .B(_2965_));
 sg13g2_xor2_1 _6987_ (.B(net1130),
    .A(net1126),
    .X(_2968_));
 sg13g2_nand2b_1 _6988_ (.Y(_2969_),
    .B(_2968_),
    .A_N(_2967_));
 sg13g2_xnor2_1 _6989_ (.Y(_2970_),
    .A(_2967_),
    .B(_2968_));
 sg13g2_nand2_1 _6990_ (.Y(_2971_),
    .A(_2964_),
    .B(_2970_));
 sg13g2_xnor2_1 _6991_ (.Y(_2972_),
    .A(_2964_),
    .B(_2970_));
 sg13g2_inv_1 _6992_ (.Y(_2973_),
    .A(_2972_));
 sg13g2_xor2_1 _6993_ (.B(_2972_),
    .A(_2954_),
    .X(_2974_));
 sg13g2_a21oi_1 _6994_ (.A1(_2956_),
    .A2(_2958_),
    .Y(_2975_),
    .B1(_2974_));
 sg13g2_xor2_1 _6995_ (.B(_2974_),
    .A(_2963_),
    .X(_2976_));
 sg13g2_a21oi_1 _6996_ (.A1(net1008),
    .A2(_2976_),
    .Y(_2977_),
    .B1(net971));
 sg13g2_a22oi_1 _6997_ (.Y(_2978_),
    .B1(_2962_),
    .B2(_2977_),
    .A2(net971),
    .A1(net378));
 sg13g2_inv_1 _6998_ (.Y(_0341_),
    .A(net379));
 sg13g2_a21oi_1 _6999_ (.A1(_2954_),
    .A2(_2973_),
    .Y(_2979_),
    .B1(_2975_));
 sg13g2_o21ai_1 _7000_ (.B1(_2969_),
    .Y(_2980_),
    .A1(net1126),
    .A2(_3251_));
 sg13g2_xnor2_1 _7001_ (.Y(_2981_),
    .A(net1124),
    .B(_2966_));
 sg13g2_nor2b_1 _7002_ (.A(net1125),
    .B_N(net1129),
    .Y(_2982_));
 sg13g2_xnor2_1 _7003_ (.Y(_2983_),
    .A(net1125),
    .B(net1129));
 sg13g2_xnor2_1 _7004_ (.Y(_2984_),
    .A(_2981_),
    .B(_2983_));
 sg13g2_nor2b_1 _7005_ (.A(_2984_),
    .B_N(_2980_),
    .Y(_2985_));
 sg13g2_xnor2_1 _7006_ (.Y(_2986_),
    .A(_2980_),
    .B(_2984_));
 sg13g2_nand2b_1 _7007_ (.Y(_2987_),
    .B(_2986_),
    .A_N(_2971_));
 sg13g2_xnor2_1 _7008_ (.Y(_2988_),
    .A(_2971_),
    .B(_2986_));
 sg13g2_nand2b_1 _7009_ (.Y(_2989_),
    .B(_2988_),
    .A_N(_2979_));
 sg13g2_nand2b_1 _7010_ (.Y(_2990_),
    .B(_2979_),
    .A_N(_2988_));
 sg13g2_nand3_1 _7011_ (.B(_2989_),
    .C(_2990_),
    .A(net1008),
    .Y(_2991_));
 sg13g2_and3_2 _7012_ (.X(_2992_),
    .A(\vgademo.plane_u[12] ),
    .B(\vgademo.plane_u[13] ),
    .C(_2941_));
 sg13g2_a21oi_1 _7013_ (.A1(net378),
    .A2(_2941_),
    .Y(_2993_),
    .B1(net482));
 sg13g2_nor3_1 _7014_ (.A(net1008),
    .B(_2992_),
    .C(_2993_),
    .Y(_2994_));
 sg13g2_nor2_1 _7015_ (.A(net971),
    .B(_2994_),
    .Y(_2995_));
 sg13g2_a22oi_1 _7016_ (.Y(_0342_),
    .B1(_2991_),
    .B2(_2995_),
    .A2(net971),
    .A1(_3262_));
 sg13g2_a21oi_1 _7017_ (.A1(_2981_),
    .A2(_2983_),
    .Y(_2996_),
    .B1(_2982_));
 sg13g2_nand3_1 _7018_ (.B(net1124),
    .C(_2966_),
    .A(net1122),
    .Y(_2997_));
 sg13g2_a21o_1 _7019_ (.A2(_2966_),
    .A1(net1124),
    .B1(net1122),
    .X(_2998_));
 sg13g2_nand2_1 _7020_ (.Y(_2999_),
    .A(_2997_),
    .B(_2998_));
 sg13g2_xor2_1 _7021_ (.B(net1127),
    .A(net1123),
    .X(_3000_));
 sg13g2_nand2_1 _7022_ (.Y(_3001_),
    .A(_2999_),
    .B(_3000_));
 sg13g2_xnor2_1 _7023_ (.Y(_3002_),
    .A(_2999_),
    .B(_3000_));
 sg13g2_nor2_1 _7024_ (.A(_2996_),
    .B(_3002_),
    .Y(_3003_));
 sg13g2_xor2_1 _7025_ (.B(_3002_),
    .A(_2996_),
    .X(_3004_));
 sg13g2_and2_1 _7026_ (.A(_2985_),
    .B(_3004_),
    .X(_3005_));
 sg13g2_xnor2_1 _7027_ (.Y(_3006_),
    .A(_2985_),
    .B(_3004_));
 sg13g2_a21oi_1 _7028_ (.A1(_2987_),
    .A2(_2989_),
    .Y(_3007_),
    .B1(_3006_));
 sg13g2_and3_1 _7029_ (.X(_3008_),
    .A(_2987_),
    .B(_2989_),
    .C(_3006_));
 sg13g2_o21ai_1 _7030_ (.B1(net1008),
    .Y(_3009_),
    .A1(_3007_),
    .A2(_3008_));
 sg13g2_xnor2_1 _7031_ (.Y(_3010_),
    .A(\vgademo.plane_u[14] ),
    .B(_2992_));
 sg13g2_a21oi_1 _7032_ (.A1(net1005),
    .A2(_3010_),
    .Y(_3011_),
    .B1(net969));
 sg13g2_a22oi_1 _7033_ (.Y(_3012_),
    .B1(_3009_),
    .B2(_3011_),
    .A2(net969),
    .A1(net463));
 sg13g2_inv_1 _7034_ (.Y(_0343_),
    .A(net464));
 sg13g2_nor2b_1 _7035_ (.A(_0028_),
    .B_N(_2992_),
    .Y(_3013_));
 sg13g2_xnor2_1 _7036_ (.Y(_3014_),
    .A(_3263_),
    .B(_3013_));
 sg13g2_a21oi_1 _7037_ (.A1(net1001),
    .A2(_3014_),
    .Y(_3015_),
    .B1(net969));
 sg13g2_o21ai_1 _7038_ (.B1(_3001_),
    .Y(_3016_),
    .A1(net1123),
    .A2(net1127));
 sg13g2_or2_1 _7039_ (.X(_3017_),
    .B(net1126),
    .A(net1121));
 sg13g2_xnor2_1 _7040_ (.Y(_3018_),
    .A(net1121),
    .B(net1126));
 sg13g2_xor2_1 _7041_ (.B(_2997_),
    .A(net1119),
    .X(_3019_));
 sg13g2_nand2b_1 _7042_ (.Y(_3020_),
    .B(_3019_),
    .A_N(_3018_));
 sg13g2_xnor2_1 _7043_ (.Y(_3021_),
    .A(_3018_),
    .B(_3019_));
 sg13g2_nand2_1 _7044_ (.Y(_3022_),
    .A(_3016_),
    .B(_3021_));
 sg13g2_xor2_1 _7045_ (.B(_3021_),
    .A(_3016_),
    .X(_3023_));
 sg13g2_nand2_1 _7046_ (.Y(_3024_),
    .A(_3003_),
    .B(_3023_));
 sg13g2_xor2_1 _7047_ (.B(_3023_),
    .A(_3003_),
    .X(_3025_));
 sg13g2_o21ai_1 _7048_ (.B1(_3025_),
    .Y(_3026_),
    .A1(_3005_),
    .A2(_3007_));
 sg13g2_or3_1 _7049_ (.A(_3005_),
    .B(_3007_),
    .C(_3025_),
    .X(_3027_));
 sg13g2_nand3_1 _7050_ (.B(_3026_),
    .C(_3027_),
    .A(net1008),
    .Y(_3028_));
 sg13g2_a22oi_1 _7051_ (.Y(_0344_),
    .B1(_3015_),
    .B2(_3028_),
    .A2(net969),
    .A1(_3263_));
 sg13g2_a21oi_1 _7052_ (.A1(net1119),
    .A2(_2997_),
    .Y(_3029_),
    .B1(_3164_));
 sg13g2_a21o_1 _7053_ (.A2(_3164_),
    .A1(net1119),
    .B1(_3029_),
    .X(_3030_));
 sg13g2_a21oi_2 _7054_ (.B1(_3030_),
    .Y(_3031_),
    .A2(_3020_),
    .A1(_3017_));
 sg13g2_nand3_1 _7055_ (.B(_3020_),
    .C(_3030_),
    .A(_3017_),
    .Y(_3032_));
 sg13g2_nand2b_1 _7056_ (.Y(_3033_),
    .B(_3032_),
    .A_N(_3031_));
 sg13g2_or2_1 _7057_ (.X(_3034_),
    .B(_3033_),
    .A(_3022_));
 sg13g2_xnor2_1 _7058_ (.Y(_3035_),
    .A(_3022_),
    .B(_3033_));
 sg13g2_a21o_1 _7059_ (.A2(_3026_),
    .A1(_3024_),
    .B1(_3035_),
    .X(_3036_));
 sg13g2_nand3_1 _7060_ (.B(_3026_),
    .C(_3035_),
    .A(_3024_),
    .Y(_3037_));
 sg13g2_and3_1 _7061_ (.X(_3038_),
    .A(\vgademo.plane_u[14] ),
    .B(\vgademo.plane_u[15] ),
    .C(_2992_));
 sg13g2_a21o_1 _7062_ (.A2(_3037_),
    .A1(_3036_),
    .B1(net1005),
    .X(_3039_));
 sg13g2_xor2_1 _7063_ (.B(_3038_),
    .A(_0029_),
    .X(_3040_));
 sg13g2_a21oi_1 _7064_ (.A1(net1002),
    .A2(_3040_),
    .Y(_3041_),
    .B1(net968));
 sg13g2_a22oi_1 _7065_ (.Y(_3042_),
    .B1(_3039_),
    .B2(_3041_),
    .A2(net968),
    .A1(net418));
 sg13g2_inv_1 _7066_ (.Y(_0345_),
    .A(net419));
 sg13g2_a21oi_2 _7067_ (.B1(net1123),
    .Y(_3043_),
    .A2(net1125),
    .A1(net1120));
 sg13g2_nand3_1 _7068_ (.B(net1123),
    .C(net1125),
    .A(net1119),
    .Y(_3044_));
 sg13g2_nor2b_1 _7069_ (.A(_3043_),
    .B_N(_3044_),
    .Y(_3045_));
 sg13g2_xnor2_1 _7070_ (.Y(_3046_),
    .A(_3031_),
    .B(_3045_));
 sg13g2_a21oi_1 _7071_ (.A1(_3034_),
    .A2(_3036_),
    .Y(_3047_),
    .B1(_3046_));
 sg13g2_nand3_1 _7072_ (.B(_3036_),
    .C(_3046_),
    .A(_3034_),
    .Y(_3048_));
 sg13g2_nand2b_1 _7073_ (.Y(_3049_),
    .B(_3048_),
    .A_N(_3047_));
 sg13g2_nand3_1 _7074_ (.B(\vgademo.plane_u[17] ),
    .C(_3038_),
    .A(\vgademo.plane_u[16] ),
    .Y(_3050_));
 sg13g2_a21o_1 _7075_ (.A2(_3038_),
    .A1(\vgademo.plane_u[16] ),
    .B1(\vgademo.plane_u[17] ),
    .X(_3051_));
 sg13g2_a21oi_1 _7076_ (.A1(_3050_),
    .A2(_3051_),
    .Y(_3052_),
    .B1(net1010));
 sg13g2_a21oi_1 _7077_ (.A1(net1010),
    .A2(_3049_),
    .Y(_3053_),
    .B1(_3052_));
 sg13g2_mux2_1 _7078_ (.A0(net475),
    .A1(_3053_),
    .S(_2799_),
    .X(_0346_));
 sg13g2_a21oi_1 _7079_ (.A1(_3031_),
    .A2(_3045_),
    .Y(_3054_),
    .B1(_3047_));
 sg13g2_xnor2_1 _7080_ (.Y(_3055_),
    .A(net1121),
    .B(_3043_));
 sg13g2_nor2_1 _7081_ (.A(_3054_),
    .B(_3055_),
    .Y(_3056_));
 sg13g2_a21oi_1 _7082_ (.A1(_3054_),
    .A2(_3055_),
    .Y(_3057_),
    .B1(net1002));
 sg13g2_nand2b_1 _7083_ (.Y(_3058_),
    .B(_3057_),
    .A_N(_3056_));
 sg13g2_xnor2_1 _7084_ (.Y(_3059_),
    .A(net508),
    .B(_3050_));
 sg13g2_a21oi_1 _7085_ (.A1(net1001),
    .A2(_3059_),
    .Y(_3060_),
    .B1(net968));
 sg13g2_a22oi_1 _7086_ (.Y(_0347_),
    .B1(_3058_),
    .B2(_3060_),
    .A2(net968),
    .A1(_3264_));
 sg13g2_a21oi_1 _7087_ (.A1(net1121),
    .A2(_3043_),
    .Y(_3061_),
    .B1(_3056_));
 sg13g2_nor2_1 _7088_ (.A(net1119),
    .B(net1121),
    .Y(_3062_));
 sg13g2_xnor2_1 _7089_ (.Y(_3063_),
    .A(net1119),
    .B(net1121));
 sg13g2_xnor2_1 _7090_ (.Y(_3064_),
    .A(_3061_),
    .B(_3063_));
 sg13g2_nor2_1 _7091_ (.A(_0030_),
    .B(_3050_),
    .Y(_3065_));
 sg13g2_xnor2_1 _7092_ (.Y(_3066_),
    .A(net414),
    .B(_3065_));
 sg13g2_a21oi_1 _7093_ (.A1(net1001),
    .A2(_3066_),
    .Y(_3067_),
    .B1(net968));
 sg13g2_o21ai_1 _7094_ (.B1(_3067_),
    .Y(_3068_),
    .A1(net1001),
    .A2(_3064_));
 sg13g2_o21ai_1 _7095_ (.B1(_3068_),
    .Y(_0348_),
    .A1(_3265_),
    .A2(_2799_));
 sg13g2_or3_1 _7096_ (.A(_3264_),
    .B(_3265_),
    .C(_3050_),
    .X(_3069_));
 sg13g2_xnor2_1 _7097_ (.Y(_3070_),
    .A(net266),
    .B(_3069_));
 sg13g2_nand3_1 _7098_ (.B(net1121),
    .C(_3061_),
    .A(net1119),
    .Y(_3071_));
 sg13g2_a21oi_1 _7099_ (.A1(_3056_),
    .A2(_3062_),
    .Y(_3072_),
    .B1(net1001));
 sg13g2_a21o_1 _7100_ (.A2(_3062_),
    .A1(_3056_),
    .B1(net1001),
    .X(_3073_));
 sg13g2_a221oi_1 _7101_ (.B2(_3072_),
    .C1(net969),
    .B1(_3071_),
    .A1(net1001),
    .Y(_3074_),
    .A2(_3070_));
 sg13g2_a21oi_1 _7102_ (.A1(_3266_),
    .A2(net968),
    .Y(_0349_),
    .B1(_3074_));
 sg13g2_nor2_1 _7103_ (.A(_0031_),
    .B(_3069_),
    .Y(_3075_));
 sg13g2_xnor2_1 _7104_ (.Y(_3076_),
    .A(_3267_),
    .B(_3075_));
 sg13g2_a21oi_1 _7105_ (.A1(net1001),
    .A2(_3076_),
    .Y(_3077_),
    .B1(net968));
 sg13g2_a22oi_1 _7106_ (.Y(_0350_),
    .B1(_3073_),
    .B2(_3077_),
    .A2(net968),
    .A1(_3267_));
 sg13g2_o21ai_1 _7107_ (.B1(_1914_),
    .Y(_3078_),
    .A1(_1858_),
    .A2(_1880_));
 sg13g2_nand2_1 _7108_ (.Y(_3079_),
    .A(net955),
    .B(_3078_));
 sg13g2_o21ai_1 _7109_ (.B1(_2196_),
    .Y(_3080_),
    .A1(_1824_),
    .A2(_3079_));
 sg13g2_a21oi_2 _7110_ (.B1(_2238_),
    .Y(_3081_),
    .A2(_3080_),
    .A1(net898));
 sg13g2_nor2_1 _7111_ (.A(_1317_),
    .B(_3081_),
    .Y(_3082_));
 sg13g2_a22oi_1 _7112_ (.Y(_3083_),
    .B1(net905),
    .B2(_2222_),
    .A2(_1912_),
    .A1(_1857_));
 sg13g2_o21ai_1 _7113_ (.B1(net955),
    .Y(_3084_),
    .A1(_1824_),
    .A2(_3083_));
 sg13g2_nand3_1 _7114_ (.B(_2205_),
    .C(_2211_),
    .A(_2204_),
    .Y(_3085_));
 sg13g2_a221oi_1 _7115_ (.B2(_2666_),
    .C1(net963),
    .B1(_3085_),
    .A1(_2664_),
    .Y(_3086_),
    .A2(_3084_));
 sg13g2_nor2_1 _7116_ (.A(_1317_),
    .B(_3086_),
    .Y(_3087_));
 sg13g2_o21ai_1 _7117_ (.B1(_2228_),
    .Y(_3088_),
    .A1(_1317_),
    .A2(_3086_));
 sg13g2_nand2_1 _7118_ (.Y(_3089_),
    .A(_3082_),
    .B(_3088_));
 sg13g2_or3_1 _7119_ (.A(_1317_),
    .B(_2228_),
    .C(_3086_),
    .X(_3090_));
 sg13g2_nand2b_1 _7120_ (.Y(_3091_),
    .B(_3090_),
    .A_N(_3082_));
 sg13g2_and2_1 _7121_ (.A(_3089_),
    .B(_3091_),
    .X(_3092_));
 sg13g2_xnor2_1 _7122_ (.Y(_3093_),
    .A(_1838_),
    .B(_1851_));
 sg13g2_a22oi_1 _7123_ (.Y(_3094_),
    .B1(_3093_),
    .B2(_2243_),
    .A2(_2248_),
    .A1(net905));
 sg13g2_nor4_1 _7124_ (.A(net902),
    .B(net899),
    .C(net947),
    .D(_3078_),
    .Y(_3095_));
 sg13g2_a221oi_1 _7125_ (.B2(_3094_),
    .C1(_3095_),
    .B1(net896),
    .A1(net957),
    .Y(_3096_),
    .A2(net960));
 sg13g2_nand2_1 _7126_ (.Y(_3097_),
    .A(net898),
    .B(_2253_));
 sg13g2_o21ai_1 _7127_ (.B1(_2692_),
    .Y(_3098_),
    .A1(_3096_),
    .A2(_3097_));
 sg13g2_nand2_1 _7128_ (.Y(_3099_),
    .A(net961),
    .B(_3098_));
 sg13g2_a21oi_1 _7129_ (.A1(net961),
    .A2(_3098_),
    .Y(_3100_),
    .B1(net1040));
 sg13g2_a21o_1 _7130_ (.A2(_3098_),
    .A1(net961),
    .B1(net1040),
    .X(_3101_));
 sg13g2_nand3_1 _7131_ (.B(net1040),
    .C(_3098_),
    .A(net961),
    .Y(_3102_));
 sg13g2_and3_1 _7132_ (.X(_3103_),
    .A(_3087_),
    .B(_3101_),
    .C(_3102_));
 sg13g2_a21oi_1 _7133_ (.A1(_3087_),
    .A2(_3102_),
    .Y(_3104_),
    .B1(_3100_));
 sg13g2_a21oi_1 _7134_ (.A1(_3088_),
    .A2(_3090_),
    .Y(_3105_),
    .B1(_3082_));
 sg13g2_and3_1 _7135_ (.X(_3106_),
    .A(_3082_),
    .B(_3088_),
    .C(_3090_));
 sg13g2_nor3_1 _7136_ (.A(_3104_),
    .B(_3105_),
    .C(_3106_),
    .Y(_3107_));
 sg13g2_o21ai_1 _7137_ (.B1(_3104_),
    .Y(_3108_),
    .A1(_3105_),
    .A2(_3106_));
 sg13g2_xor2_1 _7138_ (.B(\vgademo.plane_u[14] ),
    .A(\vgademo.a_cos[9] ),
    .X(_3109_));
 sg13g2_xnor2_1 _7139_ (.Y(_3110_),
    .A(_1849_),
    .B(_3109_));
 sg13g2_o21ai_1 _7140_ (.B1(_2271_),
    .Y(_3111_),
    .A1(_2244_),
    .A2(_3110_));
 sg13g2_inv_1 _7141_ (.Y(_3112_),
    .A(_3111_));
 sg13g2_nor4_1 _7142_ (.A(net902),
    .B(net899),
    .C(net947),
    .D(_3083_),
    .Y(_3113_));
 sg13g2_a221oi_1 _7143_ (.B2(_3111_),
    .C1(_3113_),
    .B1(net897),
    .A1(net957),
    .Y(_3114_),
    .A2(net960));
 sg13g2_o21ai_1 _7144_ (.B1(_2215_),
    .Y(_3115_),
    .A1(_2301_),
    .A2(_3114_));
 sg13g2_nand2_1 _7145_ (.Y(_3116_),
    .A(_1318_),
    .B(_3115_));
 sg13g2_and3_1 _7146_ (.X(_3117_),
    .A(_1318_),
    .B(_2307_),
    .C(_3115_));
 sg13g2_nand3_1 _7147_ (.B(_2307_),
    .C(_3115_),
    .A(_1318_),
    .Y(_3118_));
 sg13g2_a21o_1 _7148_ (.A2(_3115_),
    .A1(_1318_),
    .B1(_2307_),
    .X(_3119_));
 sg13g2_and3_1 _7149_ (.X(_3120_),
    .A(_3099_),
    .B(_3118_),
    .C(_3119_));
 sg13g2_a21oi_1 _7150_ (.A1(_3099_),
    .A2(_3119_),
    .Y(_3121_),
    .B1(_3117_));
 sg13g2_a21oi_1 _7151_ (.A1(_3101_),
    .A2(_3102_),
    .Y(_3122_),
    .B1(_3087_));
 sg13g2_o21ai_1 _7152_ (.B1(_3121_),
    .Y(_3123_),
    .A1(_3103_),
    .A2(_3122_));
 sg13g2_xnor2_1 _7153_ (.Y(_3124_),
    .A(_1841_),
    .B(_1845_));
 sg13g2_o21ai_1 _7154_ (.B1(_2267_),
    .Y(_3125_),
    .A1(_2244_),
    .A2(_3124_));
 sg13g2_nor4_1 _7155_ (.A(net904),
    .B(net901),
    .C(net948),
    .D(_3112_),
    .Y(_3126_));
 sg13g2_a221oi_1 _7156_ (.B2(_3125_),
    .C1(_3126_),
    .B1(net897),
    .A1(net957),
    .Y(_3127_),
    .A2(net960));
 sg13g2_o21ai_1 _7157_ (.B1(net962),
    .Y(_3128_),
    .A1(_2278_),
    .A2(_3127_));
 sg13g2_and2_1 _7158_ (.A(_2266_),
    .B(_3128_),
    .X(_3129_));
 sg13g2_xnor2_1 _7159_ (.Y(_3130_),
    .A(_1846_),
    .B(_1848_));
 sg13g2_nand2_1 _7160_ (.Y(_3131_),
    .A(_2243_),
    .B(_3130_));
 sg13g2_and2_1 _7161_ (.A(_2290_),
    .B(_3131_),
    .X(_3132_));
 sg13g2_mux2_1 _7162_ (.A0(_3094_),
    .A1(_3132_),
    .S(net896),
    .X(_3133_));
 sg13g2_a21oi_1 _7163_ (.A1(net955),
    .A2(_3133_),
    .Y(_3134_),
    .B1(_2285_));
 sg13g2_or2_1 _7164_ (.X(_3135_),
    .B(_3134_),
    .A(net963));
 sg13g2_xor2_1 _7165_ (.B(_3128_),
    .A(_2266_),
    .X(_3136_));
 sg13g2_a21oi_1 _7166_ (.A1(_3135_),
    .A2(_3136_),
    .Y(_3137_),
    .B1(_3129_));
 sg13g2_a21oi_1 _7167_ (.A1(_3118_),
    .A2(_3119_),
    .Y(_3138_),
    .B1(_3099_));
 sg13g2_o21ai_1 _7168_ (.B1(_3137_),
    .Y(_3139_),
    .A1(_3120_),
    .A2(_3138_));
 sg13g2_o21ai_1 _7169_ (.B1(_2313_),
    .Y(_3140_),
    .A1(_1317_),
    .A2(_3081_));
 sg13g2_nor2_1 _7170_ (.A(_2313_),
    .B(_3081_),
    .Y(_3141_));
 sg13g2_o21ai_1 _7171_ (.B1(_3140_),
    .Y(_3142_),
    .A1(_3135_),
    .A2(_3141_));
 sg13g2_nand2_1 _7172_ (.Y(_3143_),
    .A(_3116_),
    .B(_3142_));
 sg13g2_xnor2_1 _7173_ (.Y(_3144_),
    .A(_3135_),
    .B(_3136_));
 sg13g2_o21ai_1 _7174_ (.B1(_3144_),
    .Y(_3145_),
    .A1(_3116_),
    .A2(_3142_));
 sg13g2_nand3_1 _7175_ (.B(_3143_),
    .C(_3145_),
    .A(_3139_),
    .Y(_3146_));
 sg13g2_nor3_1 _7176_ (.A(_3103_),
    .B(_3121_),
    .C(_3122_),
    .Y(_3147_));
 sg13g2_nor3_1 _7177_ (.A(_3120_),
    .B(_3137_),
    .C(_3138_),
    .Y(_3148_));
 sg13g2_a21oi_1 _7178_ (.A1(_3108_),
    .A2(_3123_),
    .Y(_3149_),
    .B1(_3107_));
 sg13g2_nor3_1 _7179_ (.A(_3107_),
    .B(_3147_),
    .C(_3148_),
    .Y(_3150_));
 sg13g2_a21oi_1 _7180_ (.A1(_3146_),
    .A2(_3150_),
    .Y(_3151_),
    .B1(_3149_));
 sg13g2_nand2_1 _7181_ (.Y(_3152_),
    .A(_3092_),
    .B(_3151_));
 sg13g2_o21ai_1 _7182_ (.B1(_2335_),
    .Y(_3153_),
    .A1(_3092_),
    .A2(_3151_));
 sg13g2_nor2b_1 _7183_ (.A(_3153_),
    .B_N(_3152_),
    .Y(_0351_));
 sg13g2_a21oi_1 _7184_ (.A1(_3089_),
    .A2(_3152_),
    .Y(_0352_),
    .B1(_2336_));
 sg13g2_nor2_1 _7185_ (.A(net287),
    .B(net990),
    .Y(_3154_));
 sg13g2_a21oi_1 _7186_ (.A1(_3166_),
    .A2(net990),
    .Y(_0353_),
    .B1(_3154_));
 sg13g2_nor2_1 _7187_ (.A(net305),
    .B(net990),
    .Y(_3155_));
 sg13g2_a21oi_1 _7188_ (.A1(_3165_),
    .A2(net990),
    .Y(_0354_),
    .B1(_3155_));
 sg13g2_mux2_1 _7189_ (.A0(net435),
    .A1(\vgademo.plane_dx[2] ),
    .S(net990),
    .X(_0355_));
 sg13g2_nand2_1 _7190_ (.Y(_3156_),
    .A(net1130),
    .B(net991));
 sg13g2_o21ai_1 _7191_ (.B1(_3156_),
    .Y(_0356_),
    .A1(_3247_),
    .A2(net989));
 sg13g2_nor2_1 _7192_ (.A(\vgademo.plane_du[4] ),
    .B(net989),
    .Y(_3157_));
 sg13g2_a21oi_1 _7193_ (.A1(net1129),
    .A2(net991),
    .Y(_0357_),
    .B1(_3157_));
 sg13g2_nand2_1 _7194_ (.Y(_3158_),
    .A(net1127),
    .B(net989));
 sg13g2_o21ai_1 _7195_ (.B1(_3158_),
    .Y(_0358_),
    .A1(_3250_),
    .A2(net989));
 sg13g2_mux2_1 _7196_ (.A0(net578),
    .A1(net1126),
    .S(net989),
    .X(_0359_));
 sg13g2_nor2_1 _7197_ (.A(\vgademo.plane_du[7] ),
    .B(net989),
    .Y(_3159_));
 sg13g2_a21oi_1 _7198_ (.A1(_3164_),
    .A2(net989),
    .Y(_0360_),
    .B1(_3159_));
 sg13g2_mux2_1 _7199_ (.A0(net579),
    .A1(net1123),
    .S(net989),
    .X(_0361_));
 sg13g2_nand2_1 _7200_ (.Y(_3160_),
    .A(net1122),
    .B(net990));
 sg13g2_o21ai_1 _7201_ (.B1(_3160_),
    .Y(_0362_),
    .A1(_3259_),
    .A2(net990));
 sg13g2_mux2_1 _7202_ (.A0(net534),
    .A1(net1120),
    .S(net990),
    .X(_0363_));
 sg13g2_a21oi_1 _7203_ (.A1(\vgademo.plane_du[0] ),
    .A2(_2799_),
    .Y(_3161_),
    .B1(net233));
 sg13g2_a21oi_1 _7204_ (.A1(net1004),
    .A2(_2800_),
    .Y(_3162_),
    .B1(net972));
 sg13g2_nor2_1 _7205_ (.A(net234),
    .B(_3162_),
    .Y(_0364_));
 sg13g2_dfrbp_1 _7206_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net37),
    .D(_0111_),
    .Q_N(_3632_),
    .Q(\vgademo.linelfsr[0] ));
 sg13g2_dfrbp_1 _7207_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net119),
    .D(_0112_),
    .Q_N(_3631_),
    .Q(\vgademo.linelfsr[1] ));
 sg13g2_dfrbp_1 _7208_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net117),
    .D(net371),
    .Q_N(_3630_),
    .Q(\vgademo.linelfsr[2] ));
 sg13g2_dfrbp_1 _7209_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net115),
    .D(_0114_),
    .Q_N(_3629_),
    .Q(\vgademo.linelfsr[3] ));
 sg13g2_dfrbp_1 _7210_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net113),
    .D(_0115_),
    .Q_N(_3628_),
    .Q(\vgademo.linelfsr[4] ));
 sg13g2_dfrbp_1 _7211_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net111),
    .D(_0116_),
    .Q_N(_3627_),
    .Q(\vgademo.linelfsr[5] ));
 sg13g2_dfrbp_1 _7212_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net109),
    .D(net320),
    .Q_N(_3626_),
    .Q(\vgademo.linelfsr[6] ));
 sg13g2_dfrbp_1 _7213_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net107),
    .D(net369),
    .Q_N(_3625_),
    .Q(\vgademo.linelfsr[7] ));
 sg13g2_dfrbp_1 _7214_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net105),
    .D(net377),
    .Q_N(_3624_),
    .Q(\vgademo.linelfsr[8] ));
 sg13g2_dfrbp_1 _7215_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net103),
    .D(net404),
    .Q_N(_3623_),
    .Q(\vgademo.linelfsr[9] ));
 sg13g2_dfrbp_1 _7216_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net101),
    .D(net402),
    .Q_N(_3622_),
    .Q(\vgademo.linelfsr[10] ));
 sg13g2_dfrbp_1 _7217_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net99),
    .D(_0122_),
    .Q_N(_3621_),
    .Q(\vgademo.linelfsr[11] ));
 sg13g2_dfrbp_1 _7218_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net97),
    .D(_0123_),
    .Q_N(_3620_),
    .Q(\vgademo.linelfsr[12] ));
 sg13g2_dfrbp_1 _7219_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1158),
    .D(net272),
    .Q_N(\vgademo.audio_songpos[0] ),
    .Q(_0085_));
 sg13g2_dfrbp_1 _7220_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1158),
    .D(_0125_),
    .Q_N(\vgademo.audio_songpos[1] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _7221_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1159),
    .D(_0126_),
    .Q_N(\vgademo.audio_songpos[2] ),
    .Q(_0087_));
 sg13g2_dfrbp_1 _7222_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1158),
    .D(_0127_),
    .Q_N(\vgademo.audio_songpos[3] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 _7223_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1159),
    .D(_0128_),
    .Q_N(\vgademo.audio_songpos[4] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _7224_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1159),
    .D(_0129_),
    .Q_N(\vgademo.audio_songpos[5] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _7225_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1159),
    .D(_0130_),
    .Q_N(\vgademo.audio_songpos[6] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _7226_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1159),
    .D(net190),
    .Q_N(\vgademo.audio_songpos[7] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 _7227_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net76),
    .D(_0132_),
    .Q_N(_0024_),
    .Q(\vgademo.plane_dx[1] ));
 sg13g2_dfrbp_1 _7228_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net74),
    .D(_0133_),
    .Q_N(_0025_),
    .Q(\vgademo.plane_dx[2] ));
 sg13g2_dfrbp_1 _7229_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net72),
    .D(_0134_),
    .Q_N(_0022_),
    .Q(\vgademo.plane_dx[3] ));
 sg13g2_dfrbp_1 _7230_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net70),
    .D(_0135_),
    .Q_N(_0023_),
    .Q(\vgademo.plane_dx_div.q[3] ));
 sg13g2_dfrbp_1 _7231_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net68),
    .D(_0136_),
    .Q_N(_3619_),
    .Q(\vgademo.plane_dx_div.q[4] ));
 sg13g2_dfrbp_1 _7232_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net66),
    .D(_0137_),
    .Q_N(_3618_),
    .Q(\vgademo.plane_dx_div.q[5] ));
 sg13g2_dfrbp_1 _7233_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net64),
    .D(_0138_),
    .Q_N(_3617_),
    .Q(\vgademo.plane_dx_div.q[6] ));
 sg13g2_dfrbp_1 _7234_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net62),
    .D(_0139_),
    .Q_N(_3616_),
    .Q(\vgademo.plane_dx_div.q[7] ));
 sg13g2_dfrbp_1 _7235_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net60),
    .D(_0140_),
    .Q_N(_3615_),
    .Q(\vgademo.plane_dx_div.q[8] ));
 sg13g2_dfrbp_1 _7236_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net58),
    .D(_0141_),
    .Q_N(_3614_),
    .Q(\vgademo.plane_dx_div.q[9] ));
 sg13g2_dfrbp_1 _7237_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0142_),
    .Q_N(_0084_),
    .Q(\vgademo.plane_dx_div.i[0] ));
 sg13g2_dfrbp_1 _7238_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net54),
    .D(net329),
    .Q_N(_3613_),
    .Q(\vgademo.plane_dx_div.i[1] ));
 sg13g2_dfrbp_1 _7239_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net52),
    .D(_0144_),
    .Q_N(_3612_),
    .Q(\vgademo.plane_dx_div.i[2] ));
 sg13g2_dfrbp_1 _7240_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net38),
    .D(_0145_),
    .Q_N(_3633_),
    .Q(\vgademo.plane_dx_div.i[3] ));
 sg13g2_dfrbp_1 _7241_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1161),
    .D(\vgademo.soundtrack.sigma_delta_accum_[0] ),
    .Q_N(_3634_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[0] ));
 sg13g2_dfrbp_1 _7242_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1161),
    .D(\vgademo.soundtrack.sigma_delta_accum_[1] ),
    .Q_N(_3635_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[1] ));
 sg13g2_dfrbp_1 _7243_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1161),
    .D(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .Q_N(_3636_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[2] ));
 sg13g2_dfrbp_1 _7244_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1161),
    .D(net528),
    .Q_N(_3637_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[3] ));
 sg13g2_dfrbp_1 _7245_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1171),
    .D(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .Q_N(_3638_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[4] ));
 sg13g2_dfrbp_1 _7246_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1171),
    .D(\vgademo.soundtrack.sigma_delta_accum_[5] ),
    .Q_N(_3639_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[5] ));
 sg13g2_dfrbp_1 _7247_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1171),
    .D(net521),
    .Q_N(_3640_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[6] ));
 sg13g2_dfrbp_1 _7248_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1171),
    .D(net500),
    .Q_N(_3641_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[7] ));
 sg13g2_dfrbp_1 _7249_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1171),
    .D(\vgademo.soundtrack.sigma_delta_accum_[8] ),
    .Q_N(_3642_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[8] ));
 sg13g2_dfrbp_1 _7250_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1172),
    .D(net526),
    .Q_N(_3643_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[9] ));
 sg13g2_dfrbp_1 _7251_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1172),
    .D(net511),
    .Q_N(_3644_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[10] ));
 sg13g2_dfrbp_1 _7252_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1172),
    .D(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .Q_N(_3645_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[11] ));
 sg13g2_dfrbp_1 _7253_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1163),
    .D(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .Q_N(_3646_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[12] ));
 sg13g2_dfrbp_1 _7254_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1163),
    .D(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .Q_N(_3647_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[13] ));
 sg13g2_dfrbp_1 _7255_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1164),
    .D(\vgademo.soundtrack.sigma_delta_accum_[14] ),
    .Q_N(_3648_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[14] ));
 sg13g2_dfrbp_1 _7256_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1164),
    .D(\vgademo.soundtrack.sigma_delta_accum_[15] ),
    .Q_N(_3611_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[15] ));
 sg13g2_dfrbp_1 _7257_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1163),
    .D(_0146_),
    .Q_N(_0057_),
    .Q(\vgademo.audio_beat_out[0] ));
 sg13g2_dfrbp_1 _7258_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1163),
    .D(_0147_),
    .Q_N(_0058_),
    .Q(\vgademo.audio_beat_out[1] ));
 sg13g2_dfrbp_1 _7259_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1162),
    .D(_0148_),
    .Q_N(_0061_),
    .Q(\vgademo.audio_beat_out[2] ));
 sg13g2_dfrbp_1 _7260_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1163),
    .D(net408),
    .Q_N(_0056_),
    .Q(\vgademo.audio_beat_out[3] ));
 sg13g2_dfrbp_1 _7261_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1162),
    .D(_0150_),
    .Q_N(_0054_),
    .Q(\vgademo.audio_beat_out[4] ));
 sg13g2_dfrbp_1 _7262_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1158),
    .D(_0151_),
    .Q_N(_3610_),
    .Q(\vgademo.soundtrack.tri_osc_i[0] ));
 sg13g2_dfrbp_1 _7263_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1158),
    .D(_0152_),
    .Q_N(_3609_),
    .Q(\vgademo.soundtrack.tri_osc_i[1] ));
 sg13g2_dfrbp_1 _7264_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1158),
    .D(_0153_),
    .Q_N(_3608_),
    .Q(\vgademo.soundtrack.tri_osc_i[2] ));
 sg13g2_dfrbp_1 _7265_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1158),
    .D(net517),
    .Q_N(_3607_),
    .Q(\vgademo.soundtrack.tri_osc_i[3] ));
 sg13g2_dfrbp_1 _7266_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1158),
    .D(_0155_),
    .Q_N(_3606_),
    .Q(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_dfrbp_1 _7267_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1160),
    .D(_0156_),
    .Q_N(_3605_),
    .Q(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_dfrbp_1 _7268_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1160),
    .D(_0157_),
    .Q_N(_3604_),
    .Q(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_dfrbp_1 _7269_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1160),
    .D(_0158_),
    .Q_N(_3603_),
    .Q(\vgademo.soundtrack.tri_osc_i[7] ));
 sg13g2_dfrbp_1 _7270_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1160),
    .D(_0159_),
    .Q_N(_3602_),
    .Q(\vgademo.soundtrack.tri_osc_i[8] ));
 sg13g2_dfrbp_1 _7271_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net49),
    .D(net249),
    .Q_N(_3601_),
    .Q(audio));
 sg13g2_dfrbp_1 _7272_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1176),
    .D(net176),
    .Q_N(\vgademo.soundtrack.tick_div_[0] ),
    .Q(\vgademo.soundtrack.tick_div[0] ));
 sg13g2_dfrbp_1 _7273_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1176),
    .D(net491),
    .Q_N(_3600_),
    .Q(\vgademo.soundtrack.tick_div[1] ));
 sg13g2_dfrbp_1 _7274_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1176),
    .D(net243),
    .Q_N(_3599_),
    .Q(\vgademo.soundtrack.tick_div[2] ));
 sg13g2_dfrbp_1 _7275_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1176),
    .D(net253),
    .Q_N(_3598_),
    .Q(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_dfrbp_1 _7276_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1179),
    .D(net227),
    .Q_N(_3597_),
    .Q(\vgademo.soundtrack.tick_div[4] ));
 sg13g2_dfrbp_1 _7277_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1173),
    .D(net265),
    .Q_N(_3596_),
    .Q(\vgademo.soundtrack.tick_div[5] ));
 sg13g2_dfrbp_1 _7278_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1174),
    .D(net201),
    .Q_N(_3595_),
    .Q(\vgademo.soundtrack.tick_div[6] ));
 sg13g2_dfrbp_1 _7279_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1173),
    .D(net221),
    .Q_N(_3594_),
    .Q(\vgademo.soundtrack.tick_div[7] ));
 sg13g2_dfrbp_1 _7280_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1169),
    .D(net170),
    .Q_N(\vgademo.soundtrack.noise_lfsr[0] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 _7281_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1169),
    .D(net188),
    .Q_N(\vgademo.soundtrack.noise_lfsr[1] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 _7282_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1169),
    .D(net194),
    .Q_N(\vgademo.soundtrack.noise_lfsr[2] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 _7283_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1169),
    .D(net223),
    .Q_N(\vgademo.soundtrack.noise_lfsr[3] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 _7284_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1169),
    .D(net241),
    .Q_N(_0039_),
    .Q(\vgademo.soundtrack.noise_lfsr[4] ));
 sg13g2_dfrbp_1 _7285_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1173),
    .D(net174),
    .Q_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 _7286_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1173),
    .D(net261),
    .Q_N(_0083_),
    .Q(\vgademo.soundtrack.noise_lfsr[6] ));
 sg13g2_dfrbp_1 _7287_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1172),
    .D(net178),
    .Q_N(\vgademo.soundtrack.noise_lfsr[7] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 _7288_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1172),
    .D(net331),
    .Q_N(_0082_),
    .Q(\vgademo.soundtrack.noise_lfsr[8] ));
 sg13g2_dfrbp_1 _7289_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1170),
    .D(net205),
    .Q_N(_3593_),
    .Q(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_dfrbp_1 _7290_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1169),
    .D(net168),
    .Q_N(\vgademo.soundtrack.noise_lfsr[10] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 _7291_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1169),
    .D(net198),
    .Q_N(\vgademo.soundtrack.noise_lfsr[11] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _7292_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1170),
    .D(net172),
    .Q_N(\vgademo.soundtrack.noise_lfsr[12] ),
    .Q(_0101_));
 sg13g2_dfrbp_1 _7293_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1170),
    .D(net245),
    .Q_N(_0081_),
    .Q(\vgademo.soundtrack.noise_lfsr[13] ));
 sg13g2_dfrbp_1 _7294_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1169),
    .D(net293),
    .Q_N(_3592_),
    .Q(\vgademo.soundtrack.noise_lfsr[14] ));
 sg13g2_dfrbp_1 _7295_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1162),
    .D(net184),
    .Q_N(\vgademo.audio_snare_frames[0] ),
    .Q(_0102_));
 sg13g2_dfrbp_1 _7296_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1162),
    .D(net182),
    .Q_N(\vgademo.audio_snare_frames[1] ),
    .Q(_0103_));
 sg13g2_dfrbp_1 _7297_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1162),
    .D(net212),
    .Q_N(\vgademo.audio_snare_frames[2] ),
    .Q(_0104_));
 sg13g2_dfrbp_1 _7298_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1162),
    .D(net180),
    .Q_N(\vgademo.audio_snare_frames[3] ),
    .Q(_0105_));
 sg13g2_dfrbp_1 _7299_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net20),
    .D(_0188_),
    .Q_N(_3591_),
    .Q(\vgademo.soundtrack.pulse_osc_p[0] ));
 sg13g2_dfrbp_1 _7300_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net19),
    .D(net219),
    .Q_N(_0041_),
    .Q(\vgademo.soundtrack.pulse_osc_p[1] ));
 sg13g2_dfrbp_1 _7301_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net18),
    .D(net362),
    .Q_N(_3590_),
    .Q(\vgademo.soundtrack.pulse_osc_p[2] ));
 sg13g2_dfrbp_1 _7302_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net17),
    .D(_0191_),
    .Q_N(_3589_),
    .Q(\vgademo.soundtrack.pulse_osc_p[3] ));
 sg13g2_dfrbp_1 _7303_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net16),
    .D(net317),
    .Q_N(_3588_),
    .Q(\vgademo.soundtrack.pulse_osc_p[4] ));
 sg13g2_dfrbp_1 _7304_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net15),
    .D(_0193_),
    .Q_N(_3587_),
    .Q(\vgademo.soundtrack.pulse_osc_p[5] ));
 sg13g2_dfrbp_1 _7305_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net163),
    .D(net346),
    .Q_N(_3586_),
    .Q(\vgademo.soundtrack.pulse_osc_p[6] ));
 sg13g2_dfrbp_1 _7306_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net162),
    .D(_0195_),
    .Q_N(_3585_),
    .Q(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_dfrbp_1 _7307_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net161),
    .D(net268),
    .Q_N(_3584_),
    .Q(\vgademo.soundtrack.pulse_osc_p[8] ));
 sg13g2_dfrbp_1 _7308_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net160),
    .D(net232),
    .Q_N(_3583_),
    .Q(\vgademo.soundtrack.pulse_osc_p[9] ));
 sg13g2_dfrbp_1 _7309_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net159),
    .D(net210),
    .Q_N(_3582_),
    .Q(\vgademo.soundtrack.pulse_osc_p[10] ));
 sg13g2_dfrbp_1 _7310_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net158),
    .D(_0199_),
    .Q_N(_3581_),
    .Q(\vgademo.soundtrack.pulse_osc_p[11] ));
 sg13g2_dfrbp_1 _7311_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net157),
    .D(_0200_),
    .Q_N(_3580_),
    .Q(\vgademo.soundtrack.pulse_osc_p[12] ));
 sg13g2_dfrbp_1 _7312_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net156),
    .D(net239),
    .Q_N(_3579_),
    .Q(\vgademo.soundtrack.pulse_osc_p[13] ));
 sg13g2_dfrbp_1 _7313_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1160),
    .D(_0202_),
    .Q_N(_3578_),
    .Q(\vgademo.audio_kick_frames[0] ));
 sg13g2_dfrbp_1 _7314_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1162),
    .D(_0203_),
    .Q_N(_0067_),
    .Q(\vgademo.audio_kick_frames[1] ));
 sg13g2_dfrbp_1 _7315_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1160),
    .D(net281),
    .Q_N(_0059_),
    .Q(\vgademo.audio_kick_frames[2] ));
 sg13g2_dfrbp_1 _7316_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1161),
    .D(_0205_),
    .Q_N(\vgademo.soundtrack.pulse_vol[0] ),
    .Q(_0106_));
 sg13g2_dfrbp_1 _7317_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1161),
    .D(_0206_),
    .Q_N(\vgademo.soundtrack.pulse_vol[1] ),
    .Q(_0107_));
 sg13g2_dfrbp_1 _7318_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1161),
    .D(_0207_),
    .Q_N(\vgademo.soundtrack.pulse_vol[2] ),
    .Q(_0108_));
 sg13g2_dfrbp_1 _7319_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1164),
    .D(net203),
    .Q_N(\vgademo.soundtrack.pulse_vol[3] ),
    .Q(_0109_));
 sg13g2_dfrbp_1 _7320_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1177),
    .D(net165),
    .Q_N(\vgademo.soundtrack.sample_div_[0] ),
    .Q(\vgademo.soundtrack.sample_div[0] ));
 sg13g2_dfrbp_1 _7321_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1177),
    .D(net259),
    .Q_N(_3649_),
    .Q(\vgademo.soundtrack.sample_div[1] ));
 sg13g2_dfrbp_1 _7322_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1176),
    .D(net467),
    .Q_N(_3650_),
    .Q(\vgademo.soundtrack.sample_div[2] ));
 sg13g2_dfrbp_1 _7323_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1176),
    .D(net255),
    .Q_N(_3651_),
    .Q(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_dfrbp_1 _7324_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1176),
    .D(net216),
    .Q_N(_3652_),
    .Q(\vgademo.soundtrack.sample_div[4] ));
 sg13g2_dfrbp_1 _7325_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1176),
    .D(\vgademo.soundtrack.sample_div_[5] ),
    .Q_N(_3653_),
    .Q(\vgademo.soundtrack.sample_div[5] ));
 sg13g2_dfrbp_1 _7326_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1177),
    .D(\vgademo.soundtrack.sample_div_[6] ),
    .Q_N(_3654_),
    .Q(\vgademo.soundtrack.sample_div[6] ));
 sg13g2_dfrbp_1 _7327_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1177),
    .D(net229),
    .Q_N(_3655_),
    .Q(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_dfrbp_1 _7328_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1177),
    .D(net225),
    .Q_N(_3656_),
    .Q(\vgademo.soundtrack.sample_div[8] ));
 sg13g2_dfrbp_1 _7329_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net1170),
    .D(\vgademo.soundtrack.sample_div_[9] ),
    .Q_N(_3577_),
    .Q(\vgademo.soundtrack.sample_div[9] ));
 sg13g2_dfrbp_1 _7330_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net147),
    .D(net247),
    .Q_N(_3576_),
    .Q(\vgademo.soundtrack.tri_osc_p[0] ));
 sg13g2_dfrbp_1 _7331_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net146),
    .D(_0210_),
    .Q_N(_3575_),
    .Q(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_dfrbp_1 _7332_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net145),
    .D(_0211_),
    .Q_N(_3574_),
    .Q(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_dfrbp_1 _7333_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net144),
    .D(net432),
    .Q_N(_3573_),
    .Q(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_dfrbp_1 _7334_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net143),
    .D(_0213_),
    .Q_N(_3572_),
    .Q(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_dfrbp_1 _7335_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net142),
    .D(net434),
    .Q_N(_3571_),
    .Q(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_dfrbp_1 _7336_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net141),
    .D(_0215_),
    .Q_N(_3570_),
    .Q(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_dfrbp_1 _7337_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net140),
    .D(_0216_),
    .Q_N(_3569_),
    .Q(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_dfrbp_1 _7338_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net139),
    .D(_0217_),
    .Q_N(_3568_),
    .Q(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_dfrbp_1 _7339_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net138),
    .D(net337),
    .Q_N(_0040_),
    .Q(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_dfrbp_1 _7340_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net137),
    .D(net310),
    .Q_N(_3567_),
    .Q(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_dfrbp_1 _7341_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net136),
    .D(net295),
    .Q_N(_3566_),
    .Q(\vgademo.soundtrack.tri_osc_p[11] ));
 sg13g2_dfrbp_1 _7342_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net135),
    .D(_0221_),
    .Q_N(_3565_),
    .Q(\vgademo.soundtrack.tri_osc_p[12] ));
 sg13g2_dfrbp_1 _7343_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net134),
    .D(_0222_),
    .Q_N(_3564_),
    .Q(\vgademo.soundtrack.tri_osc_p[13] ));
 sg13g2_dfrbp_1 _7344_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net133),
    .D(net367),
    .Q_N(_3563_),
    .Q(\vgademo.soundtrack.tri_osc_p[14] ));
 sg13g2_dfrbp_1 _7345_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net132),
    .D(net400),
    .Q_N(_3562_),
    .Q(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_dfrbp_1 _7346_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net131),
    .D(_0225_),
    .Q_N(_3561_),
    .Q(\vgademo.plane_dx_div.d[16] ));
 sg13g2_dfrbp_1 _7347_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net130),
    .D(_0226_),
    .Q_N(_0069_),
    .Q(\vgademo.plane_dx_div.d[17] ));
 sg13g2_dfrbp_1 _7348_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net129),
    .D(_0227_),
    .Q_N(_0072_),
    .Q(\vgademo.plane_dx_div.d[18] ));
 sg13g2_dfrbp_1 _7349_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net128),
    .D(_0228_),
    .Q_N(_0075_),
    .Q(\vgademo.plane_dx_div.d[19] ));
 sg13g2_dfrbp_1 _7350_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net127),
    .D(_0229_),
    .Q_N(_0078_),
    .Q(\vgademo.plane_dx_div.d[20] ));
 sg13g2_dfrbp_1 _7351_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net126),
    .D(_0230_),
    .Q_N(_0080_),
    .Q(\vgademo.plane_dx_div.d[21] ));
 sg13g2_dfrbp_1 _7352_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net125),
    .D(_0231_),
    .Q_N(_0013_),
    .Q(\vgademo.plane_dx_div.d[22] ));
 sg13g2_dfrbp_1 _7353_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net124),
    .D(_0232_),
    .Q_N(_0017_),
    .Q(\vgademo.plane_dx_div.d[23] ));
 sg13g2_dfrbp_1 _7354_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net91),
    .D(_0233_),
    .Q_N(_0020_),
    .Q(\vgademo.plane_dx_div.d[24] ));
 sg13g2_dfrbp_1 _7355_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net92),
    .D(_0012_),
    .Q_N(_3657_),
    .Q(\vgademo.vsync ));
 sg13g2_dfrbp_1 _7356_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net93),
    .D(_0011_),
    .Q_N(_3658_),
    .Q(hsync));
 sg13g2_dfrbp_1 _7357_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1181),
    .D(_0000_),
    .Q_N(_3659_),
    .Q(\vgademo.h_count[0] ));
 sg13g2_dfrbp_1 _7358_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1175),
    .D(_0002_),
    .Q_N(_3660_),
    .Q(\vgademo.h_count[1] ));
 sg13g2_dfrbp_1 _7359_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1172),
    .D(_0003_),
    .Q_N(_0032_),
    .Q(\vgademo.h_count[2] ));
 sg13g2_dfrbp_1 _7360_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1181),
    .D(_0004_),
    .Q_N(_0033_),
    .Q(\vgademo.h_count[3] ));
 sg13g2_dfrbp_1 _7361_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1163),
    .D(_0005_),
    .Q_N(_0043_),
    .Q(\vgademo.h_count[4] ));
 sg13g2_dfrbp_1 _7362_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1163),
    .D(net301),
    .Q_N(_0034_),
    .Q(\vgademo.h_count[5] ));
 sg13g2_dfrbp_1 _7363_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1168),
    .D(_0007_),
    .Q_N(_0035_),
    .Q(\vgademo.h_count[6] ));
 sg13g2_dfrbp_1 _7364_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1168),
    .D(net560),
    .Q_N(_0036_),
    .Q(\vgademo.h_count[7] ));
 sg13g2_dfrbp_1 _7365_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1167),
    .D(_0009_),
    .Q_N(_0037_),
    .Q(\vgademo.h_count[8] ));
 sg13g2_dfrbp_1 _7366_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1167),
    .D(net387),
    .Q_N(_0038_),
    .Q(\vgademo.h_count[9] ));
 sg13g2_dfrbp_1 _7367_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1167),
    .D(_0001_),
    .Q_N(_0060_),
    .Q(\vgademo.h_count[10] ));
 sg13g2_dfrbp_1 _7368_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1165),
    .D(_0234_),
    .Q_N(_0063_),
    .Q(\vgademo.a_scrolly[3] ));
 sg13g2_dfrbp_1 _7369_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1165),
    .D(_0235_),
    .Q_N(_0068_),
    .Q(\vgademo.a_scrolly[4] ));
 sg13g2_dfrbp_1 _7370_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1165),
    .D(_0236_),
    .Q_N(_0055_),
    .Q(\vgademo.a_scrolly[5] ));
 sg13g2_dfrbp_1 _7371_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1165),
    .D(net581),
    .Q_N(_0074_),
    .Q(\vgademo.a_scrolly[6] ));
 sg13g2_dfrbp_1 _7372_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1166),
    .D(net547),
    .Q_N(_0077_),
    .Q(\vgademo.a_scrolly[7] ));
 sg13g2_dfrbp_1 _7373_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1165),
    .D(_0239_),
    .Q_N(_0079_),
    .Q(\vgademo.a_scrolly[8] ));
 sg13g2_dfrbp_1 _7374_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1166),
    .D(_0240_),
    .Q_N(_0064_),
    .Q(\vgademo.a_scrolly[9] ));
 sg13g2_dfrbp_1 _7375_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1166),
    .D(_0241_),
    .Q_N(_0015_),
    .Q(\vgademo.a_scrolly[10] ));
 sg13g2_dfrbp_1 _7376_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1165),
    .D(net572),
    .Q_N(_0019_),
    .Q(\vgademo.a_scrolly[11] ));
 sg13g2_dfrbp_1 _7377_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1165),
    .D(net557),
    .Q_N(_0066_),
    .Q(\vgademo.a_scrolly[12] ));
 sg13g2_dfrbp_1 _7378_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net1165),
    .D(net555),
    .Q_N(_0065_),
    .Q(\vgademo.a_scrolly[13] ));
 sg13g2_dfrbp_1 _7379_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1181),
    .D(_0245_),
    .Q_N(_3560_),
    .Q(\vgademo.bayer_j[0] ));
 sg13g2_dfrbp_1 _7380_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1181),
    .D(_0246_),
    .Q_N(_0071_),
    .Q(\vgademo.bayer_j[1] ));
 sg13g2_dfrbp_1 _7381_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1182),
    .D(net257),
    .Q_N(_0070_),
    .Q(\vgademo.v_count[2] ));
 sg13g2_dfrbp_1 _7382_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1182),
    .D(net457),
    .Q_N(_0073_),
    .Q(\vgademo.v_count[3] ));
 sg13g2_dfrbp_1 _7383_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1181),
    .D(net488),
    .Q_N(_0076_),
    .Q(\vgademo.v_count[4] ));
 sg13g2_dfrbp_1 _7384_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1181),
    .D(net504),
    .Q_N(_0062_),
    .Q(\vgademo.v_count[5] ));
 sg13g2_dfrbp_1 _7385_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1181),
    .D(net566),
    .Q_N(_0016_),
    .Q(\vgademo.v_count[6] ));
 sg13g2_dfrbp_1 _7386_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1167),
    .D(_0252_),
    .Q_N(_0014_),
    .Q(\vgademo.v_count[7] ));
 sg13g2_dfrbp_1 _7387_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1167),
    .D(net453),
    .Q_N(_0018_),
    .Q(\vgademo.v_count[8] ));
 sg13g2_dfrbp_1 _7388_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1167),
    .D(net341),
    .Q_N(_0021_),
    .Q(\vgademo.v_count[9] ));
 sg13g2_dfrbp_1 _7389_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net123),
    .D(_0255_),
    .Q_N(_3559_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7390_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net122),
    .D(_0256_),
    .Q_N(_3558_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7391_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1179),
    .D(net251),
    .Q_N(_3557_),
    .Q(\vgademo.a_cos[0] ));
 sg13g2_dfrbp_1 _7392_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1179),
    .D(net314),
    .Q_N(_3556_),
    .Q(\vgademo.a_cos[1] ));
 sg13g2_dfrbp_1 _7393_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1178),
    .D(_0259_),
    .Q_N(_3555_),
    .Q(\vgademo.a_cos[2] ));
 sg13g2_dfrbp_1 _7394_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1178),
    .D(_0260_),
    .Q_N(_3554_),
    .Q(\vgademo.a_cos[3] ));
 sg13g2_dfrbp_1 _7395_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1178),
    .D(_0261_),
    .Q_N(_3553_),
    .Q(\vgademo.a_cos[4] ));
 sg13g2_dfrbp_1 _7396_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1183),
    .D(_0262_),
    .Q_N(_3552_),
    .Q(\vgademo.a_cos[5] ));
 sg13g2_dfrbp_1 _7397_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1183),
    .D(_0263_),
    .Q_N(_3551_),
    .Q(\vgademo.a_cos[6] ));
 sg13g2_dfrbp_1 _7398_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1183),
    .D(_0264_),
    .Q_N(_3550_),
    .Q(\vgademo.a_cos[7] ));
 sg13g2_dfrbp_1 _7399_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1179),
    .D(_0265_),
    .Q_N(_3549_),
    .Q(\vgademo.a_cos[8] ));
 sg13g2_dfrbp_1 _7400_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1179),
    .D(_0266_),
    .Q_N(_3548_),
    .Q(\vgademo.a_cos[9] ));
 sg13g2_dfrbp_1 _7401_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1174),
    .D(_0267_),
    .Q_N(_3547_),
    .Q(\vgademo.a_cos[10] ));
 sg13g2_dfrbp_1 _7402_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1174),
    .D(_0268_),
    .Q_N(_3546_),
    .Q(\vgademo.a_cos[11] ));
 sg13g2_dfrbp_1 _7403_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1174),
    .D(_0269_),
    .Q_N(_3545_),
    .Q(\vgademo.a_cos[12] ));
 sg13g2_dfrbp_1 _7404_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1172),
    .D(_0270_),
    .Q_N(\vgademo.a_cos[13] ),
    .Q(_0110_));
 sg13g2_dfrbp_1 _7405_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1172),
    .D(_0271_),
    .Q_N(_3544_),
    .Q(\vgademo.a_cos[14] ));
 sg13g2_dfrbp_1 _7406_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1183),
    .D(_0272_),
    .Q_N(_3543_),
    .Q(\vgademo.a_sin[0] ));
 sg13g2_dfrbp_1 _7407_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1183),
    .D(net348),
    .Q_N(_3542_),
    .Q(\vgademo.a_sin[1] ));
 sg13g2_dfrbp_1 _7408_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1179),
    .D(_0274_),
    .Q_N(_3541_),
    .Q(\vgademo.a_sin[2] ));
 sg13g2_dfrbp_1 _7409_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1179),
    .D(_0275_),
    .Q_N(_3540_),
    .Q(\vgademo.a_sin[3] ));
 sg13g2_dfrbp_1 _7410_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1174),
    .D(net356),
    .Q_N(_3539_),
    .Q(\vgademo.a_sin[4] ));
 sg13g2_dfrbp_1 _7411_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1173),
    .D(_0277_),
    .Q_N(_3538_),
    .Q(\vgademo.a_sin[5] ));
 sg13g2_dfrbp_1 _7412_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1173),
    .D(_0278_),
    .Q_N(_3537_),
    .Q(\vgademo.a_sin[6] ));
 sg13g2_dfrbp_1 _7413_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1173),
    .D(_0279_),
    .Q_N(_3536_),
    .Q(\vgademo.a_sin[7] ));
 sg13g2_dfrbp_1 _7414_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1173),
    .D(_0280_),
    .Q_N(_3535_),
    .Q(\vgademo.a_sin[8] ));
 sg13g2_dfrbp_1 _7415_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1178),
    .D(_0281_),
    .Q_N(_3534_),
    .Q(\vgademo.a_sin[9] ));
 sg13g2_dfrbp_1 _7416_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1178),
    .D(_0282_),
    .Q_N(_3533_),
    .Q(\vgademo.a_sin[10] ));
 sg13g2_dfrbp_1 _7417_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1178),
    .D(_0283_),
    .Q_N(_3532_),
    .Q(\vgademo.a_sin[11] ));
 sg13g2_dfrbp_1 _7418_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1178),
    .D(_0284_),
    .Q_N(_3531_),
    .Q(\vgademo.a_sin[12] ));
 sg13g2_dfrbp_1 _7419_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1178),
    .D(_0285_),
    .Q_N(_3530_),
    .Q(\vgademo.a_sin[13] ));
 sg13g2_dfrbp_1 _7420_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1180),
    .D(_0286_),
    .Q_N(_3529_),
    .Q(\vgademo.a_sin[14] ));
 sg13g2_dfrbp_1 _7421_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net120),
    .D(_0287_),
    .Q_N(_3528_),
    .Q(\vgademo.scanline_audio_sample[0] ));
 sg13g2_dfrbp_1 _7422_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net118),
    .D(_0288_),
    .Q_N(_3527_),
    .Q(\vgademo.scanline_audio_sample[1] ));
 sg13g2_dfrbp_1 _7423_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net116),
    .D(_0289_),
    .Q_N(_3526_),
    .Q(\vgademo.scanline_audio_sample[2] ));
 sg13g2_dfrbp_1 _7424_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net114),
    .D(_0290_),
    .Q_N(_3525_),
    .Q(\vgademo.scanline_audio_sample[3] ));
 sg13g2_dfrbp_1 _7425_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net112),
    .D(_0291_),
    .Q_N(_3524_),
    .Q(\vgademo.scanline_audio_sample[4] ));
 sg13g2_dfrbp_1 _7426_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net110),
    .D(_0292_),
    .Q_N(_0042_),
    .Q(\vgademo.scanline_audio_sample[5] ));
 sg13g2_dfrbp_1 _7427_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net108),
    .D(_0293_),
    .Q_N(_3523_),
    .Q(\vgademo.scanline_audio_sample[6] ));
 sg13g2_dfrbp_1 _7428_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net106),
    .D(net326),
    .Q_N(_3522_),
    .Q(\vgademo.b_cos[0] ));
 sg13g2_dfrbp_1 _7429_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net104),
    .D(_0295_),
    .Q_N(_3521_),
    .Q(\vgademo.b_cos[1] ));
 sg13g2_dfrbp_1 _7430_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net102),
    .D(net450),
    .Q_N(_3520_),
    .Q(\vgademo.b_cos[2] ));
 sg13g2_dfrbp_1 _7431_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net100),
    .D(net358),
    .Q_N(_3519_),
    .Q(\vgademo.b_cos[3] ));
 sg13g2_dfrbp_1 _7432_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net98),
    .D(net393),
    .Q_N(_3518_),
    .Q(\vgademo.b_cos[4] ));
 sg13g2_dfrbp_1 _7433_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net96),
    .D(_0299_),
    .Q_N(_3517_),
    .Q(\vgademo.b_cos[5] ));
 sg13g2_dfrbp_1 _7434_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net95),
    .D(_0300_),
    .Q_N(_3516_),
    .Q(\vgademo.b_cos[6] ));
 sg13g2_dfrbp_1 _7435_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net94),
    .D(net462),
    .Q_N(_3515_),
    .Q(\vgademo.b_cos[7] ));
 sg13g2_dfrbp_1 _7436_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net90),
    .D(net440),
    .Q_N(_3514_),
    .Q(\vgademo.b_cos[8] ));
 sg13g2_dfrbp_1 _7437_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net89),
    .D(net438),
    .Q_N(_3513_),
    .Q(\vgademo.b_cos[9] ));
 sg13g2_dfrbp_1 _7438_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net88),
    .D(_0304_),
    .Q_N(_3512_),
    .Q(\vgademo.b_cos[10] ));
 sg13g2_dfrbp_1 _7439_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net87),
    .D(net423),
    .Q_N(_3511_),
    .Q(\vgademo.b_cos[11] ));
 sg13g2_dfrbp_1 _7440_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net86),
    .D(net335),
    .Q_N(_3510_),
    .Q(\vgademo.plane_dx_div.r[16] ));
 sg13g2_dfrbp_1 _7441_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net85),
    .D(net360),
    .Q_N(_3509_),
    .Q(\vgademo.plane_dx_div.r[17] ));
 sg13g2_dfrbp_1 _7442_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net84),
    .D(net339),
    .Q_N(_3508_),
    .Q(\vgademo.plane_dx_div.r[18] ));
 sg13g2_dfrbp_1 _7443_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net83),
    .D(_0309_),
    .Q_N(_3507_),
    .Q(\vgademo.plane_dx_div.r[19] ));
 sg13g2_dfrbp_1 _7444_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net82),
    .D(net263),
    .Q_N(_3506_),
    .Q(\vgademo.plane_dx_div.r[20] ));
 sg13g2_dfrbp_1 _7445_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net81),
    .D(_0311_),
    .Q_N(_3505_),
    .Q(\vgademo.plane_dx_div.r[21] ));
 sg13g2_dfrbp_1 _7446_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net80),
    .D(net384),
    .Q_N(_3504_),
    .Q(\vgademo.plane_dx_div.r[22] ));
 sg13g2_dfrbp_1 _7447_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net79),
    .D(_0313_),
    .Q_N(_3503_),
    .Q(\vgademo.plane_dx_div.r[23] ));
 sg13g2_dfrbp_1 _7448_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net78),
    .D(_0314_),
    .Q_N(_3502_),
    .Q(\vgademo.plane_dx_div.r[24] ));
 sg13g2_dfrbp_1 _7449_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net77),
    .D(_0315_),
    .Q_N(\vgademo.plane_dx[0] ),
    .Q(\vgademo.plane_dx_div.r[25] ));
 sg13g2_dfrbp_1 _7450_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net75),
    .D(_0316_),
    .Q_N(_3501_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7451_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net73),
    .D(_0317_),
    .Q_N(_3500_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7452_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net71),
    .D(_0318_),
    .Q_N(_3499_),
    .Q(\vgademo.b_sin[0] ));
 sg13g2_dfrbp_1 _7453_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net69),
    .D(net364),
    .Q_N(_3498_),
    .Q(\vgademo.b_sin[1] ));
 sg13g2_dfrbp_1 _7454_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net67),
    .D(_0320_),
    .Q_N(_3497_),
    .Q(\vgademo.b_sin[2] ));
 sg13g2_dfrbp_1 _7455_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net65),
    .D(_0321_),
    .Q_N(_3496_),
    .Q(\vgademo.b_sin[3] ));
 sg13g2_dfrbp_1 _7456_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net63),
    .D(_0322_),
    .Q_N(_3495_),
    .Q(\vgademo.b_sin[4] ));
 sg13g2_dfrbp_1 _7457_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net61),
    .D(_0323_),
    .Q_N(_3494_),
    .Q(\vgademo.b_sin[5] ));
 sg13g2_dfrbp_1 _7458_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net59),
    .D(_0324_),
    .Q_N(_3493_),
    .Q(\vgademo.b_sin[6] ));
 sg13g2_dfrbp_1 _7459_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net57),
    .D(net308),
    .Q_N(_3492_),
    .Q(\vgademo.b_sin[7] ));
 sg13g2_dfrbp_1 _7460_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net55),
    .D(_0326_),
    .Q_N(_3491_),
    .Q(\vgademo.b_sin[8] ));
 sg13g2_dfrbp_1 _7461_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net53),
    .D(_0327_),
    .Q_N(_3490_),
    .Q(\vgademo.b_sin[9] ));
 sg13g2_dfrbp_1 _7462_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net51),
    .D(_0328_),
    .Q_N(_3489_),
    .Q(\vgademo.b_sin[10] ));
 sg13g2_dfrbp_1 _7463_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net50),
    .D(_0329_),
    .Q_N(_3488_),
    .Q(\vgademo.b_sin[11] ));
 sg13g2_dfrbp_1 _7464_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net48),
    .D(net291),
    .Q_N(_3487_),
    .Q(\vgademo.plane_u[1] ));
 sg13g2_dfrbp_1 _7465_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net47),
    .D(_0331_),
    .Q_N(_3486_),
    .Q(\vgademo.plane_u[2] ));
 sg13g2_dfrbp_1 _7466_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net46),
    .D(_0332_),
    .Q_N(_3485_),
    .Q(\vgademo.plane_u[3] ));
 sg13g2_dfrbp_1 _7467_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net45),
    .D(_0333_),
    .Q_N(_3484_),
    .Q(\vgademo.plane_u[4] ));
 sg13g2_dfrbp_1 _7468_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net44),
    .D(_0334_),
    .Q_N(_3483_),
    .Q(\vgademo.plane_u[5] ));
 sg13g2_dfrbp_1 _7469_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net43),
    .D(_0335_),
    .Q_N(_3482_),
    .Q(\vgademo.plane_u[6] ));
 sg13g2_dfrbp_1 _7470_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net42),
    .D(_0336_),
    .Q_N(_3481_),
    .Q(\vgademo.plane_u[7] ));
 sg13g2_dfrbp_1 _7471_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net41),
    .D(_0337_),
    .Q_N(_3480_),
    .Q(\vgademo.plane_u[8] ));
 sg13g2_dfrbp_1 _7472_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net40),
    .D(_0338_),
    .Q_N(_3479_),
    .Q(\vgademo.plane_u[9] ));
 sg13g2_dfrbp_1 _7473_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net39),
    .D(_0339_),
    .Q_N(_3478_),
    .Q(\vgademo.plane_u[10] ));
 sg13g2_dfrbp_1 _7474_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net36),
    .D(net343),
    .Q_N(_0026_),
    .Q(\vgademo.plane_u[11] ));
 sg13g2_dfrbp_1 _7475_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net35),
    .D(_0341_),
    .Q_N(_0027_),
    .Q(\vgademo.plane_u[12] ));
 sg13g2_dfrbp_1 _7476_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net34),
    .D(net483),
    .Q_N(_0047_),
    .Q(\vgademo.plane_u[13] ));
 sg13g2_dfrbp_1 _7477_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net33),
    .D(_0343_),
    .Q_N(_0028_),
    .Q(\vgademo.plane_u[14] ));
 sg13g2_dfrbp_1 _7478_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net32),
    .D(_0344_),
    .Q_N(_0046_),
    .Q(\vgademo.plane_u[15] ));
 sg13g2_dfrbp_1 _7479_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net31),
    .D(_0345_),
    .Q_N(_0029_),
    .Q(\vgademo.plane_u[16] ));
 sg13g2_dfrbp_1 _7480_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net30),
    .D(_0346_),
    .Q_N(_0045_),
    .Q(\vgademo.plane_u[17] ));
 sg13g2_dfrbp_1 _7481_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net29),
    .D(_0347_),
    .Q_N(_0030_),
    .Q(\vgademo.plane_u[18] ));
 sg13g2_dfrbp_1 _7482_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net28),
    .D(net415),
    .Q_N(_0044_),
    .Q(\vgademo.plane_u[19] ));
 sg13g2_dfrbp_1 _7483_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net27),
    .D(_0349_),
    .Q_N(_0031_),
    .Q(\vgademo.plane_u[20] ));
 sg13g2_dfrbp_1 _7484_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net26),
    .D(net304),
    .Q_N(_3477_),
    .Q(\vgademo.plane_u[21] ));
 sg13g2_dfrbp_1 _7485_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net25),
    .D(_0351_),
    .Q_N(_3476_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7486_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net24),
    .D(_0352_),
    .Q_N(_3475_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7487_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net23),
    .D(net288),
    .Q_N(_3474_),
    .Q(\vgademo.plane_du[0] ));
 sg13g2_dfrbp_1 _7488_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net22),
    .D(net306),
    .Q_N(_3473_),
    .Q(\vgademo.plane_du[1] ));
 sg13g2_dfrbp_1 _7489_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net21),
    .D(net436),
    .Q_N(_3472_),
    .Q(\vgademo.plane_du[2] ));
 sg13g2_dfrbp_1 _7490_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net155),
    .D(net473),
    .Q_N(_0049_),
    .Q(\vgademo.plane_du[3] ));
 sg13g2_dfrbp_1 _7491_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net154),
    .D(net485),
    .Q_N(_0048_),
    .Q(\vgademo.plane_du[4] ));
 sg13g2_dfrbp_1 _7492_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net153),
    .D(_0358_),
    .Q_N(_0050_),
    .Q(\vgademo.plane_du[5] ));
 sg13g2_dfrbp_1 _7493_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0359_),
    .Q_N(_0051_),
    .Q(\vgademo.plane_du[6] ));
 sg13g2_dfrbp_1 _7494_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net151),
    .D(net352),
    .Q_N(_0052_),
    .Q(\vgademo.plane_du[7] ));
 sg13g2_dfrbp_1 _7495_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net150),
    .D(_0361_),
    .Q_N(_0053_),
    .Q(\vgademo.plane_du[8] ));
 sg13g2_dfrbp_1 _7496_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net149),
    .D(_0362_),
    .Q_N(_3471_),
    .Q(\vgademo.plane_du[9] ));
 sg13g2_dfrbp_1 _7497_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net148),
    .D(net535),
    .Q_N(_3470_),
    .Q(\vgademo.plane_du[10] ));
 sg13g2_dfrbp_1 _7498_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net121),
    .D(net235),
    .Q_N(_3469_),
    .Q(\vgademo.plane_u[0] ));
 sg13g2_tiehi _7303__16 (.L_HI(net16));
 sg13g2_tiehi _7302__17 (.L_HI(net17));
 sg13g2_tiehi _7301__18 (.L_HI(net18));
 sg13g2_tiehi _7300__19 (.L_HI(net19));
 sg13g2_tiehi _7299__20 (.L_HI(net20));
 sg13g2_tiehi _7489__21 (.L_HI(net21));
 sg13g2_tiehi _7488__22 (.L_HI(net22));
 sg13g2_tiehi _7487__23 (.L_HI(net23));
 sg13g2_tiehi _7486__24 (.L_HI(net24));
 sg13g2_tiehi _7485__25 (.L_HI(net25));
 sg13g2_tiehi _7484__26 (.L_HI(net26));
 sg13g2_tiehi _7483__27 (.L_HI(net27));
 sg13g2_tiehi _7482__28 (.L_HI(net28));
 sg13g2_tiehi _7481__29 (.L_HI(net29));
 sg13g2_tiehi _7480__30 (.L_HI(net30));
 sg13g2_tiehi _7479__31 (.L_HI(net31));
 sg13g2_tiehi _7478__32 (.L_HI(net32));
 sg13g2_tiehi _7477__33 (.L_HI(net33));
 sg13g2_tiehi _7476__34 (.L_HI(net34));
 sg13g2_tiehi _7475__35 (.L_HI(net35));
 sg13g2_tiehi _7474__36 (.L_HI(net36));
 sg13g2_tiehi _7206__37 (.L_HI(net37));
 sg13g2_tiehi _7240__38 (.L_HI(net38));
 sg13g2_tiehi _7473__39 (.L_HI(net39));
 sg13g2_tiehi _7472__40 (.L_HI(net40));
 sg13g2_tiehi _7471__41 (.L_HI(net41));
 sg13g2_tiehi _7470__42 (.L_HI(net42));
 sg13g2_tiehi _7469__43 (.L_HI(net43));
 sg13g2_tiehi _7468__44 (.L_HI(net44));
 sg13g2_tiehi _7467__45 (.L_HI(net45));
 sg13g2_tiehi _7466__46 (.L_HI(net46));
 sg13g2_tiehi _7465__47 (.L_HI(net47));
 sg13g2_tiehi _7464__48 (.L_HI(net48));
 sg13g2_tiehi _7271__49 (.L_HI(net49));
 sg13g2_tiehi _7463__50 (.L_HI(net50));
 sg13g2_tiehi _7462__51 (.L_HI(net51));
 sg13g2_tiehi _7239__52 (.L_HI(net52));
 sg13g2_tiehi _7461__53 (.L_HI(net53));
 sg13g2_tiehi _7238__54 (.L_HI(net54));
 sg13g2_tiehi _7460__55 (.L_HI(net55));
 sg13g2_tiehi _7237__56 (.L_HI(net56));
 sg13g2_tiehi _7459__57 (.L_HI(net57));
 sg13g2_tiehi _7236__58 (.L_HI(net58));
 sg13g2_tiehi _7458__59 (.L_HI(net59));
 sg13g2_tiehi _7235__60 (.L_HI(net60));
 sg13g2_tiehi _7457__61 (.L_HI(net61));
 sg13g2_tiehi _7234__62 (.L_HI(net62));
 sg13g2_tiehi _7456__63 (.L_HI(net63));
 sg13g2_tiehi _7233__64 (.L_HI(net64));
 sg13g2_tiehi _7455__65 (.L_HI(net65));
 sg13g2_tiehi _7232__66 (.L_HI(net66));
 sg13g2_tiehi _7454__67 (.L_HI(net67));
 sg13g2_tiehi _7231__68 (.L_HI(net68));
 sg13g2_tiehi _7453__69 (.L_HI(net69));
 sg13g2_tiehi _7230__70 (.L_HI(net70));
 sg13g2_tiehi _7452__71 (.L_HI(net71));
 sg13g2_tiehi _7229__72 (.L_HI(net72));
 sg13g2_tiehi _7451__73 (.L_HI(net73));
 sg13g2_tiehi _7228__74 (.L_HI(net74));
 sg13g2_tiehi _7450__75 (.L_HI(net75));
 sg13g2_tiehi _7227__76 (.L_HI(net76));
 sg13g2_tiehi _7449__77 (.L_HI(net77));
 sg13g2_tiehi _7448__78 (.L_HI(net78));
 sg13g2_tiehi _7447__79 (.L_HI(net79));
 sg13g2_tiehi _7446__80 (.L_HI(net80));
 sg13g2_tiehi _7445__81 (.L_HI(net81));
 sg13g2_tiehi _7444__82 (.L_HI(net82));
 sg13g2_tiehi _7443__83 (.L_HI(net83));
 sg13g2_tiehi _7442__84 (.L_HI(net84));
 sg13g2_tiehi _7441__85 (.L_HI(net85));
 sg13g2_tiehi _7440__86 (.L_HI(net86));
 sg13g2_tiehi _7439__87 (.L_HI(net87));
 sg13g2_tiehi _7438__88 (.L_HI(net88));
 sg13g2_tiehi _7437__89 (.L_HI(net89));
 sg13g2_tiehi _7436__90 (.L_HI(net90));
 sg13g2_tiehi _7354__91 (.L_HI(net91));
 sg13g2_tiehi _7355__92 (.L_HI(net92));
 sg13g2_tiehi _7356__93 (.L_HI(net93));
 sg13g2_tiehi _7435__94 (.L_HI(net94));
 sg13g2_tiehi _7434__95 (.L_HI(net95));
 sg13g2_tiehi _7433__96 (.L_HI(net96));
 sg13g2_tiehi _7218__97 (.L_HI(net97));
 sg13g2_tiehi _7432__98 (.L_HI(net98));
 sg13g2_tiehi _7217__99 (.L_HI(net99));
 sg13g2_tiehi _7431__100 (.L_HI(net100));
 sg13g2_tiehi _7216__101 (.L_HI(net101));
 sg13g2_tiehi _7430__102 (.L_HI(net102));
 sg13g2_tiehi _7215__103 (.L_HI(net103));
 sg13g2_tiehi _7429__104 (.L_HI(net104));
 sg13g2_tiehi _7214__105 (.L_HI(net105));
 sg13g2_tiehi _7428__106 (.L_HI(net106));
 sg13g2_tiehi _7213__107 (.L_HI(net107));
 sg13g2_tiehi _7427__108 (.L_HI(net108));
 sg13g2_tiehi _7212__109 (.L_HI(net109));
 sg13g2_tiehi _7426__110 (.L_HI(net110));
 sg13g2_tiehi _7211__111 (.L_HI(net111));
 sg13g2_tiehi _7425__112 (.L_HI(net112));
 sg13g2_tiehi _7210__113 (.L_HI(net113));
 sg13g2_tiehi _7424__114 (.L_HI(net114));
 sg13g2_tiehi _7209__115 (.L_HI(net115));
 sg13g2_tiehi _7423__116 (.L_HI(net116));
 sg13g2_tiehi _7208__117 (.L_HI(net117));
 sg13g2_tiehi _7422__118 (.L_HI(net118));
 sg13g2_tiehi _7207__119 (.L_HI(net119));
 sg13g2_tiehi _7421__120 (.L_HI(net120));
 sg13g2_tiehi _7498__121 (.L_HI(net121));
 sg13g2_tiehi _7390__122 (.L_HI(net122));
 sg13g2_tiehi _7389__123 (.L_HI(net123));
 sg13g2_tiehi _7353__124 (.L_HI(net124));
 sg13g2_tiehi _7352__125 (.L_HI(net125));
 sg13g2_tiehi _7351__126 (.L_HI(net126));
 sg13g2_tiehi _7350__127 (.L_HI(net127));
 sg13g2_tiehi _7349__128 (.L_HI(net128));
 sg13g2_tiehi _7348__129 (.L_HI(net129));
 sg13g2_tiehi _7347__130 (.L_HI(net130));
 sg13g2_tiehi _7346__131 (.L_HI(net131));
 sg13g2_tiehi _7345__132 (.L_HI(net132));
 sg13g2_tiehi _7344__133 (.L_HI(net133));
 sg13g2_tiehi _7343__134 (.L_HI(net134));
 sg13g2_tiehi _7342__135 (.L_HI(net135));
 sg13g2_tiehi _7341__136 (.L_HI(net136));
 sg13g2_tiehi _7340__137 (.L_HI(net137));
 sg13g2_tiehi _7339__138 (.L_HI(net138));
 sg13g2_tiehi _7338__139 (.L_HI(net139));
 sg13g2_tiehi _7337__140 (.L_HI(net140));
 sg13g2_tiehi _7336__141 (.L_HI(net141));
 sg13g2_tiehi _7335__142 (.L_HI(net142));
 sg13g2_tiehi _7334__143 (.L_HI(net143));
 sg13g2_tiehi _7333__144 (.L_HI(net144));
 sg13g2_tiehi _7332__145 (.L_HI(net145));
 sg13g2_tiehi _7331__146 (.L_HI(net146));
 sg13g2_tiehi _7330__147 (.L_HI(net147));
 sg13g2_tiehi _7497__148 (.L_HI(net148));
 sg13g2_tiehi _7496__149 (.L_HI(net149));
 sg13g2_tiehi _7495__150 (.L_HI(net150));
 sg13g2_tiehi _7494__151 (.L_HI(net151));
 sg13g2_tiehi _7493__152 (.L_HI(net152));
 sg13g2_tiehi _7492__153 (.L_HI(net153));
 sg13g2_tiehi _7491__154 (.L_HI(net154));
 sg13g2_tiehi _7490__155 (.L_HI(net155));
 sg13g2_tiehi _7312__156 (.L_HI(net156));
 sg13g2_tiehi _7311__157 (.L_HI(net157));
 sg13g2_tiehi _7310__158 (.L_HI(net158));
 sg13g2_tiehi _7309__159 (.L_HI(net159));
 sg13g2_tiehi _7308__160 (.L_HI(net160));
 sg13g2_tiehi _7307__161 (.L_HI(net161));
 sg13g2_tiehi _7306__162 (.L_HI(net162));
 sg13g2_tiehi _7305__163 (.L_HI(net163));
 sg13g2_tiehi tt_um_a1k0n_demo_164 (.L_HI(net164));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_a1k0n_demo_2 (.L_LO(net2));
 sg13g2_tielo tt_um_a1k0n_demo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_a1k0n_demo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_a1k0n_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_a1k0n_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_a1k0n_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_a1k0n_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_a1k0n_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_a1k0n_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_a1k0n_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_a1k0n_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_a1k0n_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_a1k0n_demo_14 (.L_LO(net14));
 sg13g2_tiehi _7304__15 (.L_HI(net15));
 sg13g2_buf_2 _7663_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_1 _7664_ (.A(\vgademo.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7665_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout896 (.A(_1825_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_1825_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_1803_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net901),
    .X(net899));
 sg13g2_buf_1 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_1770_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net904),
    .X(net902));
 sg13g2_buf_1 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_1679_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_1913_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_1473_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_1 fanout908 (.A(net909),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_1493_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net912),
    .X(net910));
 sg13g2_buf_1 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_1492_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net915),
    .X(net913));
 sg13g2_buf_1 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_2556_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_1619_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net921),
    .X(net917));
 sg13g2_buf_1 fanout918 (.A(net921),
    .X(net918));
 sg13g2_buf_4 fanout919 (.X(net919),
    .A(net921));
 sg13g2_buf_1 fanout920 (.A(net921),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_1502_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_1501_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_1501_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_1 fanout925 (.A(net926),
    .X(net925));
 sg13g2_buf_1 fanout926 (.A(_1501_),
    .X(net926));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(_2411_));
 sg13g2_buf_2 fanout928 (.A(_1476_),
    .X(net928));
 sg13g2_buf_1 fanout929 (.A(_1476_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_1476_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(net934),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_1475_));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(_1372_));
 sg13g2_buf_1 fanout936 (.A(_1372_),
    .X(net936));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_1511_));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(_1478_));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(net940));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(_1477_));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(_1479_));
 sg13g2_buf_2 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_0703_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_0633_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_1823_),
    .X(net947));
 sg13g2_buf_1 fanout948 (.A(_1823_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_0629_),
    .X(net949));
 sg13g2_buf_1 fanout950 (.A(_0629_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(net954),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(net954),
    .X(net952));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(net954));
 sg13g2_buf_2 fanout954 (.A(_1340_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_4 fanout956 (.X(net956),
    .A(_1341_));
 sg13g2_buf_2 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_1 fanout958 (.A(_1337_),
    .X(net958));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(_0861_));
 sg13g2_buf_2 fanout960 (.A(_1339_),
    .X(net960));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(_1296_));
 sg13g2_buf_2 fanout962 (.A(_1296_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_1295_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(net965),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_0828_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_0828_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net969),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_2798_),
    .X(net969));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(net971));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(net973));
 sg13g2_buf_2 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_2798_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net976),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_0596_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_0578_),
    .X(net978));
 sg13g2_buf_1 fanout979 (.A(_0578_),
    .X(net979));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(net982));
 sg13g2_buf_2 fanout981 (.A(net982),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_0577_),
    .X(net982));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(net984));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(_2491_));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(net987));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(net987));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(_0584_));
 sg13g2_buf_2 fanout988 (.A(net992),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(net991),
    .X(net989));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(net991));
 sg13g2_buf_2 fanout991 (.A(net992),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_2485_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_1391_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_1208_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_1079_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(net999),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_4 fanout999 (.X(net999),
    .A(_0595_));
 sg13g2_buf_2 fanout1000 (.A(net1007),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(net1007),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(net1005),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(net1005),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(net1007),
    .X(net1006));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(_0581_));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(net1009));
 sg13g2_buf_4 fanout1009 (.X(net1009),
    .A(net1010));
 sg13g2_buf_4 fanout1010 (.X(net1010),
    .A(net1011));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(_0580_));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(net1013));
 sg13g2_buf_2 fanout1013 (.A(_0665_),
    .X(net1013));
 sg13g2_buf_4 fanout1014 (.X(net1014),
    .A(net1015));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(_0664_));
 sg13g2_buf_2 fanout1016 (.A(net1017),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_0648_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(net1020),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(net1020));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(_0594_));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(net1023),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_0593_),
    .X(net1023));
 sg13g2_buf_4 fanout1024 (.X(net1024),
    .A(net1026));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_0583_),
    .X(net1026));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(_0582_));
 sg13g2_buf_2 fanout1028 (.A(_1078_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_1078_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(net1032),
    .X(net1031));
 sg13g2_buf_4 fanout1032 (.X(net1032),
    .A(_0661_));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(_3289_));
 sg13g2_buf_4 fanout1034 (.X(net1034),
    .A(_3289_));
 sg13g2_buf_2 fanout1035 (.A(_3288_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_3288_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_0705_),
    .X(net1037));
 sg13g2_buf_4 fanout1038 (.X(net1038),
    .A(_0632_));
 sg13g2_buf_2 fanout1039 (.A(_0631_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_2227_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_1056_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_3225_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(net1044),
    .X(net1043));
 sg13g2_buf_1 fanout1044 (.A(_3224_),
    .X(net1044));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(_3199_));
 sg13g2_buf_2 fanout1046 (.A(net1047),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_3180_),
    .X(net1047));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(_3178_));
 sg13g2_buf_2 fanout1049 (.A(_3178_),
    .X(net1049));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(\vgademo.b_sin[11] ));
 sg13g2_buf_2 fanout1051 (.A(net551),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(\vgademo.plane_dx_div.r[25] ));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(\vgademo.b_cos[10] ));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(\vgademo.b_cos[9] ));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(\vgademo.b_cos[6] ));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(net1058));
 sg13g2_buf_2 fanout1058 (.A(net507),
    .X(net1058));
 sg13g2_buf_4 fanout1059 (.X(net1059),
    .A(\vgademo.v_count[9] ));
 sg13g2_buf_2 fanout1060 (.A(\vgademo.v_count[7] ),
    .X(net1060));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(\vgademo.v_count[6] ));
 sg13g2_buf_2 fanout1062 (.A(net1063),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(net487),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(\vgademo.v_count[3] ),
    .X(net1064));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(\vgademo.v_count[2] ));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(net556));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(\vgademo.a_scrolly[11] ));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(net1069));
 sg13g2_buf_4 fanout1069 (.X(net1069),
    .A(\vgademo.a_scrolly[10] ));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(net1071));
 sg13g2_buf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(net1073),
    .X(net1072));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(\vgademo.a_scrolly[9] ));
 sg13g2_buf_2 fanout1074 (.A(net1075),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(\vgademo.a_scrolly[8] ),
    .X(net1076));
 sg13g2_buf_4 fanout1077 (.X(net1077),
    .A(net546));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(\vgademo.a_scrolly[7] ));
 sg13g2_buf_2 fanout1079 (.A(net1080),
    .X(net1079));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1081));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(\vgademo.a_scrolly[6] ));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net564));
 sg13g2_buf_2 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(\vgademo.a_scrolly[5] ));
 sg13g2_buf_2 fanout1085 (.A(net1087),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_4 fanout1087 (.X(net1087),
    .A(\vgademo.a_scrolly[4] ));
 sg13g2_buf_2 fanout1088 (.A(net1089),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(\vgademo.a_scrolly[3] ),
    .X(net1089));
 sg13g2_buf_4 fanout1090 (.X(net1090),
    .A(\vgademo.a_scrolly[3] ));
 sg13g2_buf_2 fanout1091 (.A(\vgademo.a_scrolly[3] ),
    .X(net1091));
 sg13g2_buf_4 fanout1092 (.X(net1092),
    .A(net530));
 sg13g2_buf_2 fanout1093 (.A(\vgademo.h_count[3] ),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(\vgademo.h_count[3] ),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(\vgademo.h_count[2] ),
    .X(net1095));
 sg13g2_buf_4 fanout1096 (.X(net1096),
    .A(net1097));
 sg13g2_buf_4 fanout1097 (.X(net1097),
    .A(net541));
 sg13g2_buf_4 fanout1098 (.X(net1098),
    .A(net166));
 sg13g2_buf_4 fanout1099 (.X(net1099),
    .A(net1100));
 sg13g2_buf_4 fanout1100 (.X(net1100),
    .A(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_buf_2 fanout1101 (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(net1102));
 sg13g2_buf_4 fanout1103 (.X(net1103),
    .A(\vgademo.soundtrack.pulse_vol[2] ));
 sg13g2_buf_2 fanout1104 (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(\vgademo.audio_snare_frames[3] ),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(net1110),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(net1110),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(\vgademo.audio_snare_frames[2] ),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_1 fanout1113 (.A(net1114),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(\vgademo.audio_snare_frames[1] ),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(\vgademo.audio_snare_frames[0] ),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(net1120),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(\vgademo.plane_dx_div.q[9] ),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(net539),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(net539),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(net552),
    .X(net1123));
 sg13g2_buf_1 fanout1124 (.A(\vgademo.plane_dx_div.q[7] ),
    .X(net1124));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(net351));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(net421));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(net278));
 sg13g2_buf_2 fanout1128 (.A(net278),
    .X(net1128));
 sg13g2_buf_4 fanout1129 (.X(net1129),
    .A(net484));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(net523));
 sg13g2_buf_4 fanout1131 (.X(net1131),
    .A(\vgademo.audio_songpos[7] ));
 sg13g2_buf_4 fanout1132 (.X(net1132),
    .A(\vgademo.audio_songpos[6] ));
 sg13g2_buf_2 fanout1133 (.A(\vgademo.audio_songpos[6] ),
    .X(net1133));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(net1136));
 sg13g2_buf_2 fanout1135 (.A(net1136),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(\vgademo.audio_songpos[5] ),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(net1139),
    .X(net1137));
 sg13g2_buf_1 fanout1138 (.A(net1139),
    .X(net1138));
 sg13g2_buf_4 fanout1139 (.X(net1139),
    .A(\vgademo.audio_songpos[4] ));
 sg13g2_buf_4 fanout1140 (.X(net1140),
    .A(net1142));
 sg13g2_buf_2 fanout1141 (.A(net1143),
    .X(net1141));
 sg13g2_buf_1 fanout1142 (.A(net1143),
    .X(net1142));
 sg13g2_buf_4 fanout1143 (.X(net1143),
    .A(\vgademo.audio_songpos[3] ));
 sg13g2_buf_4 fanout1144 (.X(net1144),
    .A(net1146));
 sg13g2_buf_2 fanout1145 (.A(net1146),
    .X(net1145));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(\vgademo.audio_songpos[2] ));
 sg13g2_buf_2 fanout1147 (.A(net1149),
    .X(net1147));
 sg13g2_buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(\vgademo.audio_songpos[1] ),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(net1151),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(\vgademo.audio_songpos[0] ),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sg13g2_buf_1 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_buf_2 fanout1154 (.A(net569),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(net1157),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(\vgademo.linelfsr[0] ),
    .X(net1157));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(net1168));
 sg13g2_buf_4 fanout1159 (.X(net1159),
    .A(net1168));
 sg13g2_buf_4 fanout1160 (.X(net1160),
    .A(net1164));
 sg13g2_buf_4 fanout1161 (.X(net1161),
    .A(net1164));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(net1163));
 sg13g2_buf_4 fanout1163 (.X(net1163),
    .A(net1164));
 sg13g2_buf_4 fanout1164 (.X(net1164),
    .A(net1168));
 sg13g2_buf_4 fanout1165 (.X(net1165),
    .A(net1167));
 sg13g2_buf_2 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_buf_4 fanout1167 (.X(net1167),
    .A(net1168));
 sg13g2_buf_4 fanout1168 (.X(net1168),
    .A(rst_n));
 sg13g2_buf_4 fanout1169 (.X(net1169),
    .A(net1170));
 sg13g2_buf_2 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_4 fanout1171 (.X(net1171),
    .A(net1175));
 sg13g2_buf_4 fanout1172 (.X(net1172),
    .A(net1175));
 sg13g2_buf_4 fanout1173 (.X(net1173),
    .A(net1174));
 sg13g2_buf_4 fanout1174 (.X(net1174),
    .A(net1175));
 sg13g2_buf_2 fanout1175 (.A(net1180),
    .X(net1175));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(net1177));
 sg13g2_buf_4 fanout1177 (.X(net1177),
    .A(net1180));
 sg13g2_buf_4 fanout1178 (.X(net1178),
    .A(net1179));
 sg13g2_buf_4 fanout1179 (.X(net1179),
    .A(net1180));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(rst_n));
 sg13g2_buf_4 fanout1181 (.X(net1181),
    .A(net1182));
 sg13g2_buf_2 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_4 fanout1183 (.X(net1183),
    .A(rst_n));
 sg13g2_tielo tt_um_a1k0n_demo_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_0_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_49_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_50_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_52_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_53_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_3_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_46_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_48_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_8_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_12_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_13_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_14_clk));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_30_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_32_clk));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_40_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_34_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_37_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_38_clk));
 sg13g2_inv_4 clkload32 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_21_clk));
 sg13g2_inv_1 clkload36 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload37 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_23_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload41 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload42 (.A(clknet_leaf_28_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vgademo.soundtrack.sample_div_[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold2 (.A(\vgademo.h_count[0] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold3 (.A(\vgademo.soundtrack.noise_lfsr[11] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0179_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold5 (.A(\vgademo.soundtrack.noise_lfsr[1] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0169_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0081_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0181_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0083_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0174_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold11 (.A(\vgademo.soundtrack.tick_div_[0] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0161_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0082_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0176_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0105_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0187_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0103_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0185_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0102_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0184_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0087_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0094_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0800_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0170_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0092_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0131_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0086_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0095_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0801_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0171_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0089_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0100_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0803_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0180_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold35 (.A(\vgademo.soundtrack.tick_div[6] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0798_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0167_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0109_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0208_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold40 (.A(\vgademo.soundtrack.noise_lfsr[10] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0178_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vgademo.plane_dx_div.q[3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0669_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0090_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold45 (.A(\vgademo.soundtrack.pulse_osc_p[10] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0198_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0104_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0186_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0088_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vgademo.soundtrack.sigma_delta_accum[0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold51 (.A(\vgademo.soundtrack.sample_div[4] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold52 (.A(\vgademo.soundtrack.sample_div_[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0084_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vgademo.soundtrack.pulse_osc_p[1] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0189_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold56 (.A(\vgademo.soundtrack.tick_div[7] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0168_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0096_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0172_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold60 (.A(\vgademo.soundtrack.sample_div[8] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold61 (.A(\vgademo.soundtrack.sample_div_[8] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold62 (.A(\vgademo.soundtrack.tick_div[4] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0165_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold64 (.A(\vgademo.soundtrack.sample_div[7] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold65 (.A(\vgademo.soundtrack.sample_div_[7] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold66 (.A(\vgademo.soundtrack.pulse_osc_p[9] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0941_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0197_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold69 (.A(\vgademo.plane_u[0] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold70 (.A(_3161_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0364_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0110_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold73 (.A(\vgademo.a_sin[0] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold74 (.A(\vgademo.soundtrack.pulse_osc_p[13] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0201_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold76 (.A(\vgademo.soundtrack.noise_lfsr[4] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0173_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold78 (.A(\vgademo.soundtrack.tick_div[2] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0163_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold80 (.A(\vgademo.soundtrack.noise_lfsr[13] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0182_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold82 (.A(\vgademo.soundtrack.tri_osc_p[0] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0209_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold84 (.A(audio),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0160_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold86 (.A(\vgademo.a_cos[0] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0257_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold88 (.A(\vgademo.soundtrack.tick_div[3] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0164_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold90 (.A(\vgademo.soundtrack.sample_div[3] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold91 (.A(\vgademo.soundtrack.sample_div_[3] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold92 (.A(\vgademo.v_count[2] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0247_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold94 (.A(\vgademo.soundtrack.sample_div[1] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold95 (.A(\vgademo.soundtrack.sample_div_[1] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold96 (.A(\vgademo.soundtrack.noise_lfsr[7] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0175_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold98 (.A(\vgademo.plane_dx_div.r[20] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0310_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold100 (.A(\vgademo.soundtrack.tick_div[5] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0166_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold102 (.A(\vgademo.plane_u[20] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vgademo.soundtrack.pulse_osc_p[8] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0196_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold105 (.A(\vgademo.soundtrack.pulse_osc_p[11] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold106 (.A(\vgademo.soundtrack.pulse_osc_p[0] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0085_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0124_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold109 (.A(\vgademo.soundtrack.sample_div[5] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0108_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0106_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0091_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0107_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold114 (.A(\vgademo.plane_dx_div.q[4] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold115 (.A(\vgademo.plane_dx_div.d[22] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold116 (.A(\vgademo.audio_kick_frames[2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0204_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold118 (.A(\vgademo.plane_dx_div.r[24] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold119 (.A(\vgademo.b_sin[5] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold120 (.A(\vgademo.soundtrack.sample_div[9] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold121 (.A(\vgademo.plane_dx_div.d[20] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold122 (.A(\vgademo.plane_dx_div.d[18] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold123 (.A(\vgademo.plane_du[0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0353_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold125 (.A(\vgademo.plane_u[4] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold126 (.A(\vgademo.plane_u[1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0330_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold128 (.A(\vgademo.soundtrack.noise_lfsr[0] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0183_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold130 (.A(\vgademo.soundtrack.tri_osc_p[11] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0220_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold132 (.A(\vgademo.plane_dx_div.d[23] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold133 (.A(\vgademo.plane_u[6] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold134 (.A(\vgademo.plane_dx_div.d[24] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold135 (.A(\vgademo.plane_dx_div.r[21] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0034_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0006_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold138 (.A(\vgademo.a_cos[2] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold139 (.A(\vgademo.plane_u[21] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0350_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold141 (.A(\vgademo.plane_du[1] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0354_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold143 (.A(\vgademo.b_sin[7] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0325_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold145 (.A(\vgademo.soundtrack.tri_osc_p[10] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0219_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold147 (.A(\vgademo.a_sin[5] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold148 (.A(\vgademo.scanline_audio_sample[0] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold149 (.A(\vgademo.a_cos[1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0258_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold151 (.A(\vgademo.soundtrack.pulse_osc_p[7] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold152 (.A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0192_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold154 (.A(\vgademo.audio_beat_out[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold155 (.A(\vgademo.linelfsr[6] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0117_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0033_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold158 (.A(_3293_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold159 (.A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold160 (.A(\vgademo.a_sin[3] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold161 (.A(\vgademo.b_cos[0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0294_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold163 (.A(\vgademo.plane_dx_div.i[0] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0658_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0143_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold166 (.A(\vgademo.soundtrack.noise_lfsr[8] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0177_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold168 (.A(\vgademo.scanline_audio_sample[2] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold169 (.A(\vgademo.soundtrack.tri_osc_p[12] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold170 (.A(\vgademo.plane_dx_div.r[16] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0306_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold172 (.A(\vgademo.soundtrack.tri_osc_p[9] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0218_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold174 (.A(\vgademo.plane_dx_div.r[18] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0308_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0021_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0254_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold178 (.A(\vgademo.plane_u[11] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0340_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold180 (.A(\vgademo.plane_dx_div.r[19] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold181 (.A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0194_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold183 (.A(\vgademo.a_sin[1] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0273_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold185 (.A(\vgademo.a_sin[2] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold186 (.A(\vgademo.scanline_audio_sample[5] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold187 (.A(\vgademo.plane_dx_div.q[6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0360_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold189 (.A(\vgademo.scanline_audio_sample[1] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold190 (.A(\vgademo.plane_u[2] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold191 (.A(\vgademo.a_sin[4] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0276_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold193 (.A(\vgademo.b_cos[3] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0297_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold195 (.A(\vgademo.plane_dx_div.r[17] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0307_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold197 (.A(\vgademo.soundtrack.pulse_osc_p[2] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0190_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold199 (.A(\vgademo.b_sin[1] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0319_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold201 (.A(\vgademo.plane_u[7] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold202 (.A(\vgademo.soundtrack.tri_osc_p[14] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0223_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold204 (.A(\vgademo.linelfsr[7] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0118_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold206 (.A(\vgademo.linelfsr[3] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0113_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold208 (.A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold209 (.A(\vgademo.plane_dx_div.d[19] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold210 (.A(\vgademo.plane_u[10] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold211 (.A(\vgademo.audio_beat_out[1] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold212 (.A(\vgademo.linelfsr[8] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0119_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold214 (.A(\vgademo.plane_u[12] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold215 (.A(_2978_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0014_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold217 (.A(_1261_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold218 (.A(\vgademo.b_sin[2] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold219 (.A(\vgademo.plane_dx_div.r[22] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0312_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0038_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold222 (.A(_3307_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0010_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold224 (.A(\vgademo.plane_u[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold225 (.A(\vgademo.b_sin[3] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold226 (.A(_2745_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold227 (.A(\vgademo.plane_dx_div.d[17] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold228 (.A(\vgademo.b_cos[4] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0298_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold230 (.A(\vgademo.a_cos[3] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold231 (.A(\vgademo.linelfsr[4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold232 (.A(\vgademo.plane_u[8] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold233 (.A(\vgademo.plane_dx_div.r[23] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold234 (.A(\vgademo.soundtrack.tri_osc_p[7] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold235 (.A(\vgademo.soundtrack.tri_osc_p[13] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0224_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold237 (.A(\vgademo.linelfsr[11] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0121_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold239 (.A(\vgademo.linelfsr[9] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0120_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold241 (.A(\vgademo.plane_dx_div.i[3] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0680_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold243 (.A(\vgademo.audio_beat_out[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0149_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold245 (.A(\vgademo.linelfsr[12] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold246 (.A(\vgademo.plane_dx_div.d[21] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold247 (.A(\vgademo.b_sin[0] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold248 (.A(\vgademo.linelfsr[5] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold249 (.A(\vgademo.soundtrack.tri_osc_p[4] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold250 (.A(\vgademo.plane_u[19] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0348_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold252 (.A(\vgademo.plane_dx_div.r[25] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold253 (.A(\vgademo.h_count[4] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold254 (.A(\vgademo.plane_u[16] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold255 (.A(_3042_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold256 (.A(\vgademo.plane_u[5] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold257 (.A(\vgademo.plane_dx_div.q[5] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold258 (.A(\vgademo.a_cos[14] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0305_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold260 (.A(\vgademo.soundtrack.tri_osc_p[2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold261 (.A(\vgademo.scanline_audio_sample[4] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold262 (.A(\vgademo.b_sin[6] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold263 (.A(_2764_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold264 (.A(\vgademo.soundtrack.tri_osc_p[8] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold265 (.A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold266 (.A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold267 (.A(\vgademo.soundtrack.tri_osc_p[3] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0212_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold269 (.A(\vgademo.soundtrack.tri_osc_p[5] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0214_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold271 (.A(\vgademo.plane_du[2] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0355_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold273 (.A(\vgademo.a_cos[12] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0303_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold275 (.A(\vgademo.a_cos[11] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0302_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold277 (.A(\vgademo.b_cos[1] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold278 (.A(_2498_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold279 (.A(\vgademo.a_cos[5] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold280 (.A(\vgademo.a_cos[4] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold281 (.A(\vgademo.soundtrack.tri_osc_i[8] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold282 (.A(\vgademo.plane_u[9] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold283 (.A(\vgademo.scanline_audio_sample[6] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold284 (.A(\vgademo.soundtrack.tri_osc_p[6] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold285 (.A(\vgademo.b_cos[2] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0296_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold287 (.A(\vgademo.a_sin[11] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0018_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0253_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold290 (.A(\vgademo.soundtrack.tri_osc_i[2] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0073_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold292 (.A(_1249_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0248_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold294 (.A(\vgademo.plane_dx_div.d[16] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold295 (.A(\vgademo.soundtrack.sample_div[6] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold296 (.A(\vgademo.audio_kick_frames[1] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold297 (.A(\vgademo.a_cos[10] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0301_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold299 (.A(\vgademo.plane_u[14] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold300 (.A(_3012_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold301 (.A(\vgademo.soundtrack.sample_div[2] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0570_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold303 (.A(\vgademo.soundtrack.sample_div_[2] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold304 (.A(\vgademo.soundtrack.tri_osc_p[1] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold305 (.A(\vgademo.b_cos[5] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0015_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold307 (.A(_1230_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold308 (.A(\vgademo.plane_du[3] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0356_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold310 (.A(\vgademo.a_sin[9] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold311 (.A(\vgademo.plane_u[17] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold312 (.A(\vgademo.bayer_j[1] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold313 (.A(\vgademo.plane_dx_div.i[2] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0679_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold315 (.A(\vgademo.a_sin[10] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold316 (.A(\vgademo.b_sin[10] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold317 (.A(_2790_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold318 (.A(\vgademo.plane_u[13] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0342_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0023_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0357_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold322 (.A(\vgademo.b_sin[8] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold323 (.A(\vgademo.v_count[4] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0249_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold325 (.A(\vgademo.soundtrack.tick_div[1] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0797_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0162_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0064_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold329 (.A(\vgademo.b_sin[4] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold330 (.A(_2751_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold331 (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold332 (.A(\vgademo.a_cos[7] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold333 (.A(\vgademo.a_sin[12] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold334 (.A(_2784_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold335 (.A(\vgademo.soundtrack.sigma_delta_accum[7] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold336 (.A(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold337 (.A(\vgademo.a_sin[13] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold338 (.A(\vgademo.plane_u[15] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold339 (.A(\vgademo.v_count[5] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0250_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold341 (.A(\vgademo.audio_beat_out[4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0691_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold343 (.A(\vgademo.a_sin[14] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold344 (.A(\vgademo.plane_u[18] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold345 (.A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold346 (.A(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold347 (.A(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold348 (.A(\vgademo.a_sin[6] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold349 (.A(\vgademo.soundtrack.sigma_delta_accum[11] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold350 (.A(\vgademo.soundtrack.sigma_delta_accum[12] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold351 (.A(\vgademo.a_cos[6] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold352 (.A(\vgademo.soundtrack.tri_osc_i[3] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0154_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold354 (.A(\vgademo.v_count[9] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold355 (.A(\vgademo.soundtrack.sigma_delta_accum[13] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold356 (.A(\vgademo.soundtrack.sigma_delta_accum[6] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold357 (.A(\vgademo.soundtrack.sigma_delta_accum_[6] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold358 (.A(\vgademo.a_cos[9] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold359 (.A(\vgademo.plane_dx[3] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0668_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold361 (.A(\vgademo.soundtrack.sigma_delta_accum[9] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold362 (.A(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold363 (.A(\vgademo.soundtrack.sigma_delta_accum[3] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold364 (.A(\vgademo.soundtrack.sigma_delta_accum_[3] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold365 (.A(\vgademo.soundtrack.sigma_delta_accum[8] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0060_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold367 (.A(\vgademo.plane_dx[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0667_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold369 (.A(\vgademo.soundtrack.sigma_delta_accum[4] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold370 (.A(\vgademo.plane_du[10] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0363_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0032_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold373 (.A(\vgademo.linelfsr[2] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold374 (.A(\vgademo.soundtrack.sigma_delta_accum[1] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold375 (.A(\vgademo.plane_dx_div.q[8] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0674_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold377 (.A(\vgademo.h_count[1] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold378 (.A(\vgademo.a_cos[13] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold379 (.A(\vgademo.plane_dx_div.i[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold380 (.A(\vgademo.plane_dx[0] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold381 (.A(\vgademo.plane_du[5] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold382 (.A(\vgademo.a_scrolly[7] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0238_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold384 (.A(\vgademo.soundtrack.pulse_osc_p[12] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold385 (.A(\vgademo.soundtrack.sigma_delta_accum[2] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0061_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold387 (.A(\vgademo.b_sin[11] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold388 (.A(\vgademo.plane_dx_div.q[7] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold389 (.A(\vgademo.a_sin[7] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold390 (.A(\vgademo.a_scrolly[13] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0244_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold392 (.A(\vgademo.a_scrolly[12] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0243_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0036_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold395 (.A(_3302_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0008_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold397 (.A(\vgademo.soundtrack.sigma_delta_accum[14] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0037_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold399 (.A(\vgademo.scanline_audio_sample[3] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold400 (.A(\vgademo.a_scrolly[5] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0016_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0251_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold403 (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold404 (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold405 (.A(\vgademo.linelfsr[1] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold406 (.A(\vgademo.soundtrack.sigma_delta_accum[5] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0019_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0242_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold409 (.A(\vgademo.a_cos[8] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold410 (.A(\vgademo.a_sin[8] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0035_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold412 (.A(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0079_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold414 (.A(\vgademo.plane_du[6] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold415 (.A(\vgademo.plane_du[8] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0074_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0237_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold418 (.A(\vgademo.bayer_j[0] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold419 (.A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .X(net583));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_fill_2 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_fill_1 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_4 FILLER_8_67 ();
 sg13g2_fill_2 FILLER_8_71 ();
 sg13g2_fill_2 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_96 ();
 sg13g2_decap_4 FILLER_8_103 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_128 ();
 sg13g2_decap_8 FILLER_8_135 ();
 sg13g2_decap_8 FILLER_8_142 ();
 sg13g2_decap_8 FILLER_8_149 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_decap_8 FILLER_8_163 ();
 sg13g2_decap_8 FILLER_8_170 ();
 sg13g2_decap_8 FILLER_8_177 ();
 sg13g2_decap_8 FILLER_8_184 ();
 sg13g2_decap_8 FILLER_8_191 ();
 sg13g2_decap_8 FILLER_8_198 ();
 sg13g2_decap_8 FILLER_8_205 ();
 sg13g2_decap_8 FILLER_8_212 ();
 sg13g2_decap_8 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_decap_8 FILLER_8_240 ();
 sg13g2_decap_8 FILLER_8_247 ();
 sg13g2_decap_8 FILLER_8_254 ();
 sg13g2_decap_8 FILLER_8_261 ();
 sg13g2_decap_8 FILLER_8_268 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_decap_8 FILLER_8_289 ();
 sg13g2_decap_8 FILLER_8_296 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_317 ();
 sg13g2_fill_1 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_decap_8 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_8_414 ();
 sg13g2_decap_8 FILLER_8_421 ();
 sg13g2_decap_8 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_8_435 ();
 sg13g2_decap_8 FILLER_8_442 ();
 sg13g2_decap_8 FILLER_8_449 ();
 sg13g2_decap_8 FILLER_8_456 ();
 sg13g2_decap_8 FILLER_8_463 ();
 sg13g2_decap_8 FILLER_8_470 ();
 sg13g2_decap_8 FILLER_8_477 ();
 sg13g2_decap_8 FILLER_8_484 ();
 sg13g2_decap_8 FILLER_8_491 ();
 sg13g2_decap_8 FILLER_8_498 ();
 sg13g2_decap_8 FILLER_8_505 ();
 sg13g2_decap_8 FILLER_8_512 ();
 sg13g2_decap_8 FILLER_8_519 ();
 sg13g2_decap_8 FILLER_8_526 ();
 sg13g2_decap_8 FILLER_8_533 ();
 sg13g2_decap_8 FILLER_8_540 ();
 sg13g2_decap_8 FILLER_8_547 ();
 sg13g2_decap_8 FILLER_8_554 ();
 sg13g2_decap_8 FILLER_8_561 ();
 sg13g2_decap_8 FILLER_8_568 ();
 sg13g2_decap_8 FILLER_8_575 ();
 sg13g2_decap_8 FILLER_8_582 ();
 sg13g2_decap_8 FILLER_8_589 ();
 sg13g2_decap_8 FILLER_8_596 ();
 sg13g2_decap_8 FILLER_8_603 ();
 sg13g2_decap_8 FILLER_8_610 ();
 sg13g2_decap_8 FILLER_8_617 ();
 sg13g2_decap_8 FILLER_8_624 ();
 sg13g2_decap_8 FILLER_8_631 ();
 sg13g2_decap_8 FILLER_8_638 ();
 sg13g2_decap_8 FILLER_8_645 ();
 sg13g2_decap_8 FILLER_8_652 ();
 sg13g2_decap_8 FILLER_8_659 ();
 sg13g2_decap_8 FILLER_8_666 ();
 sg13g2_decap_8 FILLER_8_673 ();
 sg13g2_decap_8 FILLER_8_680 ();
 sg13g2_decap_8 FILLER_8_687 ();
 sg13g2_decap_8 FILLER_8_694 ();
 sg13g2_decap_8 FILLER_8_701 ();
 sg13g2_decap_8 FILLER_8_708 ();
 sg13g2_decap_8 FILLER_8_715 ();
 sg13g2_decap_8 FILLER_8_722 ();
 sg13g2_decap_8 FILLER_8_729 ();
 sg13g2_decap_8 FILLER_8_736 ();
 sg13g2_decap_8 FILLER_8_743 ();
 sg13g2_decap_8 FILLER_8_750 ();
 sg13g2_decap_8 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_764 ();
 sg13g2_decap_8 FILLER_8_771 ();
 sg13g2_decap_8 FILLER_8_778 ();
 sg13g2_decap_8 FILLER_8_785 ();
 sg13g2_decap_8 FILLER_8_792 ();
 sg13g2_decap_8 FILLER_8_799 ();
 sg13g2_decap_8 FILLER_8_806 ();
 sg13g2_decap_8 FILLER_8_813 ();
 sg13g2_decap_8 FILLER_8_820 ();
 sg13g2_decap_8 FILLER_8_827 ();
 sg13g2_decap_8 FILLER_8_834 ();
 sg13g2_decap_8 FILLER_8_841 ();
 sg13g2_decap_8 FILLER_8_848 ();
 sg13g2_decap_8 FILLER_8_855 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_44 ();
 sg13g2_fill_2 FILLER_9_58 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_decap_4 FILLER_9_91 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_decap_4 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_142 ();
 sg13g2_decap_8 FILLER_9_149 ();
 sg13g2_decap_8 FILLER_9_156 ();
 sg13g2_decap_8 FILLER_9_163 ();
 sg13g2_decap_8 FILLER_9_170 ();
 sg13g2_decap_8 FILLER_9_177 ();
 sg13g2_decap_8 FILLER_9_184 ();
 sg13g2_decap_8 FILLER_9_191 ();
 sg13g2_decap_8 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_fill_2 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_8 FILLER_9_262 ();
 sg13g2_decap_8 FILLER_9_269 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_fill_1 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_283 ();
 sg13g2_fill_2 FILLER_9_290 ();
 sg13g2_fill_1 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_decap_8 FILLER_9_416 ();
 sg13g2_decap_8 FILLER_9_423 ();
 sg13g2_decap_8 FILLER_9_430 ();
 sg13g2_decap_8 FILLER_9_437 ();
 sg13g2_decap_8 FILLER_9_444 ();
 sg13g2_decap_8 FILLER_9_451 ();
 sg13g2_decap_8 FILLER_9_458 ();
 sg13g2_decap_8 FILLER_9_465 ();
 sg13g2_decap_8 FILLER_9_472 ();
 sg13g2_decap_8 FILLER_9_479 ();
 sg13g2_decap_8 FILLER_9_486 ();
 sg13g2_decap_8 FILLER_9_493 ();
 sg13g2_decap_8 FILLER_9_500 ();
 sg13g2_decap_8 FILLER_9_507 ();
 sg13g2_decap_8 FILLER_9_514 ();
 sg13g2_decap_8 FILLER_9_521 ();
 sg13g2_decap_8 FILLER_9_528 ();
 sg13g2_decap_8 FILLER_9_535 ();
 sg13g2_decap_8 FILLER_9_542 ();
 sg13g2_decap_8 FILLER_9_549 ();
 sg13g2_decap_8 FILLER_9_556 ();
 sg13g2_decap_8 FILLER_9_563 ();
 sg13g2_decap_8 FILLER_9_570 ();
 sg13g2_decap_8 FILLER_9_577 ();
 sg13g2_decap_8 FILLER_9_584 ();
 sg13g2_decap_8 FILLER_9_591 ();
 sg13g2_decap_8 FILLER_9_598 ();
 sg13g2_decap_8 FILLER_9_605 ();
 sg13g2_decap_8 FILLER_9_612 ();
 sg13g2_decap_8 FILLER_9_619 ();
 sg13g2_decap_8 FILLER_9_626 ();
 sg13g2_decap_8 FILLER_9_633 ();
 sg13g2_decap_8 FILLER_9_640 ();
 sg13g2_decap_8 FILLER_9_647 ();
 sg13g2_decap_8 FILLER_9_654 ();
 sg13g2_decap_8 FILLER_9_661 ();
 sg13g2_decap_8 FILLER_9_668 ();
 sg13g2_decap_8 FILLER_9_675 ();
 sg13g2_decap_8 FILLER_9_682 ();
 sg13g2_decap_8 FILLER_9_689 ();
 sg13g2_decap_8 FILLER_9_696 ();
 sg13g2_decap_8 FILLER_9_703 ();
 sg13g2_decap_8 FILLER_9_710 ();
 sg13g2_decap_8 FILLER_9_717 ();
 sg13g2_decap_8 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_745 ();
 sg13g2_decap_8 FILLER_9_752 ();
 sg13g2_decap_8 FILLER_9_759 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_decap_8 FILLER_9_773 ();
 sg13g2_decap_8 FILLER_9_780 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_decap_8 FILLER_9_822 ();
 sg13g2_decap_8 FILLER_9_829 ();
 sg13g2_decap_8 FILLER_9_836 ();
 sg13g2_decap_8 FILLER_9_843 ();
 sg13g2_decap_8 FILLER_9_850 ();
 sg13g2_decap_4 FILLER_9_857 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_4 FILLER_10_35 ();
 sg13g2_fill_2 FILLER_10_78 ();
 sg13g2_decap_8 FILLER_10_90 ();
 sg13g2_fill_1 FILLER_10_97 ();
 sg13g2_fill_2 FILLER_10_115 ();
 sg13g2_fill_1 FILLER_10_127 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_decap_8 FILLER_10_155 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_171 ();
 sg13g2_fill_2 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_decap_4 FILLER_10_264 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_fill_2 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_310 ();
 sg13g2_decap_4 FILLER_10_316 ();
 sg13g2_fill_2 FILLER_10_320 ();
 sg13g2_fill_2 FILLER_10_326 ();
 sg13g2_decap_4 FILLER_10_333 ();
 sg13g2_fill_2 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_fill_2 FILLER_10_418 ();
 sg13g2_fill_1 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_10_433 ();
 sg13g2_decap_8 FILLER_10_440 ();
 sg13g2_decap_8 FILLER_10_447 ();
 sg13g2_decap_8 FILLER_10_454 ();
 sg13g2_decap_8 FILLER_10_461 ();
 sg13g2_decap_8 FILLER_10_468 ();
 sg13g2_decap_8 FILLER_10_475 ();
 sg13g2_decap_8 FILLER_10_482 ();
 sg13g2_decap_8 FILLER_10_489 ();
 sg13g2_decap_8 FILLER_10_496 ();
 sg13g2_decap_8 FILLER_10_503 ();
 sg13g2_decap_8 FILLER_10_510 ();
 sg13g2_decap_8 FILLER_10_517 ();
 sg13g2_decap_8 FILLER_10_524 ();
 sg13g2_decap_8 FILLER_10_531 ();
 sg13g2_decap_8 FILLER_10_538 ();
 sg13g2_decap_8 FILLER_10_545 ();
 sg13g2_decap_8 FILLER_10_552 ();
 sg13g2_decap_8 FILLER_10_559 ();
 sg13g2_decap_8 FILLER_10_566 ();
 sg13g2_decap_8 FILLER_10_573 ();
 sg13g2_decap_8 FILLER_10_580 ();
 sg13g2_decap_8 FILLER_10_587 ();
 sg13g2_decap_8 FILLER_10_594 ();
 sg13g2_decap_8 FILLER_10_601 ();
 sg13g2_decap_8 FILLER_10_608 ();
 sg13g2_decap_8 FILLER_10_615 ();
 sg13g2_decap_8 FILLER_10_622 ();
 sg13g2_decap_8 FILLER_10_629 ();
 sg13g2_decap_8 FILLER_10_636 ();
 sg13g2_decap_8 FILLER_10_643 ();
 sg13g2_decap_8 FILLER_10_650 ();
 sg13g2_decap_8 FILLER_10_657 ();
 sg13g2_decap_8 FILLER_10_664 ();
 sg13g2_decap_8 FILLER_10_671 ();
 sg13g2_decap_8 FILLER_10_678 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_692 ();
 sg13g2_decap_8 FILLER_10_699 ();
 sg13g2_decap_8 FILLER_10_706 ();
 sg13g2_decap_8 FILLER_10_713 ();
 sg13g2_decap_8 FILLER_10_720 ();
 sg13g2_decap_8 FILLER_10_727 ();
 sg13g2_decap_8 FILLER_10_734 ();
 sg13g2_decap_8 FILLER_10_741 ();
 sg13g2_decap_8 FILLER_10_748 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_decap_8 FILLER_10_762 ();
 sg13g2_decap_8 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_776 ();
 sg13g2_decap_8 FILLER_10_783 ();
 sg13g2_decap_8 FILLER_10_790 ();
 sg13g2_decap_8 FILLER_10_797 ();
 sg13g2_decap_8 FILLER_10_804 ();
 sg13g2_decap_8 FILLER_10_811 ();
 sg13g2_decap_8 FILLER_10_818 ();
 sg13g2_decap_8 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_832 ();
 sg13g2_decap_8 FILLER_10_839 ();
 sg13g2_decap_8 FILLER_10_846 ();
 sg13g2_decap_8 FILLER_10_853 ();
 sg13g2_fill_2 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_4 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_65 ();
 sg13g2_fill_2 FILLER_11_80 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_104 ();
 sg13g2_fill_1 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_decap_8 FILLER_11_160 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_195 ();
 sg13g2_fill_1 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_fill_2 FILLER_11_225 ();
 sg13g2_fill_2 FILLER_11_241 ();
 sg13g2_fill_2 FILLER_11_292 ();
 sg13g2_decap_4 FILLER_11_328 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_4 FILLER_11_369 ();
 sg13g2_fill_2 FILLER_11_373 ();
 sg13g2_fill_2 FILLER_11_396 ();
 sg13g2_fill_1 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_437 ();
 sg13g2_decap_8 FILLER_11_444 ();
 sg13g2_decap_8 FILLER_11_451 ();
 sg13g2_decap_8 FILLER_11_458 ();
 sg13g2_decap_8 FILLER_11_465 ();
 sg13g2_decap_8 FILLER_11_472 ();
 sg13g2_decap_8 FILLER_11_479 ();
 sg13g2_decap_8 FILLER_11_486 ();
 sg13g2_decap_8 FILLER_11_493 ();
 sg13g2_decap_8 FILLER_11_500 ();
 sg13g2_decap_8 FILLER_11_507 ();
 sg13g2_decap_8 FILLER_11_514 ();
 sg13g2_decap_8 FILLER_11_521 ();
 sg13g2_decap_8 FILLER_11_528 ();
 sg13g2_decap_8 FILLER_11_535 ();
 sg13g2_decap_8 FILLER_11_542 ();
 sg13g2_decap_8 FILLER_11_549 ();
 sg13g2_decap_8 FILLER_11_556 ();
 sg13g2_decap_8 FILLER_11_563 ();
 sg13g2_decap_8 FILLER_11_570 ();
 sg13g2_decap_8 FILLER_11_577 ();
 sg13g2_decap_8 FILLER_11_584 ();
 sg13g2_decap_8 FILLER_11_591 ();
 sg13g2_decap_8 FILLER_11_598 ();
 sg13g2_decap_8 FILLER_11_605 ();
 sg13g2_decap_8 FILLER_11_612 ();
 sg13g2_decap_8 FILLER_11_619 ();
 sg13g2_decap_8 FILLER_11_626 ();
 sg13g2_decap_8 FILLER_11_633 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_654 ();
 sg13g2_decap_8 FILLER_11_661 ();
 sg13g2_decap_8 FILLER_11_668 ();
 sg13g2_decap_8 FILLER_11_675 ();
 sg13g2_decap_8 FILLER_11_682 ();
 sg13g2_decap_8 FILLER_11_689 ();
 sg13g2_decap_8 FILLER_11_696 ();
 sg13g2_decap_8 FILLER_11_703 ();
 sg13g2_decap_8 FILLER_11_710 ();
 sg13g2_decap_8 FILLER_11_717 ();
 sg13g2_decap_8 FILLER_11_724 ();
 sg13g2_decap_8 FILLER_11_731 ();
 sg13g2_decap_8 FILLER_11_738 ();
 sg13g2_decap_8 FILLER_11_745 ();
 sg13g2_decap_8 FILLER_11_752 ();
 sg13g2_decap_8 FILLER_11_759 ();
 sg13g2_decap_8 FILLER_11_766 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_787 ();
 sg13g2_decap_8 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_decap_8 FILLER_11_808 ();
 sg13g2_decap_8 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_8 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_4 FILLER_11_857 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_fill_1 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_127 ();
 sg13g2_decap_4 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_138 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_4 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_162 ();
 sg13g2_fill_2 FILLER_12_169 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_2 FILLER_12_296 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_decap_4 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_fill_1 FILLER_12_322 ();
 sg13g2_fill_2 FILLER_12_340 ();
 sg13g2_fill_1 FILLER_12_342 ();
 sg13g2_decap_4 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_364 ();
 sg13g2_fill_2 FILLER_12_385 ();
 sg13g2_fill_1 FILLER_12_387 ();
 sg13g2_fill_2 FILLER_12_392 ();
 sg13g2_fill_1 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_424 ();
 sg13g2_decap_8 FILLER_12_460 ();
 sg13g2_decap_8 FILLER_12_467 ();
 sg13g2_decap_8 FILLER_12_474 ();
 sg13g2_decap_8 FILLER_12_481 ();
 sg13g2_decap_8 FILLER_12_488 ();
 sg13g2_decap_8 FILLER_12_495 ();
 sg13g2_decap_8 FILLER_12_502 ();
 sg13g2_decap_8 FILLER_12_509 ();
 sg13g2_decap_8 FILLER_12_516 ();
 sg13g2_decap_8 FILLER_12_523 ();
 sg13g2_decap_8 FILLER_12_530 ();
 sg13g2_decap_8 FILLER_12_537 ();
 sg13g2_decap_8 FILLER_12_544 ();
 sg13g2_decap_8 FILLER_12_551 ();
 sg13g2_decap_8 FILLER_12_558 ();
 sg13g2_decap_8 FILLER_12_565 ();
 sg13g2_decap_8 FILLER_12_572 ();
 sg13g2_decap_8 FILLER_12_579 ();
 sg13g2_decap_8 FILLER_12_586 ();
 sg13g2_decap_8 FILLER_12_593 ();
 sg13g2_decap_8 FILLER_12_600 ();
 sg13g2_decap_8 FILLER_12_607 ();
 sg13g2_decap_8 FILLER_12_614 ();
 sg13g2_decap_8 FILLER_12_621 ();
 sg13g2_decap_8 FILLER_12_628 ();
 sg13g2_decap_8 FILLER_12_635 ();
 sg13g2_decap_8 FILLER_12_642 ();
 sg13g2_decap_8 FILLER_12_649 ();
 sg13g2_decap_8 FILLER_12_656 ();
 sg13g2_decap_8 FILLER_12_663 ();
 sg13g2_decap_8 FILLER_12_670 ();
 sg13g2_decap_8 FILLER_12_677 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_decap_8 FILLER_12_691 ();
 sg13g2_decap_8 FILLER_12_698 ();
 sg13g2_decap_8 FILLER_12_705 ();
 sg13g2_decap_8 FILLER_12_712 ();
 sg13g2_decap_8 FILLER_12_719 ();
 sg13g2_decap_8 FILLER_12_726 ();
 sg13g2_decap_8 FILLER_12_733 ();
 sg13g2_decap_8 FILLER_12_740 ();
 sg13g2_decap_8 FILLER_12_747 ();
 sg13g2_decap_8 FILLER_12_754 ();
 sg13g2_decap_8 FILLER_12_761 ();
 sg13g2_decap_8 FILLER_12_768 ();
 sg13g2_decap_8 FILLER_12_775 ();
 sg13g2_decap_8 FILLER_12_782 ();
 sg13g2_decap_8 FILLER_12_789 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_decap_8 FILLER_12_803 ();
 sg13g2_decap_8 FILLER_12_810 ();
 sg13g2_decap_8 FILLER_12_817 ();
 sg13g2_decap_8 FILLER_12_824 ();
 sg13g2_decap_8 FILLER_12_831 ();
 sg13g2_decap_8 FILLER_12_838 ();
 sg13g2_decap_8 FILLER_12_845 ();
 sg13g2_decap_8 FILLER_12_852 ();
 sg13g2_fill_2 FILLER_12_859 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_54 ();
 sg13g2_decap_4 FILLER_13_61 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_decap_8 FILLER_13_92 ();
 sg13g2_fill_1 FILLER_13_99 ();
 sg13g2_decap_4 FILLER_13_105 ();
 sg13g2_fill_2 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_115 ();
 sg13g2_decap_8 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_decap_4 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_216 ();
 sg13g2_decap_8 FILLER_13_223 ();
 sg13g2_decap_4 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_fill_2 FILLER_13_261 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_4 FILLER_13_293 ();
 sg13g2_decap_4 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_335 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_fill_2 FILLER_13_369 ();
 sg13g2_fill_1 FILLER_13_371 ();
 sg13g2_fill_2 FILLER_13_385 ();
 sg13g2_fill_1 FILLER_13_387 ();
 sg13g2_fill_2 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_436 ();
 sg13g2_decap_8 FILLER_13_456 ();
 sg13g2_decap_8 FILLER_13_463 ();
 sg13g2_decap_8 FILLER_13_470 ();
 sg13g2_decap_8 FILLER_13_477 ();
 sg13g2_decap_8 FILLER_13_484 ();
 sg13g2_decap_8 FILLER_13_491 ();
 sg13g2_decap_8 FILLER_13_498 ();
 sg13g2_decap_8 FILLER_13_505 ();
 sg13g2_decap_8 FILLER_13_512 ();
 sg13g2_decap_8 FILLER_13_519 ();
 sg13g2_decap_8 FILLER_13_526 ();
 sg13g2_decap_8 FILLER_13_533 ();
 sg13g2_decap_8 FILLER_13_540 ();
 sg13g2_decap_8 FILLER_13_547 ();
 sg13g2_decap_8 FILLER_13_554 ();
 sg13g2_decap_8 FILLER_13_561 ();
 sg13g2_decap_8 FILLER_13_568 ();
 sg13g2_decap_8 FILLER_13_575 ();
 sg13g2_decap_8 FILLER_13_582 ();
 sg13g2_decap_8 FILLER_13_589 ();
 sg13g2_decap_8 FILLER_13_596 ();
 sg13g2_decap_8 FILLER_13_603 ();
 sg13g2_decap_8 FILLER_13_610 ();
 sg13g2_decap_8 FILLER_13_617 ();
 sg13g2_decap_8 FILLER_13_624 ();
 sg13g2_decap_8 FILLER_13_631 ();
 sg13g2_decap_8 FILLER_13_638 ();
 sg13g2_decap_8 FILLER_13_645 ();
 sg13g2_decap_8 FILLER_13_652 ();
 sg13g2_decap_8 FILLER_13_659 ();
 sg13g2_decap_8 FILLER_13_666 ();
 sg13g2_decap_8 FILLER_13_673 ();
 sg13g2_decap_8 FILLER_13_680 ();
 sg13g2_decap_8 FILLER_13_687 ();
 sg13g2_decap_8 FILLER_13_694 ();
 sg13g2_decap_8 FILLER_13_701 ();
 sg13g2_decap_8 FILLER_13_708 ();
 sg13g2_decap_8 FILLER_13_715 ();
 sg13g2_decap_8 FILLER_13_722 ();
 sg13g2_decap_8 FILLER_13_729 ();
 sg13g2_decap_8 FILLER_13_736 ();
 sg13g2_decap_8 FILLER_13_743 ();
 sg13g2_decap_8 FILLER_13_750 ();
 sg13g2_decap_8 FILLER_13_757 ();
 sg13g2_decap_8 FILLER_13_764 ();
 sg13g2_decap_8 FILLER_13_771 ();
 sg13g2_decap_8 FILLER_13_778 ();
 sg13g2_decap_8 FILLER_13_785 ();
 sg13g2_decap_8 FILLER_13_792 ();
 sg13g2_decap_8 FILLER_13_799 ();
 sg13g2_decap_8 FILLER_13_806 ();
 sg13g2_decap_8 FILLER_13_813 ();
 sg13g2_decap_8 FILLER_13_820 ();
 sg13g2_decap_8 FILLER_13_827 ();
 sg13g2_decap_8 FILLER_13_834 ();
 sg13g2_decap_8 FILLER_13_841 ();
 sg13g2_decap_8 FILLER_13_848 ();
 sg13g2_decap_8 FILLER_13_855 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_51 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_decap_4 FILLER_14_153 ();
 sg13g2_fill_1 FILLER_14_157 ();
 sg13g2_fill_2 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_fill_2 FILLER_14_187 ();
 sg13g2_fill_1 FILLER_14_189 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_242 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_268 ();
 sg13g2_fill_2 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_297 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_4 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_4 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_4 FILLER_14_416 ();
 sg13g2_fill_1 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_437 ();
 sg13g2_decap_8 FILLER_14_465 ();
 sg13g2_decap_8 FILLER_14_472 ();
 sg13g2_decap_8 FILLER_14_479 ();
 sg13g2_decap_8 FILLER_14_486 ();
 sg13g2_decap_8 FILLER_14_493 ();
 sg13g2_decap_8 FILLER_14_500 ();
 sg13g2_decap_8 FILLER_14_507 ();
 sg13g2_decap_8 FILLER_14_514 ();
 sg13g2_decap_8 FILLER_14_521 ();
 sg13g2_decap_8 FILLER_14_528 ();
 sg13g2_decap_8 FILLER_14_535 ();
 sg13g2_decap_8 FILLER_14_542 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_decap_8 FILLER_14_556 ();
 sg13g2_decap_8 FILLER_14_563 ();
 sg13g2_decap_8 FILLER_14_570 ();
 sg13g2_decap_8 FILLER_14_577 ();
 sg13g2_decap_8 FILLER_14_584 ();
 sg13g2_decap_8 FILLER_14_591 ();
 sg13g2_decap_8 FILLER_14_598 ();
 sg13g2_decap_8 FILLER_14_605 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_619 ();
 sg13g2_decap_8 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_633 ();
 sg13g2_decap_8 FILLER_14_640 ();
 sg13g2_decap_8 FILLER_14_647 ();
 sg13g2_decap_8 FILLER_14_654 ();
 sg13g2_decap_8 FILLER_14_661 ();
 sg13g2_decap_8 FILLER_14_668 ();
 sg13g2_decap_8 FILLER_14_675 ();
 sg13g2_decap_8 FILLER_14_682 ();
 sg13g2_decap_8 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_696 ();
 sg13g2_decap_8 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_710 ();
 sg13g2_decap_8 FILLER_14_717 ();
 sg13g2_decap_8 FILLER_14_724 ();
 sg13g2_decap_8 FILLER_14_731 ();
 sg13g2_decap_8 FILLER_14_738 ();
 sg13g2_decap_8 FILLER_14_745 ();
 sg13g2_decap_8 FILLER_14_752 ();
 sg13g2_decap_8 FILLER_14_759 ();
 sg13g2_decap_8 FILLER_14_766 ();
 sg13g2_decap_8 FILLER_14_773 ();
 sg13g2_decap_8 FILLER_14_780 ();
 sg13g2_decap_8 FILLER_14_787 ();
 sg13g2_decap_8 FILLER_14_794 ();
 sg13g2_decap_8 FILLER_14_801 ();
 sg13g2_decap_8 FILLER_14_808 ();
 sg13g2_decap_8 FILLER_14_815 ();
 sg13g2_decap_8 FILLER_14_822 ();
 sg13g2_decap_8 FILLER_14_829 ();
 sg13g2_decap_8 FILLER_14_836 ();
 sg13g2_decap_8 FILLER_14_843 ();
 sg13g2_decap_8 FILLER_14_850 ();
 sg13g2_decap_4 FILLER_14_857 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_149 ();
 sg13g2_fill_2 FILLER_15_171 ();
 sg13g2_fill_2 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_191 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_decap_4 FILLER_15_304 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_decap_4 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_4 FILLER_15_380 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_fill_2 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_416 ();
 sg13g2_decap_4 FILLER_15_423 ();
 sg13g2_fill_1 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_437 ();
 sg13g2_fill_2 FILLER_15_444 ();
 sg13g2_decap_8 FILLER_15_464 ();
 sg13g2_decap_8 FILLER_15_471 ();
 sg13g2_decap_8 FILLER_15_478 ();
 sg13g2_decap_8 FILLER_15_485 ();
 sg13g2_decap_8 FILLER_15_492 ();
 sg13g2_decap_8 FILLER_15_499 ();
 sg13g2_decap_8 FILLER_15_506 ();
 sg13g2_decap_8 FILLER_15_513 ();
 sg13g2_decap_8 FILLER_15_520 ();
 sg13g2_decap_8 FILLER_15_527 ();
 sg13g2_decap_8 FILLER_15_534 ();
 sg13g2_decap_8 FILLER_15_541 ();
 sg13g2_decap_8 FILLER_15_548 ();
 sg13g2_decap_8 FILLER_15_555 ();
 sg13g2_decap_8 FILLER_15_562 ();
 sg13g2_decap_8 FILLER_15_569 ();
 sg13g2_decap_8 FILLER_15_576 ();
 sg13g2_decap_8 FILLER_15_583 ();
 sg13g2_decap_8 FILLER_15_590 ();
 sg13g2_decap_8 FILLER_15_597 ();
 sg13g2_decap_8 FILLER_15_604 ();
 sg13g2_decap_8 FILLER_15_611 ();
 sg13g2_decap_8 FILLER_15_618 ();
 sg13g2_decap_8 FILLER_15_625 ();
 sg13g2_decap_8 FILLER_15_632 ();
 sg13g2_decap_8 FILLER_15_639 ();
 sg13g2_decap_8 FILLER_15_646 ();
 sg13g2_decap_8 FILLER_15_653 ();
 sg13g2_decap_8 FILLER_15_660 ();
 sg13g2_decap_8 FILLER_15_667 ();
 sg13g2_decap_8 FILLER_15_674 ();
 sg13g2_decap_8 FILLER_15_681 ();
 sg13g2_decap_8 FILLER_15_688 ();
 sg13g2_decap_8 FILLER_15_695 ();
 sg13g2_decap_8 FILLER_15_702 ();
 sg13g2_decap_8 FILLER_15_709 ();
 sg13g2_decap_8 FILLER_15_716 ();
 sg13g2_decap_8 FILLER_15_723 ();
 sg13g2_decap_8 FILLER_15_730 ();
 sg13g2_decap_8 FILLER_15_737 ();
 sg13g2_decap_8 FILLER_15_744 ();
 sg13g2_decap_8 FILLER_15_751 ();
 sg13g2_decap_8 FILLER_15_758 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_8 FILLER_15_772 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_8 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_793 ();
 sg13g2_decap_8 FILLER_15_800 ();
 sg13g2_decap_8 FILLER_15_807 ();
 sg13g2_decap_8 FILLER_15_814 ();
 sg13g2_decap_8 FILLER_15_821 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_decap_8 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_849 ();
 sg13g2_decap_4 FILLER_15_856 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_96 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_decap_8 FILLER_16_157 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_decap_4 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_1 FILLER_16_207 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_246 ();
 sg13g2_decap_4 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_299 ();
 sg13g2_decap_4 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_4 FILLER_16_326 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_decap_4 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_373 ();
 sg13g2_fill_1 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_fill_1 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_466 ();
 sg13g2_decap_8 FILLER_16_473 ();
 sg13g2_decap_8 FILLER_16_480 ();
 sg13g2_decap_8 FILLER_16_487 ();
 sg13g2_decap_8 FILLER_16_494 ();
 sg13g2_decap_8 FILLER_16_501 ();
 sg13g2_decap_8 FILLER_16_508 ();
 sg13g2_decap_8 FILLER_16_515 ();
 sg13g2_decap_8 FILLER_16_522 ();
 sg13g2_decap_8 FILLER_16_529 ();
 sg13g2_decap_8 FILLER_16_536 ();
 sg13g2_decap_8 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_550 ();
 sg13g2_decap_8 FILLER_16_557 ();
 sg13g2_decap_8 FILLER_16_564 ();
 sg13g2_decap_8 FILLER_16_571 ();
 sg13g2_decap_8 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_585 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_599 ();
 sg13g2_decap_8 FILLER_16_606 ();
 sg13g2_decap_8 FILLER_16_613 ();
 sg13g2_decap_8 FILLER_16_620 ();
 sg13g2_decap_8 FILLER_16_627 ();
 sg13g2_decap_8 FILLER_16_634 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_648 ();
 sg13g2_decap_8 FILLER_16_655 ();
 sg13g2_decap_8 FILLER_16_662 ();
 sg13g2_decap_8 FILLER_16_669 ();
 sg13g2_decap_8 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_decap_8 FILLER_16_704 ();
 sg13g2_decap_8 FILLER_16_711 ();
 sg13g2_decap_8 FILLER_16_718 ();
 sg13g2_decap_8 FILLER_16_725 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_decap_8 FILLER_16_774 ();
 sg13g2_decap_8 FILLER_16_781 ();
 sg13g2_decap_8 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_795 ();
 sg13g2_decap_8 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_809 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_851 ();
 sg13g2_decap_4 FILLER_16_858 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_fill_2 FILLER_17_30 ();
 sg13g2_decap_4 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_decap_4 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_1 FILLER_17_204 ();
 sg13g2_decap_4 FILLER_17_225 ();
 sg13g2_fill_1 FILLER_17_229 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_decap_4 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_decap_4 FILLER_17_401 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_4 FILLER_17_435 ();
 sg13g2_fill_1 FILLER_17_439 ();
 sg13g2_decap_8 FILLER_17_449 ();
 sg13g2_decap_8 FILLER_17_456 ();
 sg13g2_fill_2 FILLER_17_472 ();
 sg13g2_fill_1 FILLER_17_474 ();
 sg13g2_decap_8 FILLER_17_493 ();
 sg13g2_decap_8 FILLER_17_500 ();
 sg13g2_decap_8 FILLER_17_507 ();
 sg13g2_decap_8 FILLER_17_514 ();
 sg13g2_decap_8 FILLER_17_521 ();
 sg13g2_decap_8 FILLER_17_528 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_decap_8 FILLER_17_542 ();
 sg13g2_decap_8 FILLER_17_549 ();
 sg13g2_decap_8 FILLER_17_556 ();
 sg13g2_decap_8 FILLER_17_563 ();
 sg13g2_decap_8 FILLER_17_570 ();
 sg13g2_decap_8 FILLER_17_577 ();
 sg13g2_decap_8 FILLER_17_584 ();
 sg13g2_decap_8 FILLER_17_591 ();
 sg13g2_decap_8 FILLER_17_598 ();
 sg13g2_decap_8 FILLER_17_605 ();
 sg13g2_decap_8 FILLER_17_612 ();
 sg13g2_decap_8 FILLER_17_619 ();
 sg13g2_decap_8 FILLER_17_626 ();
 sg13g2_decap_8 FILLER_17_633 ();
 sg13g2_decap_8 FILLER_17_640 ();
 sg13g2_decap_8 FILLER_17_647 ();
 sg13g2_decap_8 FILLER_17_654 ();
 sg13g2_decap_8 FILLER_17_661 ();
 sg13g2_decap_8 FILLER_17_668 ();
 sg13g2_decap_8 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_682 ();
 sg13g2_decap_8 FILLER_17_689 ();
 sg13g2_decap_8 FILLER_17_696 ();
 sg13g2_decap_8 FILLER_17_703 ();
 sg13g2_decap_8 FILLER_17_710 ();
 sg13g2_decap_8 FILLER_17_717 ();
 sg13g2_decap_8 FILLER_17_724 ();
 sg13g2_decap_8 FILLER_17_731 ();
 sg13g2_decap_8 FILLER_17_738 ();
 sg13g2_decap_8 FILLER_17_745 ();
 sg13g2_decap_8 FILLER_17_752 ();
 sg13g2_decap_8 FILLER_17_759 ();
 sg13g2_decap_8 FILLER_17_766 ();
 sg13g2_decap_8 FILLER_17_773 ();
 sg13g2_decap_8 FILLER_17_780 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_decap_8 FILLER_17_794 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_decap_8 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_decap_8 FILLER_17_836 ();
 sg13g2_decap_8 FILLER_17_843 ();
 sg13g2_decap_8 FILLER_17_850 ();
 sg13g2_decap_4 FILLER_17_857 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_23 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_39 ();
 sg13g2_fill_2 FILLER_18_76 ();
 sg13g2_fill_1 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_decap_4 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_4 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_4 FILLER_18_305 ();
 sg13g2_decap_4 FILLER_18_320 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_fill_2 FILLER_18_353 ();
 sg13g2_decap_4 FILLER_18_456 ();
 sg13g2_decap_8 FILLER_18_505 ();
 sg13g2_decap_8 FILLER_18_512 ();
 sg13g2_decap_8 FILLER_18_519 ();
 sg13g2_decap_8 FILLER_18_526 ();
 sg13g2_decap_8 FILLER_18_533 ();
 sg13g2_decap_8 FILLER_18_540 ();
 sg13g2_decap_8 FILLER_18_547 ();
 sg13g2_decap_8 FILLER_18_554 ();
 sg13g2_decap_8 FILLER_18_561 ();
 sg13g2_decap_8 FILLER_18_568 ();
 sg13g2_decap_8 FILLER_18_575 ();
 sg13g2_decap_8 FILLER_18_582 ();
 sg13g2_decap_8 FILLER_18_589 ();
 sg13g2_decap_8 FILLER_18_596 ();
 sg13g2_decap_8 FILLER_18_603 ();
 sg13g2_decap_8 FILLER_18_610 ();
 sg13g2_decap_8 FILLER_18_617 ();
 sg13g2_decap_8 FILLER_18_624 ();
 sg13g2_decap_8 FILLER_18_631 ();
 sg13g2_decap_8 FILLER_18_638 ();
 sg13g2_decap_8 FILLER_18_645 ();
 sg13g2_decap_8 FILLER_18_652 ();
 sg13g2_decap_8 FILLER_18_659 ();
 sg13g2_decap_8 FILLER_18_666 ();
 sg13g2_decap_8 FILLER_18_673 ();
 sg13g2_decap_8 FILLER_18_680 ();
 sg13g2_decap_8 FILLER_18_687 ();
 sg13g2_decap_8 FILLER_18_694 ();
 sg13g2_decap_8 FILLER_18_701 ();
 sg13g2_decap_8 FILLER_18_708 ();
 sg13g2_decap_8 FILLER_18_715 ();
 sg13g2_decap_8 FILLER_18_722 ();
 sg13g2_decap_8 FILLER_18_729 ();
 sg13g2_decap_8 FILLER_18_736 ();
 sg13g2_decap_8 FILLER_18_743 ();
 sg13g2_decap_8 FILLER_18_750 ();
 sg13g2_decap_8 FILLER_18_757 ();
 sg13g2_decap_8 FILLER_18_764 ();
 sg13g2_decap_8 FILLER_18_771 ();
 sg13g2_decap_8 FILLER_18_778 ();
 sg13g2_decap_8 FILLER_18_785 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_decap_8 FILLER_18_799 ();
 sg13g2_decap_8 FILLER_18_806 ();
 sg13g2_decap_8 FILLER_18_813 ();
 sg13g2_decap_8 FILLER_18_820 ();
 sg13g2_decap_8 FILLER_18_827 ();
 sg13g2_decap_8 FILLER_18_834 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_848 ();
 sg13g2_decap_8 FILLER_18_855 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_11 ();
 sg13g2_fill_2 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_decap_4 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_120 ();
 sg13g2_decap_8 FILLER_19_127 ();
 sg13g2_decap_8 FILLER_19_134 ();
 sg13g2_decap_4 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_4 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_fill_2 FILLER_19_251 ();
 sg13g2_fill_1 FILLER_19_253 ();
 sg13g2_fill_2 FILLER_19_290 ();
 sg13g2_fill_2 FILLER_19_297 ();
 sg13g2_decap_4 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_395 ();
 sg13g2_fill_1 FILLER_19_401 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_4 FILLER_19_417 ();
 sg13g2_decap_8 FILLER_19_425 ();
 sg13g2_fill_2 FILLER_19_432 ();
 sg13g2_decap_8 FILLER_19_439 ();
 sg13g2_decap_4 FILLER_19_446 ();
 sg13g2_fill_2 FILLER_19_450 ();
 sg13g2_fill_1 FILLER_19_478 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_536 ();
 sg13g2_decap_8 FILLER_19_543 ();
 sg13g2_decap_8 FILLER_19_550 ();
 sg13g2_decap_8 FILLER_19_557 ();
 sg13g2_decap_8 FILLER_19_564 ();
 sg13g2_decap_8 FILLER_19_571 ();
 sg13g2_decap_8 FILLER_19_578 ();
 sg13g2_decap_8 FILLER_19_585 ();
 sg13g2_decap_8 FILLER_19_592 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_decap_8 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_620 ();
 sg13g2_decap_8 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_634 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_decap_8 FILLER_19_648 ();
 sg13g2_decap_8 FILLER_19_655 ();
 sg13g2_decap_8 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_676 ();
 sg13g2_decap_8 FILLER_19_683 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_decap_8 FILLER_19_697 ();
 sg13g2_decap_8 FILLER_19_704 ();
 sg13g2_decap_8 FILLER_19_711 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_decap_8 FILLER_19_732 ();
 sg13g2_decap_8 FILLER_19_739 ();
 sg13g2_decap_8 FILLER_19_746 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_767 ();
 sg13g2_decap_8 FILLER_19_774 ();
 sg13g2_decap_8 FILLER_19_781 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_decap_8 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_8 FILLER_19_823 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_decap_8 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_844 ();
 sg13g2_decap_8 FILLER_19_851 ();
 sg13g2_decap_4 FILLER_19_858 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_48 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_decap_4 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_2 FILLER_20_195 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_229 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_fill_1 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_4 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_decap_4 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_4 FILLER_20_396 ();
 sg13g2_fill_2 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_fill_2 FILLER_20_451 ();
 sg13g2_fill_2 FILLER_20_484 ();
 sg13g2_fill_2 FILLER_20_522 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_fill_2 FILLER_20_560 ();
 sg13g2_decap_4 FILLER_20_579 ();
 sg13g2_fill_2 FILLER_20_583 ();
 sg13g2_decap_8 FILLER_20_594 ();
 sg13g2_decap_8 FILLER_20_601 ();
 sg13g2_decap_8 FILLER_20_608 ();
 sg13g2_decap_8 FILLER_20_615 ();
 sg13g2_decap_8 FILLER_20_622 ();
 sg13g2_decap_8 FILLER_20_629 ();
 sg13g2_decap_8 FILLER_20_636 ();
 sg13g2_decap_8 FILLER_20_643 ();
 sg13g2_decap_8 FILLER_20_650 ();
 sg13g2_decap_8 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_671 ();
 sg13g2_decap_8 FILLER_20_678 ();
 sg13g2_decap_8 FILLER_20_685 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_decap_8 FILLER_20_706 ();
 sg13g2_decap_8 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_720 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_decap_8 FILLER_20_734 ();
 sg13g2_decap_8 FILLER_20_741 ();
 sg13g2_decap_8 FILLER_20_748 ();
 sg13g2_decap_8 FILLER_20_755 ();
 sg13g2_decap_8 FILLER_20_762 ();
 sg13g2_decap_8 FILLER_20_769 ();
 sg13g2_decap_8 FILLER_20_776 ();
 sg13g2_decap_8 FILLER_20_783 ();
 sg13g2_decap_8 FILLER_20_790 ();
 sg13g2_decap_8 FILLER_20_797 ();
 sg13g2_decap_8 FILLER_20_804 ();
 sg13g2_decap_8 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_20_825 ();
 sg13g2_decap_8 FILLER_20_832 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_decap_4 FILLER_21_97 ();
 sg13g2_decap_8 FILLER_21_124 ();
 sg13g2_decap_8 FILLER_21_131 ();
 sg13g2_decap_4 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_142 ();
 sg13g2_decap_4 FILLER_21_155 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_decap_4 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_decap_4 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_4 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_fill_1 FILLER_21_371 ();
 sg13g2_decap_4 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_2 FILLER_21_444 ();
 sg13g2_fill_1 FILLER_21_446 ();
 sg13g2_fill_2 FILLER_21_496 ();
 sg13g2_fill_1 FILLER_21_498 ();
 sg13g2_fill_1 FILLER_21_513 ();
 sg13g2_fill_2 FILLER_21_529 ();
 sg13g2_fill_1 FILLER_21_531 ();
 sg13g2_fill_2 FILLER_21_567 ();
 sg13g2_fill_1 FILLER_21_569 ();
 sg13g2_fill_1 FILLER_21_596 ();
 sg13g2_decap_8 FILLER_21_600 ();
 sg13g2_fill_2 FILLER_21_607 ();
 sg13g2_fill_1 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_619 ();
 sg13g2_decap_8 FILLER_21_626 ();
 sg13g2_decap_8 FILLER_21_633 ();
 sg13g2_decap_8 FILLER_21_640 ();
 sg13g2_decap_8 FILLER_21_647 ();
 sg13g2_decap_8 FILLER_21_654 ();
 sg13g2_decap_8 FILLER_21_661 ();
 sg13g2_decap_8 FILLER_21_668 ();
 sg13g2_decap_8 FILLER_21_675 ();
 sg13g2_decap_8 FILLER_21_682 ();
 sg13g2_decap_8 FILLER_21_689 ();
 sg13g2_decap_8 FILLER_21_696 ();
 sg13g2_decap_8 FILLER_21_703 ();
 sg13g2_decap_8 FILLER_21_710 ();
 sg13g2_decap_8 FILLER_21_717 ();
 sg13g2_decap_8 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_731 ();
 sg13g2_decap_8 FILLER_21_738 ();
 sg13g2_decap_8 FILLER_21_745 ();
 sg13g2_decap_8 FILLER_21_752 ();
 sg13g2_decap_8 FILLER_21_759 ();
 sg13g2_decap_8 FILLER_21_766 ();
 sg13g2_decap_8 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_780 ();
 sg13g2_decap_8 FILLER_21_787 ();
 sg13g2_decap_8 FILLER_21_794 ();
 sg13g2_decap_8 FILLER_21_801 ();
 sg13g2_decap_8 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_815 ();
 sg13g2_decap_8 FILLER_21_822 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_decap_8 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_850 ();
 sg13g2_decap_4 FILLER_21_857 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_decap_4 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_decap_4 FILLER_22_162 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_4 FILLER_22_323 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_fill_1 FILLER_22_404 ();
 sg13g2_decap_4 FILLER_22_415 ();
 sg13g2_fill_2 FILLER_22_419 ();
 sg13g2_fill_1 FILLER_22_435 ();
 sg13g2_fill_2 FILLER_22_445 ();
 sg13g2_fill_1 FILLER_22_447 ();
 sg13g2_fill_1 FILLER_22_519 ();
 sg13g2_decap_4 FILLER_22_564 ();
 sg13g2_fill_1 FILLER_22_568 ();
 sg13g2_decap_4 FILLER_22_574 ();
 sg13g2_fill_2 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_decap_8 FILLER_23_82 ();
 sg13g2_fill_2 FILLER_23_89 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_decap_4 FILLER_23_102 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_decap_4 FILLER_23_138 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_decap_4 FILLER_23_351 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_370 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_decap_4 FILLER_23_396 ();
 sg13g2_fill_1 FILLER_23_400 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_fill_2 FILLER_23_430 ();
 sg13g2_fill_1 FILLER_23_432 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_fill_2 FILLER_23_462 ();
 sg13g2_decap_4 FILLER_23_518 ();
 sg13g2_fill_2 FILLER_23_531 ();
 sg13g2_fill_1 FILLER_23_533 ();
 sg13g2_decap_8 FILLER_23_578 ();
 sg13g2_fill_1 FILLER_23_585 ();
 sg13g2_fill_2 FILLER_23_609 ();
 sg13g2_fill_1 FILLER_23_642 ();
 sg13g2_decap_8 FILLER_23_652 ();
 sg13g2_decap_8 FILLER_23_659 ();
 sg13g2_decap_8 FILLER_23_666 ();
 sg13g2_decap_8 FILLER_23_673 ();
 sg13g2_decap_8 FILLER_23_680 ();
 sg13g2_decap_8 FILLER_23_687 ();
 sg13g2_decap_8 FILLER_23_694 ();
 sg13g2_decap_8 FILLER_23_701 ();
 sg13g2_decap_8 FILLER_23_708 ();
 sg13g2_decap_8 FILLER_23_715 ();
 sg13g2_decap_8 FILLER_23_722 ();
 sg13g2_decap_8 FILLER_23_729 ();
 sg13g2_decap_8 FILLER_23_736 ();
 sg13g2_decap_8 FILLER_23_743 ();
 sg13g2_decap_8 FILLER_23_750 ();
 sg13g2_decap_8 FILLER_23_757 ();
 sg13g2_decap_8 FILLER_23_764 ();
 sg13g2_decap_8 FILLER_23_771 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_8 FILLER_23_785 ();
 sg13g2_decap_8 FILLER_23_792 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_decap_8 FILLER_23_820 ();
 sg13g2_decap_8 FILLER_23_827 ();
 sg13g2_decap_8 FILLER_23_834 ();
 sg13g2_decap_8 FILLER_23_841 ();
 sg13g2_decap_8 FILLER_23_848 ();
 sg13g2_decap_8 FILLER_23_855 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_fill_2 FILLER_24_59 ();
 sg13g2_fill_1 FILLER_24_61 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_1 FILLER_24_89 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_decap_4 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_decap_4 FILLER_24_155 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_214 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_decap_4 FILLER_24_318 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_decap_4 FILLER_24_331 ();
 sg13g2_fill_2 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_4 FILLER_24_349 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_decap_4 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_449 ();
 sg13g2_fill_1 FILLER_24_456 ();
 sg13g2_fill_2 FILLER_24_471 ();
 sg13g2_decap_4 FILLER_24_517 ();
 sg13g2_fill_1 FILLER_24_529 ();
 sg13g2_decap_4 FILLER_24_563 ();
 sg13g2_fill_2 FILLER_24_626 ();
 sg13g2_fill_1 FILLER_24_628 ();
 sg13g2_decap_8 FILLER_24_655 ();
 sg13g2_decap_8 FILLER_24_662 ();
 sg13g2_decap_8 FILLER_24_669 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_690 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_704 ();
 sg13g2_decap_8 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_718 ();
 sg13g2_decap_8 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_8 FILLER_24_746 ();
 sg13g2_decap_8 FILLER_24_753 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_decap_8 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_decap_8 FILLER_24_788 ();
 sg13g2_decap_8 FILLER_24_795 ();
 sg13g2_decap_8 FILLER_24_802 ();
 sg13g2_decap_8 FILLER_24_809 ();
 sg13g2_decap_8 FILLER_24_816 ();
 sg13g2_decap_8 FILLER_24_823 ();
 sg13g2_decap_8 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_837 ();
 sg13g2_decap_8 FILLER_24_844 ();
 sg13g2_decap_8 FILLER_24_851 ();
 sg13g2_decap_4 FILLER_24_858 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_51 ();
 sg13g2_decap_8 FILLER_25_58 ();
 sg13g2_decap_8 FILLER_25_65 ();
 sg13g2_decap_4 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_decap_4 FILLER_25_90 ();
 sg13g2_fill_2 FILLER_25_94 ();
 sg13g2_decap_4 FILLER_25_101 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_decap_4 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_decap_4 FILLER_25_136 ();
 sg13g2_fill_2 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_decap_4 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_decap_4 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_4 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_fill_1 FILLER_25_390 ();
 sg13g2_decap_4 FILLER_25_415 ();
 sg13g2_fill_1 FILLER_25_419 ();
 sg13g2_fill_2 FILLER_25_435 ();
 sg13g2_fill_1 FILLER_25_437 ();
 sg13g2_decap_8 FILLER_25_443 ();
 sg13g2_fill_2 FILLER_25_450 ();
 sg13g2_fill_1 FILLER_25_452 ();
 sg13g2_decap_4 FILLER_25_488 ();
 sg13g2_fill_2 FILLER_25_518 ();
 sg13g2_fill_2 FILLER_25_595 ();
 sg13g2_fill_1 FILLER_25_597 ();
 sg13g2_decap_8 FILLER_25_603 ();
 sg13g2_decap_4 FILLER_25_610 ();
 sg13g2_fill_1 FILLER_25_614 ();
 sg13g2_fill_1 FILLER_25_627 ();
 sg13g2_decap_8 FILLER_25_654 ();
 sg13g2_decap_8 FILLER_25_661 ();
 sg13g2_decap_8 FILLER_25_668 ();
 sg13g2_decap_8 FILLER_25_675 ();
 sg13g2_decap_8 FILLER_25_682 ();
 sg13g2_decap_8 FILLER_25_689 ();
 sg13g2_decap_8 FILLER_25_696 ();
 sg13g2_decap_8 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_710 ();
 sg13g2_decap_8 FILLER_25_717 ();
 sg13g2_decap_8 FILLER_25_724 ();
 sg13g2_decap_8 FILLER_25_731 ();
 sg13g2_decap_8 FILLER_25_738 ();
 sg13g2_decap_8 FILLER_25_745 ();
 sg13g2_decap_8 FILLER_25_752 ();
 sg13g2_decap_8 FILLER_25_759 ();
 sg13g2_decap_8 FILLER_25_766 ();
 sg13g2_decap_8 FILLER_25_773 ();
 sg13g2_decap_8 FILLER_25_780 ();
 sg13g2_decap_8 FILLER_25_787 ();
 sg13g2_decap_8 FILLER_25_794 ();
 sg13g2_decap_8 FILLER_25_801 ();
 sg13g2_decap_8 FILLER_25_808 ();
 sg13g2_decap_8 FILLER_25_815 ();
 sg13g2_decap_8 FILLER_25_822 ();
 sg13g2_decap_8 FILLER_25_829 ();
 sg13g2_decap_8 FILLER_25_836 ();
 sg13g2_decap_8 FILLER_25_843 ();
 sg13g2_decap_8 FILLER_25_850 ();
 sg13g2_decap_4 FILLER_25_857 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_decap_4 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_fill_2 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_decap_8 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_299 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_4 FILLER_26_339 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_397 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_26_415 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_1 FILLER_26_449 ();
 sg13g2_decap_8 FILLER_26_459 ();
 sg13g2_fill_2 FILLER_26_466 ();
 sg13g2_decap_4 FILLER_26_487 ();
 sg13g2_fill_1 FILLER_26_491 ();
 sg13g2_fill_2 FILLER_26_534 ();
 sg13g2_fill_1 FILLER_26_536 ();
 sg13g2_decap_4 FILLER_26_582 ();
 sg13g2_fill_2 FILLER_26_586 ();
 sg13g2_fill_2 FILLER_26_638 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_fill_2 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_decap_4 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_decap_8 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_decap_4 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_216 ();
 sg13g2_decap_4 FILLER_27_233 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_346 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_2 FILLER_27_366 ();
 sg13g2_decap_4 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_400 ();
 sg13g2_fill_1 FILLER_27_402 ();
 sg13g2_decap_4 FILLER_27_412 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_fill_1 FILLER_27_430 ();
 sg13g2_fill_1 FILLER_27_511 ();
 sg13g2_fill_1 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_591 ();
 sg13g2_decap_4 FILLER_27_624 ();
 sg13g2_decap_8 FILLER_27_654 ();
 sg13g2_decap_8 FILLER_27_661 ();
 sg13g2_decap_8 FILLER_27_668 ();
 sg13g2_decap_8 FILLER_27_675 ();
 sg13g2_decap_8 FILLER_27_682 ();
 sg13g2_decap_8 FILLER_27_689 ();
 sg13g2_decap_8 FILLER_27_696 ();
 sg13g2_decap_8 FILLER_27_703 ();
 sg13g2_decap_8 FILLER_27_710 ();
 sg13g2_decap_8 FILLER_27_717 ();
 sg13g2_decap_8 FILLER_27_724 ();
 sg13g2_decap_8 FILLER_27_731 ();
 sg13g2_decap_8 FILLER_27_738 ();
 sg13g2_decap_8 FILLER_27_745 ();
 sg13g2_decap_8 FILLER_27_752 ();
 sg13g2_decap_8 FILLER_27_759 ();
 sg13g2_decap_8 FILLER_27_766 ();
 sg13g2_decap_8 FILLER_27_773 ();
 sg13g2_decap_8 FILLER_27_780 ();
 sg13g2_decap_8 FILLER_27_787 ();
 sg13g2_decap_8 FILLER_27_794 ();
 sg13g2_decap_8 FILLER_27_801 ();
 sg13g2_decap_8 FILLER_27_808 ();
 sg13g2_decap_8 FILLER_27_815 ();
 sg13g2_decap_8 FILLER_27_822 ();
 sg13g2_decap_8 FILLER_27_829 ();
 sg13g2_decap_8 FILLER_27_836 ();
 sg13g2_decap_8 FILLER_27_843 ();
 sg13g2_decap_8 FILLER_27_850 ();
 sg13g2_decap_4 FILLER_27_857 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_66 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_decap_4 FILLER_28_74 ();
 sg13g2_fill_2 FILLER_28_78 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_decap_8 FILLER_28_99 ();
 sg13g2_decap_8 FILLER_28_106 ();
 sg13g2_fill_2 FILLER_28_113 ();
 sg13g2_fill_1 FILLER_28_115 ();
 sg13g2_decap_4 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_184 ();
 sg13g2_decap_4 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_decap_4 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_28_412 ();
 sg13g2_fill_2 FILLER_28_424 ();
 sg13g2_decap_4 FILLER_28_461 ();
 sg13g2_fill_2 FILLER_28_465 ();
 sg13g2_fill_1 FILLER_28_489 ();
 sg13g2_fill_1 FILLER_28_530 ();
 sg13g2_fill_2 FILLER_28_557 ();
 sg13g2_fill_1 FILLER_28_559 ();
 sg13g2_fill_2 FILLER_28_569 ();
 sg13g2_fill_2 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_590 ();
 sg13g2_fill_2 FILLER_28_597 ();
 sg13g2_decap_8 FILLER_28_652 ();
 sg13g2_decap_8 FILLER_28_659 ();
 sg13g2_decap_8 FILLER_28_666 ();
 sg13g2_decap_8 FILLER_28_673 ();
 sg13g2_decap_8 FILLER_28_680 ();
 sg13g2_decap_8 FILLER_28_687 ();
 sg13g2_decap_8 FILLER_28_694 ();
 sg13g2_decap_8 FILLER_28_701 ();
 sg13g2_decap_8 FILLER_28_708 ();
 sg13g2_decap_8 FILLER_28_715 ();
 sg13g2_decap_8 FILLER_28_722 ();
 sg13g2_decap_8 FILLER_28_729 ();
 sg13g2_decap_8 FILLER_28_736 ();
 sg13g2_decap_8 FILLER_28_743 ();
 sg13g2_decap_8 FILLER_28_750 ();
 sg13g2_decap_8 FILLER_28_757 ();
 sg13g2_decap_8 FILLER_28_764 ();
 sg13g2_decap_8 FILLER_28_771 ();
 sg13g2_decap_8 FILLER_28_778 ();
 sg13g2_decap_8 FILLER_28_785 ();
 sg13g2_decap_8 FILLER_28_792 ();
 sg13g2_decap_8 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_806 ();
 sg13g2_decap_8 FILLER_28_813 ();
 sg13g2_decap_8 FILLER_28_820 ();
 sg13g2_decap_8 FILLER_28_827 ();
 sg13g2_decap_8 FILLER_28_834 ();
 sg13g2_decap_8 FILLER_28_841 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_fill_2 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_decap_4 FILLER_29_127 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_fill_2 FILLER_29_378 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_422 ();
 sg13g2_fill_1 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_461 ();
 sg13g2_fill_2 FILLER_29_498 ();
 sg13g2_fill_1 FILLER_29_500 ();
 sg13g2_fill_1 FILLER_29_510 ();
 sg13g2_fill_2 FILLER_29_529 ();
 sg13g2_decap_4 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_604 ();
 sg13g2_decap_8 FILLER_29_611 ();
 sg13g2_fill_2 FILLER_29_618 ();
 sg13g2_fill_2 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_646 ();
 sg13g2_decap_8 FILLER_29_653 ();
 sg13g2_decap_8 FILLER_29_660 ();
 sg13g2_decap_8 FILLER_29_667 ();
 sg13g2_decap_8 FILLER_29_674 ();
 sg13g2_decap_8 FILLER_29_681 ();
 sg13g2_decap_8 FILLER_29_688 ();
 sg13g2_decap_8 FILLER_29_695 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_709 ();
 sg13g2_decap_8 FILLER_29_716 ();
 sg13g2_decap_8 FILLER_29_723 ();
 sg13g2_decap_8 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_8 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_72 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_96 ();
 sg13g2_fill_2 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_110 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_decap_4 FILLER_30_128 ();
 sg13g2_decap_4 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_178 ();
 sg13g2_decap_4 FILLER_30_185 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_4 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_decap_4 FILLER_30_247 ();
 sg13g2_decap_4 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_4 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_419 ();
 sg13g2_decap_8 FILLER_30_429 ();
 sg13g2_fill_1 FILLER_30_436 ();
 sg13g2_decap_8 FILLER_30_472 ();
 sg13g2_fill_2 FILLER_30_479 ();
 sg13g2_decap_8 FILLER_30_486 ();
 sg13g2_fill_1 FILLER_30_493 ();
 sg13g2_fill_2 FILLER_30_538 ();
 sg13g2_fill_2 FILLER_30_544 ();
 sg13g2_fill_2 FILLER_30_555 ();
 sg13g2_fill_1 FILLER_30_557 ();
 sg13g2_fill_2 FILLER_30_580 ();
 sg13g2_fill_1 FILLER_30_582 ();
 sg13g2_fill_2 FILLER_30_644 ();
 sg13g2_fill_1 FILLER_30_646 ();
 sg13g2_decap_8 FILLER_30_673 ();
 sg13g2_fill_1 FILLER_30_680 ();
 sg13g2_fill_2 FILLER_30_685 ();
 sg13g2_fill_1 FILLER_30_687 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_44 ();
 sg13g2_fill_2 FILLER_31_50 ();
 sg13g2_fill_1 FILLER_31_52 ();
 sg13g2_decap_4 FILLER_31_57 ();
 sg13g2_decap_8 FILLER_31_66 ();
 sg13g2_decap_4 FILLER_31_73 ();
 sg13g2_decap_8 FILLER_31_82 ();
 sg13g2_fill_2 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_4 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_345 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_4 FILLER_31_415 ();
 sg13g2_fill_1 FILLER_31_424 ();
 sg13g2_fill_2 FILLER_31_433 ();
 sg13g2_decap_8 FILLER_31_487 ();
 sg13g2_decap_4 FILLER_31_494 ();
 sg13g2_fill_2 FILLER_31_504 ();
 sg13g2_fill_2 FILLER_31_526 ();
 sg13g2_fill_1 FILLER_31_528 ();
 sg13g2_fill_2 FILLER_31_555 ();
 sg13g2_fill_1 FILLER_31_557 ();
 sg13g2_fill_2 FILLER_31_571 ();
 sg13g2_fill_1 FILLER_31_573 ();
 sg13g2_fill_1 FILLER_31_595 ();
 sg13g2_fill_2 FILLER_31_618 ();
 sg13g2_fill_1 FILLER_31_620 ();
 sg13g2_decap_4 FILLER_31_655 ();
 sg13g2_fill_2 FILLER_31_659 ();
 sg13g2_fill_2 FILLER_31_702 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_fill_1 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_741 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_decap_8 FILLER_31_769 ();
 sg13g2_decap_8 FILLER_31_776 ();
 sg13g2_decap_8 FILLER_31_783 ();
 sg13g2_decap_8 FILLER_31_790 ();
 sg13g2_decap_8 FILLER_31_797 ();
 sg13g2_decap_8 FILLER_31_804 ();
 sg13g2_decap_8 FILLER_31_811 ();
 sg13g2_decap_8 FILLER_31_818 ();
 sg13g2_decap_8 FILLER_31_825 ();
 sg13g2_decap_8 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_decap_8 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_853 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_87 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_4 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_221 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_308 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_decap_8 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_32_440 ();
 sg13g2_decap_8 FILLER_32_447 ();
 sg13g2_decap_8 FILLER_32_454 ();
 sg13g2_decap_8 FILLER_32_461 ();
 sg13g2_decap_4 FILLER_32_468 ();
 sg13g2_fill_2 FILLER_32_472 ();
 sg13g2_fill_2 FILLER_32_526 ();
 sg13g2_fill_1 FILLER_32_528 ();
 sg13g2_fill_1 FILLER_32_546 ();
 sg13g2_fill_2 FILLER_32_562 ();
 sg13g2_decap_8 FILLER_32_591 ();
 sg13g2_decap_8 FILLER_32_598 ();
 sg13g2_decap_8 FILLER_32_605 ();
 sg13g2_decap_8 FILLER_32_612 ();
 sg13g2_fill_2 FILLER_32_619 ();
 sg13g2_fill_1 FILLER_32_621 ();
 sg13g2_fill_1 FILLER_32_640 ();
 sg13g2_decap_8 FILLER_32_662 ();
 sg13g2_fill_2 FILLER_32_669 ();
 sg13g2_decap_4 FILLER_32_680 ();
 sg13g2_fill_1 FILLER_32_684 ();
 sg13g2_decap_4 FILLER_32_689 ();
 sg13g2_fill_1 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_746 ();
 sg13g2_decap_8 FILLER_32_753 ();
 sg13g2_decap_8 FILLER_32_760 ();
 sg13g2_decap_8 FILLER_32_767 ();
 sg13g2_decap_8 FILLER_32_774 ();
 sg13g2_decap_8 FILLER_32_781 ();
 sg13g2_decap_8 FILLER_32_788 ();
 sg13g2_decap_8 FILLER_32_795 ();
 sg13g2_decap_8 FILLER_32_802 ();
 sg13g2_decap_8 FILLER_32_809 ();
 sg13g2_decap_8 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_823 ();
 sg13g2_decap_8 FILLER_32_830 ();
 sg13g2_decap_8 FILLER_32_837 ();
 sg13g2_decap_8 FILLER_32_844 ();
 sg13g2_decap_8 FILLER_32_851 ();
 sg13g2_decap_4 FILLER_32_858 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_decap_4 FILLER_33_68 ();
 sg13g2_fill_2 FILLER_33_72 ();
 sg13g2_decap_8 FILLER_33_96 ();
 sg13g2_decap_8 FILLER_33_103 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_181 ();
 sg13g2_decap_8 FILLER_33_188 ();
 sg13g2_decap_4 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_205 ();
 sg13g2_decap_4 FILLER_33_221 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_decap_4 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_290 ();
 sg13g2_decap_4 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_33_416 ();
 sg13g2_fill_1 FILLER_33_428 ();
 sg13g2_fill_2 FILLER_33_432 ();
 sg13g2_fill_1 FILLER_33_434 ();
 sg13g2_fill_1 FILLER_33_440 ();
 sg13g2_fill_2 FILLER_33_454 ();
 sg13g2_fill_1 FILLER_33_456 ();
 sg13g2_fill_2 FILLER_33_470 ();
 sg13g2_fill_1 FILLER_33_472 ();
 sg13g2_fill_2 FILLER_33_544 ();
 sg13g2_fill_1 FILLER_33_546 ();
 sg13g2_decap_4 FILLER_33_626 ();
 sg13g2_decap_8 FILLER_33_639 ();
 sg13g2_fill_1 FILLER_33_646 ();
 sg13g2_decap_8 FILLER_33_652 ();
 sg13g2_fill_2 FILLER_33_659 ();
 sg13g2_fill_1 FILLER_33_666 ();
 sg13g2_fill_1 FILLER_33_685 ();
 sg13g2_fill_1 FILLER_33_705 ();
 sg13g2_fill_2 FILLER_33_712 ();
 sg13g2_fill_2 FILLER_33_723 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_8 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_decap_8 FILLER_33_781 ();
 sg13g2_decap_8 FILLER_33_788 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_decap_8 FILLER_33_816 ();
 sg13g2_decap_8 FILLER_33_823 ();
 sg13g2_decap_8 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_837 ();
 sg13g2_decap_8 FILLER_33_844 ();
 sg13g2_decap_8 FILLER_33_851 ();
 sg13g2_decap_4 FILLER_33_858 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_18 ();
 sg13g2_fill_2 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_86 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_4 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_159 ();
 sg13g2_decap_4 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_fill_2 FILLER_34_176 ();
 sg13g2_fill_1 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_fill_1 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_decap_4 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_34_412 ();
 sg13g2_fill_2 FILLER_34_446 ();
 sg13g2_fill_2 FILLER_34_468 ();
 sg13g2_decap_4 FILLER_34_486 ();
 sg13g2_decap_4 FILLER_34_527 ();
 sg13g2_fill_1 FILLER_34_531 ();
 sg13g2_decap_8 FILLER_34_537 ();
 sg13g2_decap_4 FILLER_34_544 ();
 sg13g2_decap_4 FILLER_34_556 ();
 sg13g2_fill_2 FILLER_34_594 ();
 sg13g2_fill_2 FILLER_34_605 ();
 sg13g2_decap_4 FILLER_34_647 ();
 sg13g2_fill_2 FILLER_34_651 ();
 sg13g2_decap_4 FILLER_34_662 ();
 sg13g2_decap_4 FILLER_34_671 ();
 sg13g2_decap_4 FILLER_34_688 ();
 sg13g2_fill_1 FILLER_34_692 ();
 sg13g2_fill_2 FILLER_34_736 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_fill_2 FILLER_35_97 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_decap_4 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_decap_8 FILLER_35_293 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_decap_8 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_decap_4 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_decap_4 FILLER_35_358 ();
 sg13g2_fill_2 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_35_432 ();
 sg13g2_decap_4 FILLER_35_438 ();
 sg13g2_fill_1 FILLER_35_442 ();
 sg13g2_decap_4 FILLER_35_456 ();
 sg13g2_fill_2 FILLER_35_460 ();
 sg13g2_fill_2 FILLER_35_479 ();
 sg13g2_fill_2 FILLER_35_522 ();
 sg13g2_fill_1 FILLER_35_558 ();
 sg13g2_decap_8 FILLER_35_585 ();
 sg13g2_decap_4 FILLER_35_592 ();
 sg13g2_fill_2 FILLER_35_618 ();
 sg13g2_decap_8 FILLER_35_632 ();
 sg13g2_decap_4 FILLER_35_639 ();
 sg13g2_decap_4 FILLER_35_695 ();
 sg13g2_fill_1 FILLER_35_699 ();
 sg13g2_decap_8 FILLER_35_711 ();
 sg13g2_fill_2 FILLER_35_718 ();
 sg13g2_decap_4 FILLER_35_729 ();
 sg13g2_fill_2 FILLER_35_733 ();
 sg13g2_fill_1 FILLER_35_738 ();
 sg13g2_fill_1 FILLER_35_755 ();
 sg13g2_decap_8 FILLER_35_769 ();
 sg13g2_decap_8 FILLER_35_776 ();
 sg13g2_decap_8 FILLER_35_783 ();
 sg13g2_decap_8 FILLER_35_790 ();
 sg13g2_decap_8 FILLER_35_797 ();
 sg13g2_decap_8 FILLER_35_804 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_decap_8 FILLER_35_832 ();
 sg13g2_decap_8 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_846 ();
 sg13g2_decap_8 FILLER_35_853 ();
 sg13g2_fill_2 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_66 ();
 sg13g2_fill_1 FILLER_36_89 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_136 ();
 sg13g2_decap_8 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_decap_8 FILLER_36_173 ();
 sg13g2_decap_4 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_decap_8 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_decap_4 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_decap_4 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_fill_1 FILLER_36_367 ();
 sg13g2_fill_1 FILLER_36_402 ();
 sg13g2_decap_4 FILLER_36_407 ();
 sg13g2_fill_2 FILLER_36_411 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_decap_8 FILLER_36_430 ();
 sg13g2_decap_4 FILLER_36_437 ();
 sg13g2_fill_1 FILLER_36_467 ();
 sg13g2_decap_8 FILLER_36_487 ();
 sg13g2_decap_4 FILLER_36_494 ();
 sg13g2_decap_4 FILLER_36_503 ();
 sg13g2_decap_4 FILLER_36_520 ();
 sg13g2_fill_1 FILLER_36_528 ();
 sg13g2_decap_8 FILLER_36_548 ();
 sg13g2_decap_4 FILLER_36_555 ();
 sg13g2_fill_2 FILLER_36_559 ();
 sg13g2_decap_4 FILLER_36_580 ();
 sg13g2_fill_2 FILLER_36_592 ();
 sg13g2_fill_2 FILLER_36_607 ();
 sg13g2_fill_1 FILLER_36_609 ();
 sg13g2_decap_4 FILLER_36_637 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_decap_4 FILLER_36_650 ();
 sg13g2_fill_2 FILLER_36_654 ();
 sg13g2_decap_8 FILLER_36_661 ();
 sg13g2_decap_8 FILLER_36_668 ();
 sg13g2_decap_8 FILLER_36_675 ();
 sg13g2_decap_8 FILLER_36_682 ();
 sg13g2_decap_4 FILLER_36_689 ();
 sg13g2_decap_4 FILLER_36_744 ();
 sg13g2_decap_8 FILLER_36_774 ();
 sg13g2_decap_8 FILLER_36_781 ();
 sg13g2_decap_8 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_decap_8 FILLER_36_830 ();
 sg13g2_decap_8 FILLER_36_837 ();
 sg13g2_decap_8 FILLER_36_844 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_decap_4 FILLER_36_858 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_88 ();
 sg13g2_decap_4 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_106 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_decap_4 FILLER_37_230 ();
 sg13g2_decap_4 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_261 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_decap_4 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_decap_4 FILLER_37_371 ();
 sg13g2_fill_2 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_433 ();
 sg13g2_fill_2 FILLER_37_440 ();
 sg13g2_decap_8 FILLER_37_450 ();
 sg13g2_fill_1 FILLER_37_457 ();
 sg13g2_fill_1 FILLER_37_467 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_fill_2 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_513 ();
 sg13g2_decap_8 FILLER_37_520 ();
 sg13g2_decap_8 FILLER_37_540 ();
 sg13g2_fill_2 FILLER_37_547 ();
 sg13g2_fill_1 FILLER_37_554 ();
 sg13g2_fill_1 FILLER_37_570 ();
 sg13g2_decap_4 FILLER_37_587 ();
 sg13g2_decap_8 FILLER_37_603 ();
 sg13g2_decap_4 FILLER_37_610 ();
 sg13g2_fill_2 FILLER_37_614 ();
 sg13g2_decap_8 FILLER_37_632 ();
 sg13g2_decap_4 FILLER_37_647 ();
 sg13g2_fill_1 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_687 ();
 sg13g2_decap_8 FILLER_37_694 ();
 sg13g2_decap_8 FILLER_37_710 ();
 sg13g2_decap_4 FILLER_37_717 ();
 sg13g2_fill_2 FILLER_37_721 ();
 sg13g2_fill_2 FILLER_37_727 ();
 sg13g2_fill_1 FILLER_37_729 ();
 sg13g2_fill_2 FILLER_37_743 ();
 sg13g2_decap_4 FILLER_37_759 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_fill_1 FILLER_38_67 ();
 sg13g2_decap_4 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_fill_1 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_4 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_253 ();
 sg13g2_decap_4 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_decap_4 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_298 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_decap_4 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_decap_4 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_418 ();
 sg13g2_decap_8 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_432 ();
 sg13g2_decap_8 FILLER_38_449 ();
 sg13g2_decap_4 FILLER_38_456 ();
 sg13g2_fill_2 FILLER_38_460 ();
 sg13g2_fill_2 FILLER_38_493 ();
 sg13g2_fill_1 FILLER_38_495 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_fill_1 FILLER_38_511 ();
 sg13g2_fill_2 FILLER_38_527 ();
 sg13g2_decap_8 FILLER_38_564 ();
 sg13g2_decap_8 FILLER_38_607 ();
 sg13g2_fill_2 FILLER_38_614 ();
 sg13g2_fill_1 FILLER_38_633 ();
 sg13g2_decap_8 FILLER_38_650 ();
 sg13g2_decap_8 FILLER_38_657 ();
 sg13g2_decap_4 FILLER_38_664 ();
 sg13g2_fill_2 FILLER_38_692 ();
 sg13g2_decap_4 FILLER_38_715 ();
 sg13g2_fill_1 FILLER_38_719 ();
 sg13g2_decap_8 FILLER_38_724 ();
 sg13g2_fill_1 FILLER_38_731 ();
 sg13g2_fill_2 FILLER_38_737 ();
 sg13g2_fill_2 FILLER_38_756 ();
 sg13g2_fill_1 FILLER_38_758 ();
 sg13g2_decap_8 FILLER_38_785 ();
 sg13g2_decap_8 FILLER_38_792 ();
 sg13g2_decap_8 FILLER_38_799 ();
 sg13g2_decap_8 FILLER_38_806 ();
 sg13g2_decap_8 FILLER_38_813 ();
 sg13g2_decap_8 FILLER_38_820 ();
 sg13g2_decap_8 FILLER_38_827 ();
 sg13g2_decap_8 FILLER_38_834 ();
 sg13g2_decap_8 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_848 ();
 sg13g2_decap_8 FILLER_38_855 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_4 FILLER_39_42 ();
 sg13g2_fill_2 FILLER_39_46 ();
 sg13g2_fill_2 FILLER_39_58 ();
 sg13g2_decap_8 FILLER_39_86 ();
 sg13g2_decap_4 FILLER_39_93 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_146 ();
 sg13g2_fill_1 FILLER_39_148 ();
 sg13g2_fill_1 FILLER_39_154 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_decap_4 FILLER_39_192 ();
 sg13g2_fill_1 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_204 ();
 sg13g2_decap_8 FILLER_39_211 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_235 ();
 sg13g2_decap_4 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_245 ();
 sg13g2_fill_2 FILLER_39_273 ();
 sg13g2_fill_1 FILLER_39_275 ();
 sg13g2_fill_2 FILLER_39_305 ();
 sg13g2_decap_8 FILLER_39_323 ();
 sg13g2_decap_8 FILLER_39_351 ();
 sg13g2_fill_2 FILLER_39_358 ();
 sg13g2_decap_8 FILLER_39_370 ();
 sg13g2_fill_2 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_388 ();
 sg13g2_decap_4 FILLER_39_395 ();
 sg13g2_fill_2 FILLER_39_402 ();
 sg13g2_fill_1 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_409 ();
 sg13g2_decap_4 FILLER_39_415 ();
 sg13g2_fill_2 FILLER_39_419 ();
 sg13g2_decap_8 FILLER_39_459 ();
 sg13g2_decap_4 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_486 ();
 sg13g2_fill_2 FILLER_39_493 ();
 sg13g2_decap_4 FILLER_39_508 ();
 sg13g2_fill_2 FILLER_39_520 ();
 sg13g2_fill_2 FILLER_39_530 ();
 sg13g2_fill_1 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_560 ();
 sg13g2_fill_2 FILLER_39_567 ();
 sg13g2_fill_2 FILLER_39_577 ();
 sg13g2_fill_1 FILLER_39_579 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_fill_1 FILLER_39_600 ();
 sg13g2_fill_1 FILLER_39_618 ();
 sg13g2_fill_1 FILLER_39_641 ();
 sg13g2_decap_8 FILLER_39_668 ();
 sg13g2_fill_1 FILLER_39_675 ();
 sg13g2_fill_1 FILLER_39_680 ();
 sg13g2_decap_4 FILLER_39_735 ();
 sg13g2_fill_1 FILLER_39_739 ();
 sg13g2_decap_4 FILLER_39_764 ();
 sg13g2_fill_2 FILLER_39_768 ();
 sg13g2_decap_8 FILLER_39_774 ();
 sg13g2_decap_8 FILLER_39_781 ();
 sg13g2_decap_8 FILLER_39_788 ();
 sg13g2_decap_8 FILLER_39_795 ();
 sg13g2_decap_8 FILLER_39_802 ();
 sg13g2_decap_8 FILLER_39_809 ();
 sg13g2_decap_8 FILLER_39_816 ();
 sg13g2_decap_8 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_830 ();
 sg13g2_decap_8 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_4 FILLER_39_858 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_decap_8 FILLER_40_43 ();
 sg13g2_decap_8 FILLER_40_50 ();
 sg13g2_decap_4 FILLER_40_57 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_decap_4 FILLER_40_79 ();
 sg13g2_fill_2 FILLER_40_83 ();
 sg13g2_fill_2 FILLER_40_120 ();
 sg13g2_fill_1 FILLER_40_122 ();
 sg13g2_fill_1 FILLER_40_144 ();
 sg13g2_decap_8 FILLER_40_170 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_decap_8 FILLER_40_186 ();
 sg13g2_decap_4 FILLER_40_193 ();
 sg13g2_fill_1 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_202 ();
 sg13g2_fill_2 FILLER_40_222 ();
 sg13g2_decap_8 FILLER_40_229 ();
 sg13g2_decap_8 FILLER_40_236 ();
 sg13g2_fill_1 FILLER_40_243 ();
 sg13g2_fill_2 FILLER_40_249 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_fill_2 FILLER_40_287 ();
 sg13g2_fill_1 FILLER_40_289 ();
 sg13g2_fill_2 FILLER_40_294 ();
 sg13g2_fill_2 FILLER_40_313 ();
 sg13g2_decap_8 FILLER_40_323 ();
 sg13g2_decap_4 FILLER_40_330 ();
 sg13g2_fill_2 FILLER_40_334 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_fill_1 FILLER_40_419 ();
 sg13g2_fill_2 FILLER_40_425 ();
 sg13g2_fill_1 FILLER_40_427 ();
 sg13g2_fill_2 FILLER_40_458 ();
 sg13g2_decap_8 FILLER_40_477 ();
 sg13g2_decap_4 FILLER_40_484 ();
 sg13g2_fill_1 FILLER_40_488 ();
 sg13g2_fill_1 FILLER_40_519 ();
 sg13g2_fill_2 FILLER_40_536 ();
 sg13g2_fill_2 FILLER_40_576 ();
 sg13g2_fill_1 FILLER_40_578 ();
 sg13g2_decap_8 FILLER_40_659 ();
 sg13g2_fill_1 FILLER_40_671 ();
 sg13g2_fill_2 FILLER_40_688 ();
 sg13g2_fill_1 FILLER_40_690 ();
 sg13g2_decap_8 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_fill_2 FILLER_40_730 ();
 sg13g2_decap_8 FILLER_40_753 ();
 sg13g2_fill_1 FILLER_40_760 ();
 sg13g2_decap_8 FILLER_40_774 ();
 sg13g2_decap_8 FILLER_40_781 ();
 sg13g2_decap_8 FILLER_40_788 ();
 sg13g2_decap_8 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_802 ();
 sg13g2_decap_8 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_decap_8 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_16 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_fill_2 FILLER_41_28 ();
 sg13g2_fill_1 FILLER_41_30 ();
 sg13g2_fill_2 FILLER_41_65 ();
 sg13g2_fill_1 FILLER_41_76 ();
 sg13g2_decap_4 FILLER_41_125 ();
 sg13g2_decap_4 FILLER_41_132 ();
 sg13g2_decap_8 FILLER_41_141 ();
 sg13g2_fill_2 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_150 ();
 sg13g2_decap_8 FILLER_41_156 ();
 sg13g2_decap_8 FILLER_41_163 ();
 sg13g2_decap_4 FILLER_41_170 ();
 sg13g2_fill_2 FILLER_41_174 ();
 sg13g2_fill_1 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_fill_2 FILLER_41_224 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_decap_4 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_263 ();
 sg13g2_fill_2 FILLER_41_299 ();
 sg13g2_fill_1 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_fill_2 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_fill_2 FILLER_41_359 ();
 sg13g2_fill_1 FILLER_41_361 ();
 sg13g2_decap_8 FILLER_41_375 ();
 sg13g2_decap_8 FILLER_41_382 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_fill_1 FILLER_41_396 ();
 sg13g2_fill_2 FILLER_41_405 ();
 sg13g2_fill_1 FILLER_41_407 ();
 sg13g2_fill_2 FILLER_41_416 ();
 sg13g2_decap_8 FILLER_41_444 ();
 sg13g2_decap_8 FILLER_41_451 ();
 sg13g2_decap_8 FILLER_41_458 ();
 sg13g2_fill_1 FILLER_41_465 ();
 sg13g2_decap_4 FILLER_41_492 ();
 sg13g2_decap_8 FILLER_41_512 ();
 sg13g2_decap_4 FILLER_41_519 ();
 sg13g2_decap_8 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_535 ();
 sg13g2_decap_8 FILLER_41_550 ();
 sg13g2_decap_8 FILLER_41_557 ();
 sg13g2_decap_4 FILLER_41_564 ();
 sg13g2_fill_1 FILLER_41_568 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_fill_2 FILLER_41_602 ();
 sg13g2_fill_1 FILLER_41_604 ();
 sg13g2_fill_2 FILLER_41_614 ();
 sg13g2_fill_2 FILLER_41_621 ();
 sg13g2_fill_2 FILLER_41_645 ();
 sg13g2_fill_1 FILLER_41_647 ();
 sg13g2_fill_2 FILLER_41_666 ();
 sg13g2_decap_4 FILLER_41_677 ();
 sg13g2_fill_2 FILLER_41_681 ();
 sg13g2_fill_2 FILLER_41_746 ();
 sg13g2_fill_2 FILLER_41_753 ();
 sg13g2_fill_1 FILLER_41_755 ();
 sg13g2_decap_8 FILLER_41_782 ();
 sg13g2_decap_8 FILLER_41_789 ();
 sg13g2_decap_8 FILLER_41_796 ();
 sg13g2_decap_8 FILLER_41_803 ();
 sg13g2_decap_8 FILLER_41_810 ();
 sg13g2_decap_8 FILLER_41_817 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_8 FILLER_41_831 ();
 sg13g2_decap_8 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_fill_2 FILLER_41_859 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_4 ();
 sg13g2_decap_8 FILLER_42_32 ();
 sg13g2_fill_2 FILLER_42_39 ();
 sg13g2_fill_1 FILLER_42_41 ();
 sg13g2_fill_1 FILLER_42_46 ();
 sg13g2_decap_4 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_69 ();
 sg13g2_fill_1 FILLER_42_79 ();
 sg13g2_decap_4 FILLER_42_88 ();
 sg13g2_fill_2 FILLER_42_92 ();
 sg13g2_decap_4 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_102 ();
 sg13g2_decap_8 FILLER_42_122 ();
 sg13g2_fill_1 FILLER_42_129 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_fill_2 FILLER_42_174 ();
 sg13g2_decap_8 FILLER_42_194 ();
 sg13g2_decap_4 FILLER_42_201 ();
 sg13g2_fill_2 FILLER_42_205 ();
 sg13g2_fill_1 FILLER_42_220 ();
 sg13g2_fill_2 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_4 FILLER_42_259 ();
 sg13g2_fill_2 FILLER_42_263 ();
 sg13g2_fill_2 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_290 ();
 sg13g2_fill_1 FILLER_42_292 ();
 sg13g2_fill_2 FILLER_42_301 ();
 sg13g2_fill_1 FILLER_42_318 ();
 sg13g2_decap_4 FILLER_42_324 ();
 sg13g2_fill_2 FILLER_42_328 ();
 sg13g2_fill_2 FILLER_42_335 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_356 ();
 sg13g2_fill_1 FILLER_42_358 ();
 sg13g2_decap_4 FILLER_42_363 ();
 sg13g2_fill_1 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_4 FILLER_42_401 ();
 sg13g2_fill_2 FILLER_42_405 ();
 sg13g2_fill_1 FILLER_42_415 ();
 sg13g2_decap_8 FILLER_42_437 ();
 sg13g2_fill_2 FILLER_42_444 ();
 sg13g2_fill_1 FILLER_42_446 ();
 sg13g2_fill_2 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_4 FILLER_42_483 ();
 sg13g2_fill_2 FILLER_42_487 ();
 sg13g2_fill_2 FILLER_42_531 ();
 sg13g2_fill_1 FILLER_42_533 ();
 sg13g2_fill_2 FILLER_42_549 ();
 sg13g2_fill_1 FILLER_42_551 ();
 sg13g2_decap_4 FILLER_42_578 ();
 sg13g2_fill_2 FILLER_42_582 ();
 sg13g2_fill_1 FILLER_42_615 ();
 sg13g2_fill_2 FILLER_42_641 ();
 sg13g2_fill_1 FILLER_42_643 ();
 sg13g2_decap_4 FILLER_42_648 ();
 sg13g2_fill_2 FILLER_42_652 ();
 sg13g2_decap_4 FILLER_42_659 ();
 sg13g2_fill_1 FILLER_42_663 ();
 sg13g2_decap_8 FILLER_42_690 ();
 sg13g2_fill_1 FILLER_42_702 ();
 sg13g2_fill_2 FILLER_42_715 ();
 sg13g2_fill_1 FILLER_42_717 ();
 sg13g2_fill_2 FILLER_42_727 ();
 sg13g2_fill_1 FILLER_42_729 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_4 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_4 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_27 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_fill_2 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_55 ();
 sg13g2_fill_2 FILLER_43_67 ();
 sg13g2_fill_1 FILLER_43_69 ();
 sg13g2_fill_1 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_4 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_109 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_4 FILLER_43_126 ();
 sg13g2_fill_1 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_144 ();
 sg13g2_decap_8 FILLER_43_150 ();
 sg13g2_fill_2 FILLER_43_157 ();
 sg13g2_decap_4 FILLER_43_163 ();
 sg13g2_decap_8 FILLER_43_171 ();
 sg13g2_fill_2 FILLER_43_178 ();
 sg13g2_fill_1 FILLER_43_180 ();
 sg13g2_decap_8 FILLER_43_211 ();
 sg13g2_decap_8 FILLER_43_218 ();
 sg13g2_fill_1 FILLER_43_225 ();
 sg13g2_decap_8 FILLER_43_230 ();
 sg13g2_fill_2 FILLER_43_237 ();
 sg13g2_decap_4 FILLER_43_249 ();
 sg13g2_fill_1 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_290 ();
 sg13g2_decap_4 FILLER_43_326 ();
 sg13g2_fill_1 FILLER_43_330 ();
 sg13g2_decap_8 FILLER_43_339 ();
 sg13g2_fill_2 FILLER_43_346 ();
 sg13g2_fill_1 FILLER_43_348 ();
 sg13g2_decap_4 FILLER_43_357 ();
 sg13g2_fill_1 FILLER_43_372 ();
 sg13g2_decap_4 FILLER_43_382 ();
 sg13g2_fill_2 FILLER_43_398 ();
 sg13g2_fill_1 FILLER_43_400 ();
 sg13g2_decap_4 FILLER_43_408 ();
 sg13g2_decap_4 FILLER_43_443 ();
 sg13g2_fill_1 FILLER_43_447 ();
 sg13g2_fill_2 FILLER_43_465 ();
 sg13g2_decap_4 FILLER_43_493 ();
 sg13g2_fill_1 FILLER_43_497 ();
 sg13g2_fill_2 FILLER_43_515 ();
 sg13g2_decap_4 FILLER_43_539 ();
 sg13g2_fill_1 FILLER_43_543 ();
 sg13g2_decap_8 FILLER_43_556 ();
 sg13g2_fill_2 FILLER_43_567 ();
 sg13g2_fill_1 FILLER_43_569 ();
 sg13g2_decap_8 FILLER_43_604 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_628 ();
 sg13g2_decap_4 FILLER_43_635 ();
 sg13g2_fill_2 FILLER_43_639 ();
 sg13g2_fill_1 FILLER_43_646 ();
 sg13g2_decap_8 FILLER_43_667 ();
 sg13g2_fill_1 FILLER_43_674 ();
 sg13g2_decap_8 FILLER_43_684 ();
 sg13g2_fill_2 FILLER_43_703 ();
 sg13g2_fill_1 FILLER_43_722 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_4 ();
 sg13g2_fill_1 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_123 ();
 sg13g2_fill_1 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_171 ();
 sg13g2_fill_2 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_185 ();
 sg13g2_fill_2 FILLER_44_195 ();
 sg13g2_fill_1 FILLER_44_197 ();
 sg13g2_fill_2 FILLER_44_203 ();
 sg13g2_fill_1 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_223 ();
 sg13g2_decap_8 FILLER_44_251 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_fill_2 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_fill_2 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_4 FILLER_44_301 ();
 sg13g2_fill_1 FILLER_44_318 ();
 sg13g2_decap_4 FILLER_44_324 ();
 sg13g2_decap_8 FILLER_44_339 ();
 sg13g2_decap_4 FILLER_44_360 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_4 FILLER_44_389 ();
 sg13g2_fill_2 FILLER_44_393 ();
 sg13g2_fill_2 FILLER_44_416 ();
 sg13g2_fill_1 FILLER_44_418 ();
 sg13g2_fill_1 FILLER_44_447 ();
 sg13g2_decap_4 FILLER_44_473 ();
 sg13g2_fill_1 FILLER_44_477 ();
 sg13g2_decap_8 FILLER_44_482 ();
 sg13g2_fill_2 FILLER_44_489 ();
 sg13g2_fill_1 FILLER_44_491 ();
 sg13g2_decap_8 FILLER_44_514 ();
 sg13g2_fill_2 FILLER_44_521 ();
 sg13g2_fill_1 FILLER_44_523 ();
 sg13g2_decap_8 FILLER_44_538 ();
 sg13g2_fill_2 FILLER_44_545 ();
 sg13g2_fill_1 FILLER_44_547 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_8 FILLER_44_567 ();
 sg13g2_fill_1 FILLER_44_574 ();
 sg13g2_fill_1 FILLER_44_583 ();
 sg13g2_decap_4 FILLER_44_601 ();
 sg13g2_fill_1 FILLER_44_605 ();
 sg13g2_fill_1 FILLER_44_615 ();
 sg13g2_fill_1 FILLER_44_619 ();
 sg13g2_fill_1 FILLER_44_651 ();
 sg13g2_fill_1 FILLER_44_656 ();
 sg13g2_fill_2 FILLER_44_699 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_11 ();
 sg13g2_fill_2 FILLER_45_29 ();
 sg13g2_fill_1 FILLER_45_61 ();
 sg13g2_decap_8 FILLER_45_100 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_fill_1 FILLER_45_109 ();
 sg13g2_decap_8 FILLER_45_124 ();
 sg13g2_fill_2 FILLER_45_131 ();
 sg13g2_decap_8 FILLER_45_139 ();
 sg13g2_decap_4 FILLER_45_146 ();
 sg13g2_decap_4 FILLER_45_155 ();
 sg13g2_fill_1 FILLER_45_159 ();
 sg13g2_fill_1 FILLER_45_167 ();
 sg13g2_decap_4 FILLER_45_173 ();
 sg13g2_decap_8 FILLER_45_199 ();
 sg13g2_decap_8 FILLER_45_206 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_236 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_fill_2 FILLER_45_249 ();
 sg13g2_fill_1 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_296 ();
 sg13g2_decap_8 FILLER_45_304 ();
 sg13g2_fill_1 FILLER_45_311 ();
 sg13g2_decap_8 FILLER_45_316 ();
 sg13g2_fill_2 FILLER_45_323 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_fill_2 FILLER_45_336 ();
 sg13g2_fill_1 FILLER_45_338 ();
 sg13g2_fill_2 FILLER_45_359 ();
 sg13g2_fill_2 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_402 ();
 sg13g2_fill_2 FILLER_45_436 ();
 sg13g2_decap_8 FILLER_45_465 ();
 sg13g2_decap_8 FILLER_45_477 ();
 sg13g2_decap_4 FILLER_45_484 ();
 sg13g2_decap_4 FILLER_45_509 ();
 sg13g2_fill_1 FILLER_45_513 ();
 sg13g2_fill_2 FILLER_45_522 ();
 sg13g2_fill_2 FILLER_45_543 ();
 sg13g2_fill_1 FILLER_45_545 ();
 sg13g2_fill_2 FILLER_45_563 ();
 sg13g2_fill_1 FILLER_45_565 ();
 sg13g2_decap_8 FILLER_45_573 ();
 sg13g2_decap_4 FILLER_45_585 ();
 sg13g2_fill_2 FILLER_45_589 ();
 sg13g2_decap_8 FILLER_45_617 ();
 sg13g2_decap_8 FILLER_45_662 ();
 sg13g2_decap_8 FILLER_45_669 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_decap_4 FILLER_45_683 ();
 sg13g2_fill_2 FILLER_45_692 ();
 sg13g2_fill_1 FILLER_45_694 ();
 sg13g2_decap_8 FILLER_45_702 ();
 sg13g2_fill_1 FILLER_45_709 ();
 sg13g2_decap_8 FILLER_45_719 ();
 sg13g2_decap_8 FILLER_45_726 ();
 sg13g2_decap_8 FILLER_45_733 ();
 sg13g2_decap_8 FILLER_45_740 ();
 sg13g2_decap_8 FILLER_45_747 ();
 sg13g2_decap_8 FILLER_45_754 ();
 sg13g2_decap_8 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_768 ();
 sg13g2_decap_8 FILLER_45_775 ();
 sg13g2_decap_8 FILLER_45_782 ();
 sg13g2_decap_8 FILLER_45_789 ();
 sg13g2_decap_8 FILLER_45_796 ();
 sg13g2_decap_8 FILLER_45_803 ();
 sg13g2_decap_8 FILLER_45_810 ();
 sg13g2_decap_8 FILLER_45_817 ();
 sg13g2_decap_8 FILLER_45_824 ();
 sg13g2_decap_8 FILLER_45_831 ();
 sg13g2_decap_8 FILLER_45_838 ();
 sg13g2_decap_8 FILLER_45_845 ();
 sg13g2_decap_8 FILLER_45_852 ();
 sg13g2_fill_2 FILLER_45_859 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_1 FILLER_46_29 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_92 ();
 sg13g2_decap_4 FILLER_46_115 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_fill_2 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_135 ();
 sg13g2_fill_2 FILLER_46_149 ();
 sg13g2_fill_1 FILLER_46_151 ();
 sg13g2_fill_2 FILLER_46_160 ();
 sg13g2_fill_1 FILLER_46_167 ();
 sg13g2_decap_8 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_190 ();
 sg13g2_decap_8 FILLER_46_207 ();
 sg13g2_decap_8 FILLER_46_214 ();
 sg13g2_decap_4 FILLER_46_247 ();
 sg13g2_fill_2 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_271 ();
 sg13g2_fill_1 FILLER_46_273 ();
 sg13g2_fill_2 FILLER_46_283 ();
 sg13g2_fill_2 FILLER_46_290 ();
 sg13g2_fill_1 FILLER_46_292 ();
 sg13g2_decap_4 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_306 ();
 sg13g2_fill_2 FILLER_46_321 ();
 sg13g2_fill_1 FILLER_46_323 ();
 sg13g2_decap_8 FILLER_46_333 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_345 ();
 sg13g2_decap_8 FILLER_46_351 ();
 sg13g2_fill_2 FILLER_46_366 ();
 sg13g2_fill_1 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_fill_2 FILLER_46_403 ();
 sg13g2_fill_1 FILLER_46_405 ();
 sg13g2_fill_2 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_417 ();
 sg13g2_decap_4 FILLER_46_424 ();
 sg13g2_decap_8 FILLER_46_442 ();
 sg13g2_fill_2 FILLER_46_449 ();
 sg13g2_fill_2 FILLER_46_459 ();
 sg13g2_decap_4 FILLER_46_484 ();
 sg13g2_fill_1 FILLER_46_488 ();
 sg13g2_fill_2 FILLER_46_494 ();
 sg13g2_decap_8 FILLER_46_505 ();
 sg13g2_decap_8 FILLER_46_512 ();
 sg13g2_fill_1 FILLER_46_519 ();
 sg13g2_fill_1 FILLER_46_527 ();
 sg13g2_fill_2 FILLER_46_554 ();
 sg13g2_fill_1 FILLER_46_556 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_fill_1 FILLER_46_595 ();
 sg13g2_fill_1 FILLER_46_601 ();
 sg13g2_decap_8 FILLER_46_606 ();
 sg13g2_decap_4 FILLER_46_613 ();
 sg13g2_fill_1 FILLER_46_617 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_4 FILLER_46_637 ();
 sg13g2_fill_2 FILLER_46_641 ();
 sg13g2_decap_8 FILLER_46_646 ();
 sg13g2_fill_2 FILLER_46_653 ();
 sg13g2_fill_1 FILLER_46_655 ();
 sg13g2_fill_2 FILLER_46_687 ();
 sg13g2_fill_1 FILLER_46_689 ();
 sg13g2_fill_1 FILLER_46_699 ();
 sg13g2_decap_4 FILLER_46_719 ();
 sg13g2_fill_1 FILLER_46_723 ();
 sg13g2_decap_8 FILLER_46_734 ();
 sg13g2_decap_8 FILLER_46_741 ();
 sg13g2_decap_8 FILLER_46_748 ();
 sg13g2_decap_8 FILLER_46_755 ();
 sg13g2_decap_8 FILLER_46_762 ();
 sg13g2_decap_8 FILLER_46_769 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_decap_8 FILLER_46_783 ();
 sg13g2_decap_8 FILLER_46_790 ();
 sg13g2_decap_8 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_804 ();
 sg13g2_decap_8 FILLER_46_811 ();
 sg13g2_decap_8 FILLER_46_818 ();
 sg13g2_decap_8 FILLER_46_825 ();
 sg13g2_decap_8 FILLER_46_832 ();
 sg13g2_decap_8 FILLER_46_839 ();
 sg13g2_decap_8 FILLER_46_846 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_27 ();
 sg13g2_decap_8 FILLER_47_46 ();
 sg13g2_decap_8 FILLER_47_53 ();
 sg13g2_decap_8 FILLER_47_60 ();
 sg13g2_fill_2 FILLER_47_67 ();
 sg13g2_fill_1 FILLER_47_69 ();
 sg13g2_fill_2 FILLER_47_74 ();
 sg13g2_fill_1 FILLER_47_76 ();
 sg13g2_decap_8 FILLER_47_81 ();
 sg13g2_decap_8 FILLER_47_88 ();
 sg13g2_fill_2 FILLER_47_95 ();
 sg13g2_decap_8 FILLER_47_114 ();
 sg13g2_decap_4 FILLER_47_121 ();
 sg13g2_decap_8 FILLER_47_138 ();
 sg13g2_decap_8 FILLER_47_145 ();
 sg13g2_decap_4 FILLER_47_152 ();
 sg13g2_fill_1 FILLER_47_156 ();
 sg13g2_fill_1 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_167 ();
 sg13g2_fill_2 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_184 ();
 sg13g2_fill_1 FILLER_47_191 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_206 ();
 sg13g2_decap_8 FILLER_47_213 ();
 sg13g2_fill_2 FILLER_47_220 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_decap_4 FILLER_47_281 ();
 sg13g2_fill_2 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_fill_1 FILLER_47_299 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_315 ();
 sg13g2_decap_4 FILLER_47_321 ();
 sg13g2_fill_2 FILLER_47_348 ();
 sg13g2_decap_4 FILLER_47_355 ();
 sg13g2_fill_2 FILLER_47_424 ();
 sg13g2_decap_8 FILLER_47_452 ();
 sg13g2_decap_8 FILLER_47_459 ();
 sg13g2_fill_2 FILLER_47_466 ();
 sg13g2_fill_1 FILLER_47_468 ();
 sg13g2_decap_4 FILLER_47_478 ();
 sg13g2_fill_2 FILLER_47_482 ();
 sg13g2_fill_1 FILLER_47_492 ();
 sg13g2_decap_4 FILLER_47_509 ();
 sg13g2_decap_4 FILLER_47_534 ();
 sg13g2_fill_1 FILLER_47_538 ();
 sg13g2_fill_2 FILLER_47_559 ();
 sg13g2_fill_1 FILLER_47_561 ();
 sg13g2_decap_4 FILLER_47_585 ();
 sg13g2_fill_2 FILLER_47_609 ();
 sg13g2_fill_1 FILLER_47_611 ();
 sg13g2_fill_2 FILLER_47_633 ();
 sg13g2_fill_1 FILLER_47_635 ();
 sg13g2_decap_8 FILLER_47_667 ();
 sg13g2_fill_1 FILLER_47_674 ();
 sg13g2_fill_1 FILLER_47_680 ();
 sg13g2_fill_2 FILLER_47_710 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_fill_1 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_734 ();
 sg13g2_fill_1 FILLER_47_741 ();
 sg13g2_decap_8 FILLER_47_755 ();
 sg13g2_decap_8 FILLER_47_762 ();
 sg13g2_decap_8 FILLER_47_769 ();
 sg13g2_decap_8 FILLER_47_776 ();
 sg13g2_decap_8 FILLER_47_783 ();
 sg13g2_decap_8 FILLER_47_790 ();
 sg13g2_decap_8 FILLER_47_797 ();
 sg13g2_decap_8 FILLER_47_804 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_818 ();
 sg13g2_decap_8 FILLER_47_825 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_839 ();
 sg13g2_decap_8 FILLER_47_846 ();
 sg13g2_decap_8 FILLER_47_853 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_fill_2 FILLER_48_55 ();
 sg13g2_decap_4 FILLER_48_82 ();
 sg13g2_fill_1 FILLER_48_86 ();
 sg13g2_decap_8 FILLER_48_100 ();
 sg13g2_fill_2 FILLER_48_120 ();
 sg13g2_decap_4 FILLER_48_127 ();
 sg13g2_fill_1 FILLER_48_149 ();
 sg13g2_decap_4 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_decap_4 FILLER_48_185 ();
 sg13g2_fill_1 FILLER_48_189 ();
 sg13g2_fill_2 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_202 ();
 sg13g2_decap_4 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_215 ();
 sg13g2_fill_2 FILLER_48_238 ();
 sg13g2_decap_4 FILLER_48_243 ();
 sg13g2_fill_1 FILLER_48_247 ();
 sg13g2_fill_2 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_282 ();
 sg13g2_decap_8 FILLER_48_296 ();
 sg13g2_fill_1 FILLER_48_307 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_decap_4 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_344 ();
 sg13g2_fill_2 FILLER_48_351 ();
 sg13g2_fill_1 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_362 ();
 sg13g2_fill_1 FILLER_48_364 ();
 sg13g2_decap_4 FILLER_48_395 ();
 sg13g2_fill_1 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_48_410 ();
 sg13g2_decap_4 FILLER_48_419 ();
 sg13g2_decap_8 FILLER_48_426 ();
 sg13g2_decap_4 FILLER_48_433 ();
 sg13g2_fill_2 FILLER_48_441 ();
 sg13g2_fill_1 FILLER_48_443 ();
 sg13g2_decap_8 FILLER_48_478 ();
 sg13g2_decap_8 FILLER_48_485 ();
 sg13g2_fill_2 FILLER_48_492 ();
 sg13g2_fill_1 FILLER_48_494 ();
 sg13g2_fill_2 FILLER_48_503 ();
 sg13g2_decap_8 FILLER_48_510 ();
 sg13g2_decap_8 FILLER_48_517 ();
 sg13g2_decap_8 FILLER_48_524 ();
 sg13g2_decap_4 FILLER_48_531 ();
 sg13g2_fill_2 FILLER_48_535 ();
 sg13g2_fill_2 FILLER_48_567 ();
 sg13g2_fill_1 FILLER_48_569 ();
 sg13g2_fill_2 FILLER_48_609 ();
 sg13g2_fill_2 FILLER_48_626 ();
 sg13g2_fill_1 FILLER_48_628 ();
 sg13g2_fill_1 FILLER_48_640 ();
 sg13g2_fill_2 FILLER_48_660 ();
 sg13g2_fill_1 FILLER_48_688 ();
 sg13g2_fill_2 FILLER_48_702 ();
 sg13g2_fill_1 FILLER_48_718 ();
 sg13g2_fill_1 FILLER_48_727 ();
 sg13g2_decap_8 FILLER_48_757 ();
 sg13g2_decap_8 FILLER_48_764 ();
 sg13g2_decap_8 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_792 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_decap_8 FILLER_48_813 ();
 sg13g2_decap_8 FILLER_48_820 ();
 sg13g2_decap_8 FILLER_48_827 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_841 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_49 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_2 FILLER_49_65 ();
 sg13g2_fill_1 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_72 ();
 sg13g2_decap_4 FILLER_49_79 ();
 sg13g2_fill_2 FILLER_49_108 ();
 sg13g2_decap_4 FILLER_49_131 ();
 sg13g2_decap_8 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_170 ();
 sg13g2_decap_8 FILLER_49_194 ();
 sg13g2_decap_8 FILLER_49_201 ();
 sg13g2_decap_4 FILLER_49_208 ();
 sg13g2_decap_4 FILLER_49_226 ();
 sg13g2_fill_2 FILLER_49_230 ();
 sg13g2_decap_4 FILLER_49_237 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_4 FILLER_49_291 ();
 sg13g2_fill_2 FILLER_49_303 ();
 sg13g2_fill_1 FILLER_49_305 ();
 sg13g2_fill_1 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_335 ();
 sg13g2_decap_8 FILLER_49_365 ();
 sg13g2_decap_4 FILLER_49_372 ();
 sg13g2_fill_2 FILLER_49_376 ();
 sg13g2_fill_2 FILLER_49_394 ();
 sg13g2_fill_1 FILLER_49_396 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_fill_2 FILLER_49_409 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_fill_1 FILLER_49_455 ();
 sg13g2_decap_4 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_467 ();
 sg13g2_decap_4 FILLER_49_474 ();
 sg13g2_decap_4 FILLER_49_528 ();
 sg13g2_fill_2 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_568 ();
 sg13g2_decap_4 FILLER_49_575 ();
 sg13g2_fill_2 FILLER_49_579 ();
 sg13g2_decap_4 FILLER_49_585 ();
 sg13g2_fill_2 FILLER_49_589 ();
 sg13g2_decap_4 FILLER_49_596 ();
 sg13g2_fill_1 FILLER_49_600 ();
 sg13g2_decap_4 FILLER_49_606 ();
 sg13g2_decap_4 FILLER_49_619 ();
 sg13g2_fill_1 FILLER_49_643 ();
 sg13g2_fill_2 FILLER_49_658 ();
 sg13g2_fill_1 FILLER_49_660 ();
 sg13g2_decap_8 FILLER_49_688 ();
 sg13g2_decap_4 FILLER_49_695 ();
 sg13g2_fill_1 FILLER_49_711 ();
 sg13g2_decap_8 FILLER_49_717 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_4 FILLER_49_744 ();
 sg13g2_fill_2 FILLER_49_748 ();
 sg13g2_decap_8 FILLER_49_758 ();
 sg13g2_decap_8 FILLER_49_765 ();
 sg13g2_decap_8 FILLER_49_772 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_793 ();
 sg13g2_decap_8 FILLER_49_800 ();
 sg13g2_decap_8 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_decap_8 FILLER_49_821 ();
 sg13g2_decap_8 FILLER_49_828 ();
 sg13g2_decap_8 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_4 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_18 ();
 sg13g2_decap_8 FILLER_50_41 ();
 sg13g2_decap_8 FILLER_50_48 ();
 sg13g2_fill_2 FILLER_50_55 ();
 sg13g2_fill_1 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_99 ();
 sg13g2_decap_8 FILLER_50_106 ();
 sg13g2_decap_8 FILLER_50_113 ();
 sg13g2_decap_8 FILLER_50_120 ();
 sg13g2_decap_8 FILLER_50_127 ();
 sg13g2_fill_2 FILLER_50_134 ();
 sg13g2_decap_4 FILLER_50_144 ();
 sg13g2_fill_2 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_158 ();
 sg13g2_decap_4 FILLER_50_168 ();
 sg13g2_fill_2 FILLER_50_172 ();
 sg13g2_decap_4 FILLER_50_194 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_fill_2 FILLER_50_212 ();
 sg13g2_fill_1 FILLER_50_214 ();
 sg13g2_decap_4 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_260 ();
 sg13g2_fill_2 FILLER_50_279 ();
 sg13g2_decap_4 FILLER_50_291 ();
 sg13g2_fill_1 FILLER_50_295 ();
 sg13g2_decap_8 FILLER_50_312 ();
 sg13g2_decap_4 FILLER_50_319 ();
 sg13g2_fill_2 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_334 ();
 sg13g2_fill_2 FILLER_50_344 ();
 sg13g2_fill_1 FILLER_50_346 ();
 sg13g2_fill_2 FILLER_50_356 ();
 sg13g2_decap_8 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_378 ();
 sg13g2_fill_2 FILLER_50_385 ();
 sg13g2_fill_2 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_2 FILLER_50_408 ();
 sg13g2_fill_2 FILLER_50_458 ();
 sg13g2_fill_1 FILLER_50_500 ();
 sg13g2_decap_8 FILLER_50_533 ();
 sg13g2_decap_8 FILLER_50_540 ();
 sg13g2_decap_8 FILLER_50_547 ();
 sg13g2_fill_2 FILLER_50_554 ();
 sg13g2_fill_1 FILLER_50_561 ();
 sg13g2_fill_2 FILLER_50_581 ();
 sg13g2_fill_1 FILLER_50_583 ();
 sg13g2_fill_1 FILLER_50_589 ();
 sg13g2_decap_4 FILLER_50_597 ();
 sg13g2_fill_2 FILLER_50_616 ();
 sg13g2_fill_1 FILLER_50_618 ();
 sg13g2_decap_8 FILLER_50_642 ();
 sg13g2_decap_4 FILLER_50_659 ();
 sg13g2_decap_4 FILLER_50_668 ();
 sg13g2_fill_1 FILLER_50_672 ();
 sg13g2_fill_2 FILLER_50_698 ();
 sg13g2_decap_8 FILLER_50_710 ();
 sg13g2_fill_1 FILLER_50_717 ();
 sg13g2_decap_4 FILLER_50_730 ();
 sg13g2_decap_8 FILLER_50_748 ();
 sg13g2_decap_4 FILLER_50_755 ();
 sg13g2_fill_2 FILLER_50_759 ();
 sg13g2_decap_8 FILLER_50_765 ();
 sg13g2_decap_8 FILLER_50_772 ();
 sg13g2_decap_8 FILLER_50_779 ();
 sg13g2_decap_8 FILLER_50_786 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_decap_8 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_807 ();
 sg13g2_decap_8 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_821 ();
 sg13g2_decap_8 FILLER_50_828 ();
 sg13g2_decap_8 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_842 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_36 ();
 sg13g2_fill_1 FILLER_51_51 ();
 sg13g2_decap_8 FILLER_51_65 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_decap_8 FILLER_51_79 ();
 sg13g2_decap_8 FILLER_51_94 ();
 sg13g2_decap_4 FILLER_51_101 ();
 sg13g2_fill_2 FILLER_51_105 ();
 sg13g2_fill_1 FILLER_51_191 ();
 sg13g2_fill_2 FILLER_51_201 ();
 sg13g2_fill_1 FILLER_51_203 ();
 sg13g2_decap_8 FILLER_51_212 ();
 sg13g2_decap_8 FILLER_51_240 ();
 sg13g2_fill_1 FILLER_51_247 ();
 sg13g2_fill_2 FILLER_51_274 ();
 sg13g2_decap_4 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_344 ();
 sg13g2_decap_4 FILLER_51_361 ();
 sg13g2_fill_1 FILLER_51_365 ();
 sg13g2_decap_8 FILLER_51_371 ();
 sg13g2_decap_4 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_408 ();
 sg13g2_fill_2 FILLER_51_421 ();
 sg13g2_fill_1 FILLER_51_423 ();
 sg13g2_decap_8 FILLER_51_433 ();
 sg13g2_decap_4 FILLER_51_440 ();
 sg13g2_decap_4 FILLER_51_454 ();
 sg13g2_decap_4 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_491 ();
 sg13g2_fill_1 FILLER_51_493 ();
 sg13g2_fill_1 FILLER_51_497 ();
 sg13g2_decap_8 FILLER_51_503 ();
 sg13g2_decap_4 FILLER_51_515 ();
 sg13g2_fill_1 FILLER_51_519 ();
 sg13g2_fill_1 FILLER_51_525 ();
 sg13g2_decap_8 FILLER_51_531 ();
 sg13g2_fill_2 FILLER_51_538 ();
 sg13g2_fill_1 FILLER_51_540 ();
 sg13g2_fill_2 FILLER_51_556 ();
 sg13g2_decap_8 FILLER_51_571 ();
 sg13g2_decap_8 FILLER_51_578 ();
 sg13g2_decap_8 FILLER_51_597 ();
 sg13g2_fill_1 FILLER_51_604 ();
 sg13g2_decap_4 FILLER_51_615 ();
 sg13g2_decap_8 FILLER_51_627 ();
 sg13g2_decap_8 FILLER_51_634 ();
 sg13g2_fill_1 FILLER_51_641 ();
 sg13g2_decap_8 FILLER_51_668 ();
 sg13g2_fill_2 FILLER_51_675 ();
 sg13g2_fill_1 FILLER_51_677 ();
 sg13g2_decap_8 FILLER_51_681 ();
 sg13g2_fill_1 FILLER_51_688 ();
 sg13g2_decap_8 FILLER_51_693 ();
 sg13g2_fill_2 FILLER_51_700 ();
 sg13g2_fill_1 FILLER_51_702 ();
 sg13g2_fill_2 FILLER_51_726 ();
 sg13g2_decap_8 FILLER_51_776 ();
 sg13g2_decap_8 FILLER_51_783 ();
 sg13g2_decap_8 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_797 ();
 sg13g2_decap_8 FILLER_51_804 ();
 sg13g2_decap_8 FILLER_51_811 ();
 sg13g2_decap_8 FILLER_51_818 ();
 sg13g2_decap_8 FILLER_51_825 ();
 sg13g2_decap_8 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_839 ();
 sg13g2_decap_8 FILLER_51_846 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_40 ();
 sg13g2_decap_4 FILLER_52_47 ();
 sg13g2_decap_8 FILLER_52_59 ();
 sg13g2_decap_4 FILLER_52_66 ();
 sg13g2_fill_1 FILLER_52_78 ();
 sg13g2_decap_8 FILLER_52_115 ();
 sg13g2_decap_4 FILLER_52_122 ();
 sg13g2_fill_1 FILLER_52_130 ();
 sg13g2_decap_8 FILLER_52_149 ();
 sg13g2_decap_8 FILLER_52_156 ();
 sg13g2_decap_8 FILLER_52_163 ();
 sg13g2_decap_8 FILLER_52_170 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_2 FILLER_52_197 ();
 sg13g2_fill_1 FILLER_52_199 ();
 sg13g2_decap_8 FILLER_52_209 ();
 sg13g2_decap_4 FILLER_52_216 ();
 sg13g2_fill_1 FILLER_52_225 ();
 sg13g2_decap_8 FILLER_52_230 ();
 sg13g2_decap_4 FILLER_52_237 ();
 sg13g2_fill_2 FILLER_52_241 ();
 sg13g2_decap_8 FILLER_52_282 ();
 sg13g2_decap_8 FILLER_52_289 ();
 sg13g2_decap_8 FILLER_52_296 ();
 sg13g2_decap_8 FILLER_52_303 ();
 sg13g2_fill_1 FILLER_52_310 ();
 sg13g2_decap_8 FILLER_52_327 ();
 sg13g2_fill_2 FILLER_52_334 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_345 ();
 sg13g2_decap_8 FILLER_52_352 ();
 sg13g2_decap_4 FILLER_52_374 ();
 sg13g2_fill_2 FILLER_52_378 ();
 sg13g2_fill_1 FILLER_52_393 ();
 sg13g2_fill_2 FILLER_52_445 ();
 sg13g2_fill_2 FILLER_52_466 ();
 sg13g2_fill_1 FILLER_52_468 ();
 sg13g2_decap_4 FILLER_52_521 ();
 sg13g2_fill_1 FILLER_52_525 ();
 sg13g2_fill_2 FILLER_52_538 ();
 sg13g2_decap_4 FILLER_52_553 ();
 sg13g2_fill_1 FILLER_52_557 ();
 sg13g2_decap_8 FILLER_52_563 ();
 sg13g2_fill_1 FILLER_52_575 ();
 sg13g2_decap_4 FILLER_52_588 ();
 sg13g2_decap_8 FILLER_52_604 ();
 sg13g2_decap_8 FILLER_52_624 ();
 sg13g2_fill_1 FILLER_52_631 ();
 sg13g2_fill_2 FILLER_52_637 ();
 sg13g2_fill_1 FILLER_52_639 ();
 sg13g2_decap_4 FILLER_52_649 ();
 sg13g2_decap_4 FILLER_52_657 ();
 sg13g2_fill_2 FILLER_52_661 ();
 sg13g2_decap_8 FILLER_52_675 ();
 sg13g2_fill_2 FILLER_52_682 ();
 sg13g2_fill_1 FILLER_52_684 ();
 sg13g2_decap_8 FILLER_52_700 ();
 sg13g2_fill_1 FILLER_52_707 ();
 sg13g2_decap_8 FILLER_52_721 ();
 sg13g2_fill_1 FILLER_52_728 ();
 sg13g2_fill_2 FILLER_52_750 ();
 sg13g2_fill_2 FILLER_52_755 ();
 sg13g2_decap_8 FILLER_52_762 ();
 sg13g2_decap_4 FILLER_52_769 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_decap_8 FILLER_52_791 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_1 FILLER_53_21 ();
 sg13g2_fill_1 FILLER_53_34 ();
 sg13g2_fill_1 FILLER_53_51 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_4 FILLER_53_76 ();
 sg13g2_fill_2 FILLER_53_93 ();
 sg13g2_fill_1 FILLER_53_95 ();
 sg13g2_fill_1 FILLER_53_110 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_fill_2 FILLER_53_247 ();
 sg13g2_fill_1 FILLER_53_249 ();
 sg13g2_fill_1 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_335 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_357 ();
 sg13g2_fill_2 FILLER_53_376 ();
 sg13g2_fill_1 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_8 FILLER_53_406 ();
 sg13g2_decap_8 FILLER_53_417 ();
 sg13g2_decap_4 FILLER_53_424 ();
 sg13g2_fill_2 FILLER_53_436 ();
 sg13g2_fill_1 FILLER_53_438 ();
 sg13g2_decap_4 FILLER_53_453 ();
 sg13g2_fill_1 FILLER_53_465 ();
 sg13g2_fill_2 FILLER_53_492 ();
 sg13g2_fill_2 FILLER_53_510 ();
 sg13g2_decap_4 FILLER_53_526 ();
 sg13g2_fill_2 FILLER_53_530 ();
 sg13g2_fill_2 FILLER_53_550 ();
 sg13g2_decap_4 FILLER_53_565 ();
 sg13g2_decap_8 FILLER_53_585 ();
 sg13g2_decap_8 FILLER_53_592 ();
 sg13g2_fill_2 FILLER_53_599 ();
 sg13g2_fill_1 FILLER_53_601 ();
 sg13g2_fill_1 FILLER_53_620 ();
 sg13g2_decap_8 FILLER_53_642 ();
 sg13g2_fill_1 FILLER_53_657 ();
 sg13g2_decap_4 FILLER_53_671 ();
 sg13g2_fill_2 FILLER_53_675 ();
 sg13g2_fill_2 FILLER_53_690 ();
 sg13g2_fill_1 FILLER_53_692 ();
 sg13g2_decap_8 FILLER_53_701 ();
 sg13g2_decap_8 FILLER_53_708 ();
 sg13g2_decap_4 FILLER_53_715 ();
 sg13g2_fill_2 FILLER_53_732 ();
 sg13g2_decap_8 FILLER_53_788 ();
 sg13g2_decap_8 FILLER_53_795 ();
 sg13g2_decap_8 FILLER_53_802 ();
 sg13g2_decap_8 FILLER_53_809 ();
 sg13g2_decap_8 FILLER_53_816 ();
 sg13g2_decap_8 FILLER_53_823 ();
 sg13g2_decap_8 FILLER_53_830 ();
 sg13g2_decap_8 FILLER_53_837 ();
 sg13g2_decap_8 FILLER_53_844 ();
 sg13g2_decap_8 FILLER_53_851 ();
 sg13g2_decap_4 FILLER_53_858 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_4 FILLER_54_14 ();
 sg13g2_fill_1 FILLER_54_18 ();
 sg13g2_decap_8 FILLER_54_27 ();
 sg13g2_decap_8 FILLER_54_34 ();
 sg13g2_decap_8 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_48 ();
 sg13g2_fill_1 FILLER_54_50 ();
 sg13g2_decap_8 FILLER_54_65 ();
 sg13g2_decap_4 FILLER_54_114 ();
 sg13g2_fill_2 FILLER_54_118 ();
 sg13g2_fill_1 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_155 ();
 sg13g2_decap_8 FILLER_54_162 ();
 sg13g2_decap_8 FILLER_54_174 ();
 sg13g2_fill_2 FILLER_54_181 ();
 sg13g2_fill_1 FILLER_54_183 ();
 sg13g2_decap_4 FILLER_54_209 ();
 sg13g2_fill_2 FILLER_54_213 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_decap_8 FILLER_54_226 ();
 sg13g2_decap_4 FILLER_54_233 ();
 sg13g2_fill_1 FILLER_54_237 ();
 sg13g2_decap_8 FILLER_54_251 ();
 sg13g2_decap_8 FILLER_54_258 ();
 sg13g2_decap_8 FILLER_54_265 ();
 sg13g2_decap_8 FILLER_54_272 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_fill_1 FILLER_54_281 ();
 sg13g2_fill_2 FILLER_54_295 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_fill_2 FILLER_54_339 ();
 sg13g2_fill_1 FILLER_54_341 ();
 sg13g2_decap_8 FILLER_54_347 ();
 sg13g2_fill_2 FILLER_54_354 ();
 sg13g2_fill_1 FILLER_54_356 ();
 sg13g2_fill_1 FILLER_54_363 ();
 sg13g2_decap_8 FILLER_54_368 ();
 sg13g2_decap_8 FILLER_54_375 ();
 sg13g2_decap_8 FILLER_54_382 ();
 sg13g2_fill_1 FILLER_54_389 ();
 sg13g2_fill_1 FILLER_54_406 ();
 sg13g2_fill_2 FILLER_54_421 ();
 sg13g2_decap_4 FILLER_54_442 ();
 sg13g2_fill_1 FILLER_54_446 ();
 sg13g2_decap_4 FILLER_54_456 ();
 sg13g2_fill_2 FILLER_54_460 ();
 sg13g2_decap_8 FILLER_54_501 ();
 sg13g2_fill_1 FILLER_54_508 ();
 sg13g2_decap_8 FILLER_54_525 ();
 sg13g2_decap_8 FILLER_54_532 ();
 sg13g2_decap_8 FILLER_54_539 ();
 sg13g2_fill_2 FILLER_54_546 ();
 sg13g2_fill_1 FILLER_54_548 ();
 sg13g2_decap_4 FILLER_54_554 ();
 sg13g2_fill_2 FILLER_54_563 ();
 sg13g2_fill_1 FILLER_54_565 ();
 sg13g2_decap_8 FILLER_54_574 ();
 sg13g2_decap_4 FILLER_54_581 ();
 sg13g2_decap_8 FILLER_54_602 ();
 sg13g2_fill_1 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_627 ();
 sg13g2_decap_8 FILLER_54_634 ();
 sg13g2_fill_2 FILLER_54_641 ();
 sg13g2_fill_2 FILLER_54_648 ();
 sg13g2_fill_1 FILLER_54_650 ();
 sg13g2_fill_1 FILLER_54_656 ();
 sg13g2_decap_8 FILLER_54_665 ();
 sg13g2_fill_2 FILLER_54_684 ();
 sg13g2_decap_4 FILLER_54_703 ();
 sg13g2_fill_2 FILLER_54_707 ();
 sg13g2_decap_4 FILLER_54_722 ();
 sg13g2_fill_2 FILLER_54_726 ();
 sg13g2_decap_8 FILLER_54_740 ();
 sg13g2_decap_4 FILLER_54_747 ();
 sg13g2_fill_1 FILLER_54_751 ();
 sg13g2_decap_8 FILLER_54_764 ();
 sg13g2_decap_8 FILLER_54_771 ();
 sg13g2_decap_8 FILLER_54_778 ();
 sg13g2_decap_8 FILLER_54_785 ();
 sg13g2_decap_8 FILLER_54_792 ();
 sg13g2_decap_8 FILLER_54_799 ();
 sg13g2_decap_8 FILLER_54_806 ();
 sg13g2_decap_8 FILLER_54_813 ();
 sg13g2_decap_8 FILLER_54_820 ();
 sg13g2_decap_8 FILLER_54_827 ();
 sg13g2_decap_8 FILLER_54_834 ();
 sg13g2_decap_8 FILLER_54_841 ();
 sg13g2_decap_8 FILLER_54_848 ();
 sg13g2_decap_8 FILLER_54_855 ();
 sg13g2_fill_2 FILLER_55_38 ();
 sg13g2_fill_2 FILLER_55_45 ();
 sg13g2_fill_1 FILLER_55_47 ();
 sg13g2_fill_2 FILLER_55_96 ();
 sg13g2_fill_1 FILLER_55_98 ();
 sg13g2_decap_4 FILLER_55_114 ();
 sg13g2_decap_4 FILLER_55_140 ();
 sg13g2_fill_1 FILLER_55_144 ();
 sg13g2_decap_8 FILLER_55_179 ();
 sg13g2_decap_8 FILLER_55_199 ();
 sg13g2_decap_4 FILLER_55_206 ();
 sg13g2_fill_2 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_226 ();
 sg13g2_fill_2 FILLER_55_262 ();
 sg13g2_fill_1 FILLER_55_307 ();
 sg13g2_decap_8 FILLER_55_313 ();
 sg13g2_fill_1 FILLER_55_329 ();
 sg13g2_decap_4 FILLER_55_359 ();
 sg13g2_fill_1 FILLER_55_363 ();
 sg13g2_decap_4 FILLER_55_378 ();
 sg13g2_fill_2 FILLER_55_382 ();
 sg13g2_fill_2 FILLER_55_392 ();
 sg13g2_fill_1 FILLER_55_394 ();
 sg13g2_fill_2 FILLER_55_399 ();
 sg13g2_fill_1 FILLER_55_401 ();
 sg13g2_decap_4 FILLER_55_411 ();
 sg13g2_fill_2 FILLER_55_415 ();
 sg13g2_fill_2 FILLER_55_440 ();
 sg13g2_fill_1 FILLER_55_450 ();
 sg13g2_decap_8 FILLER_55_464 ();
 sg13g2_fill_2 FILLER_55_471 ();
 sg13g2_decap_8 FILLER_55_477 ();
 sg13g2_fill_2 FILLER_55_484 ();
 sg13g2_fill_2 FILLER_55_516 ();
 sg13g2_fill_1 FILLER_55_558 ();
 sg13g2_fill_1 FILLER_55_579 ();
 sg13g2_decap_4 FILLER_55_593 ();
 sg13g2_fill_2 FILLER_55_597 ();
 sg13g2_fill_2 FILLER_55_603 ();
 sg13g2_fill_2 FILLER_55_612 ();
 sg13g2_fill_1 FILLER_55_614 ();
 sg13g2_decap_8 FILLER_55_619 ();
 sg13g2_fill_1 FILLER_55_634 ();
 sg13g2_decap_8 FILLER_55_660 ();
 sg13g2_decap_4 FILLER_55_667 ();
 sg13g2_decap_8 FILLER_55_692 ();
 sg13g2_decap_8 FILLER_55_699 ();
 sg13g2_fill_1 FILLER_55_706 ();
 sg13g2_decap_4 FILLER_55_711 ();
 sg13g2_fill_1 FILLER_55_715 ();
 sg13g2_decap_4 FILLER_55_734 ();
 sg13g2_decap_8 FILLER_55_747 ();
 sg13g2_fill_2 FILLER_55_754 ();
 sg13g2_decap_8 FILLER_55_794 ();
 sg13g2_decap_8 FILLER_55_801 ();
 sg13g2_decap_8 FILLER_55_808 ();
 sg13g2_decap_8 FILLER_55_815 ();
 sg13g2_decap_8 FILLER_55_822 ();
 sg13g2_decap_8 FILLER_55_829 ();
 sg13g2_decap_8 FILLER_55_836 ();
 sg13g2_decap_8 FILLER_55_843 ();
 sg13g2_decap_8 FILLER_55_850 ();
 sg13g2_decap_4 FILLER_55_857 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_11 ();
 sg13g2_fill_2 FILLER_56_30 ();
 sg13g2_fill_2 FILLER_56_47 ();
 sg13g2_decap_8 FILLER_56_62 ();
 sg13g2_decap_8 FILLER_56_69 ();
 sg13g2_decap_8 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_83 ();
 sg13g2_decap_8 FILLER_56_115 ();
 sg13g2_fill_1 FILLER_56_122 ();
 sg13g2_fill_1 FILLER_56_131 ();
 sg13g2_decap_4 FILLER_56_137 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_decap_8 FILLER_56_146 ();
 sg13g2_decap_8 FILLER_56_153 ();
 sg13g2_decap_8 FILLER_56_160 ();
 sg13g2_decap_4 FILLER_56_167 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_decap_8 FILLER_56_177 ();
 sg13g2_fill_2 FILLER_56_184 ();
 sg13g2_fill_1 FILLER_56_186 ();
 sg13g2_decap_4 FILLER_56_191 ();
 sg13g2_fill_2 FILLER_56_195 ();
 sg13g2_fill_1 FILLER_56_205 ();
 sg13g2_decap_8 FILLER_56_218 ();
 sg13g2_decap_8 FILLER_56_233 ();
 sg13g2_decap_4 FILLER_56_240 ();
 sg13g2_decap_4 FILLER_56_247 ();
 sg13g2_fill_2 FILLER_56_251 ();
 sg13g2_fill_2 FILLER_56_257 ();
 sg13g2_decap_8 FILLER_56_288 ();
 sg13g2_fill_2 FILLER_56_295 ();
 sg13g2_fill_2 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_309 ();
 sg13g2_fill_2 FILLER_56_321 ();
 sg13g2_decap_8 FILLER_56_334 ();
 sg13g2_decap_8 FILLER_56_341 ();
 sg13g2_decap_4 FILLER_56_348 ();
 sg13g2_fill_2 FILLER_56_352 ();
 sg13g2_fill_1 FILLER_56_372 ();
 sg13g2_fill_1 FILLER_56_382 ();
 sg13g2_fill_2 FILLER_56_391 ();
 sg13g2_fill_1 FILLER_56_393 ();
 sg13g2_decap_8 FILLER_56_418 ();
 sg13g2_fill_1 FILLER_56_425 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_441 ();
 sg13g2_decap_8 FILLER_56_472 ();
 sg13g2_decap_4 FILLER_56_479 ();
 sg13g2_fill_2 FILLER_56_483 ();
 sg13g2_decap_8 FILLER_56_489 ();
 sg13g2_fill_1 FILLER_56_496 ();
 sg13g2_fill_2 FILLER_56_501 ();
 sg13g2_fill_2 FILLER_56_512 ();
 sg13g2_decap_8 FILLER_56_524 ();
 sg13g2_decap_8 FILLER_56_531 ();
 sg13g2_decap_8 FILLER_56_542 ();
 sg13g2_decap_8 FILLER_56_549 ();
 sg13g2_decap_4 FILLER_56_556 ();
 sg13g2_decap_8 FILLER_56_598 ();
 sg13g2_decap_4 FILLER_56_605 ();
 sg13g2_fill_2 FILLER_56_627 ();
 sg13g2_fill_1 FILLER_56_642 ();
 sg13g2_decap_4 FILLER_56_647 ();
 sg13g2_decap_8 FILLER_56_659 ();
 sg13g2_fill_2 FILLER_56_666 ();
 sg13g2_fill_1 FILLER_56_668 ();
 sg13g2_decap_8 FILLER_56_685 ();
 sg13g2_fill_1 FILLER_56_692 ();
 sg13g2_decap_4 FILLER_56_702 ();
 sg13g2_decap_8 FILLER_56_718 ();
 sg13g2_fill_2 FILLER_56_725 ();
 sg13g2_fill_2 FILLER_56_743 ();
 sg13g2_decap_4 FILLER_56_770 ();
 sg13g2_fill_2 FILLER_56_774 ();
 sg13g2_decap_8 FILLER_56_800 ();
 sg13g2_decap_8 FILLER_56_807 ();
 sg13g2_decap_8 FILLER_56_814 ();
 sg13g2_decap_8 FILLER_56_821 ();
 sg13g2_decap_8 FILLER_56_828 ();
 sg13g2_decap_8 FILLER_56_835 ();
 sg13g2_decap_8 FILLER_56_842 ();
 sg13g2_decap_8 FILLER_56_849 ();
 sg13g2_decap_4 FILLER_56_856 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_fill_2 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_58 ();
 sg13g2_decap_4 FILLER_57_82 ();
 sg13g2_decap_8 FILLER_57_104 ();
 sg13g2_fill_2 FILLER_57_111 ();
 sg13g2_fill_2 FILLER_57_122 ();
 sg13g2_fill_1 FILLER_57_124 ();
 sg13g2_fill_2 FILLER_57_134 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_fill_2 FILLER_57_168 ();
 sg13g2_fill_2 FILLER_57_178 ();
 sg13g2_decap_8 FILLER_57_193 ();
 sg13g2_decap_8 FILLER_57_213 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_2 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_236 ();
 sg13g2_decap_4 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_253 ();
 sg13g2_fill_1 FILLER_57_257 ();
 sg13g2_decap_8 FILLER_57_263 ();
 sg13g2_decap_4 FILLER_57_270 ();
 sg13g2_fill_2 FILLER_57_274 ();
 sg13g2_fill_2 FILLER_57_311 ();
 sg13g2_fill_2 FILLER_57_318 ();
 sg13g2_fill_1 FILLER_57_334 ();
 sg13g2_decap_8 FILLER_57_347 ();
 sg13g2_decap_4 FILLER_57_359 ();
 sg13g2_fill_1 FILLER_57_363 ();
 sg13g2_decap_8 FILLER_57_369 ();
 sg13g2_decap_8 FILLER_57_376 ();
 sg13g2_decap_4 FILLER_57_383 ();
 sg13g2_decap_8 FILLER_57_391 ();
 sg13g2_decap_4 FILLER_57_398 ();
 sg13g2_decap_8 FILLER_57_415 ();
 sg13g2_decap_8 FILLER_57_445 ();
 sg13g2_decap_8 FILLER_57_452 ();
 sg13g2_decap_4 FILLER_57_459 ();
 sg13g2_fill_1 FILLER_57_463 ();
 sg13g2_decap_8 FILLER_57_500 ();
 sg13g2_fill_2 FILLER_57_526 ();
 sg13g2_fill_1 FILLER_57_528 ();
 sg13g2_decap_4 FILLER_57_542 ();
 sg13g2_fill_1 FILLER_57_546 ();
 sg13g2_fill_1 FILLER_57_559 ();
 sg13g2_decap_4 FILLER_57_586 ();
 sg13g2_fill_1 FILLER_57_628 ();
 sg13g2_fill_2 FILLER_57_637 ();
 sg13g2_fill_1 FILLER_57_639 ();
 sg13g2_fill_2 FILLER_57_653 ();
 sg13g2_fill_1 FILLER_57_655 ();
 sg13g2_decap_4 FILLER_57_664 ();
 sg13g2_decap_8 FILLER_57_676 ();
 sg13g2_decap_4 FILLER_57_683 ();
 sg13g2_fill_2 FILLER_57_705 ();
 sg13g2_decap_4 FILLER_57_715 ();
 sg13g2_decap_4 FILLER_57_732 ();
 sg13g2_fill_1 FILLER_57_736 ();
 sg13g2_decap_8 FILLER_57_742 ();
 sg13g2_decap_4 FILLER_57_749 ();
 sg13g2_fill_1 FILLER_57_753 ();
 sg13g2_fill_2 FILLER_57_763 ();
 sg13g2_fill_1 FILLER_57_765 ();
 sg13g2_decap_8 FILLER_57_775 ();
 sg13g2_decap_8 FILLER_57_782 ();
 sg13g2_decap_8 FILLER_57_789 ();
 sg13g2_decap_8 FILLER_57_796 ();
 sg13g2_decap_8 FILLER_57_803 ();
 sg13g2_decap_8 FILLER_57_810 ();
 sg13g2_decap_8 FILLER_57_817 ();
 sg13g2_decap_8 FILLER_57_824 ();
 sg13g2_decap_8 FILLER_57_831 ();
 sg13g2_decap_8 FILLER_57_838 ();
 sg13g2_decap_8 FILLER_57_845 ();
 sg13g2_decap_8 FILLER_57_852 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_fill_2 FILLER_58_40 ();
 sg13g2_fill_1 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_72 ();
 sg13g2_decap_4 FILLER_58_78 ();
 sg13g2_decap_4 FILLER_58_87 ();
 sg13g2_fill_1 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_100 ();
 sg13g2_decap_4 FILLER_58_107 ();
 sg13g2_fill_1 FILLER_58_111 ();
 sg13g2_fill_1 FILLER_58_125 ();
 sg13g2_decap_8 FILLER_58_139 ();
 sg13g2_decap_4 FILLER_58_146 ();
 sg13g2_fill_2 FILLER_58_150 ();
 sg13g2_decap_4 FILLER_58_155 ();
 sg13g2_decap_4 FILLER_58_178 ();
 sg13g2_fill_1 FILLER_58_182 ();
 sg13g2_fill_2 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_215 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_fill_1 FILLER_58_239 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_fill_1 FILLER_58_318 ();
 sg13g2_fill_1 FILLER_58_380 ();
 sg13g2_fill_2 FILLER_58_399 ();
 sg13g2_fill_1 FILLER_58_401 ();
 sg13g2_decap_4 FILLER_58_411 ();
 sg13g2_fill_2 FILLER_58_415 ();
 sg13g2_decap_4 FILLER_58_426 ();
 sg13g2_fill_1 FILLER_58_430 ();
 sg13g2_decap_4 FILLER_58_444 ();
 sg13g2_fill_1 FILLER_58_448 ();
 sg13g2_decap_8 FILLER_58_470 ();
 sg13g2_decap_8 FILLER_58_477 ();
 sg13g2_fill_1 FILLER_58_484 ();
 sg13g2_fill_2 FILLER_58_511 ();
 sg13g2_decap_4 FILLER_58_523 ();
 sg13g2_fill_1 FILLER_58_553 ();
 sg13g2_decap_8 FILLER_58_563 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_decap_4 FILLER_58_581 ();
 sg13g2_fill_1 FILLER_58_585 ();
 sg13g2_decap_8 FILLER_58_594 ();
 sg13g2_decap_4 FILLER_58_601 ();
 sg13g2_decap_8 FILLER_58_617 ();
 sg13g2_fill_2 FILLER_58_624 ();
 sg13g2_decap_8 FILLER_58_630 ();
 sg13g2_decap_8 FILLER_58_637 ();
 sg13g2_decap_4 FILLER_58_644 ();
 sg13g2_fill_1 FILLER_58_648 ();
 sg13g2_decap_8 FILLER_58_655 ();
 sg13g2_decap_4 FILLER_58_677 ();
 sg13g2_fill_1 FILLER_58_681 ();
 sg13g2_fill_2 FILLER_58_703 ();
 sg13g2_decap_8 FILLER_58_717 ();
 sg13g2_decap_4 FILLER_58_724 ();
 sg13g2_fill_2 FILLER_58_728 ();
 sg13g2_fill_2 FILLER_58_753 ();
 sg13g2_fill_1 FILLER_58_755 ();
 sg13g2_decap_8 FILLER_58_793 ();
 sg13g2_decap_8 FILLER_58_800 ();
 sg13g2_decap_8 FILLER_58_807 ();
 sg13g2_decap_8 FILLER_58_814 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_fill_1 FILLER_59_21 ();
 sg13g2_fill_1 FILLER_59_82 ();
 sg13g2_decap_8 FILLER_59_116 ();
 sg13g2_fill_1 FILLER_59_123 ();
 sg13g2_decap_4 FILLER_59_131 ();
 sg13g2_decap_4 FILLER_59_142 ();
 sg13g2_decap_8 FILLER_59_163 ();
 sg13g2_decap_8 FILLER_59_170 ();
 sg13g2_fill_2 FILLER_59_177 ();
 sg13g2_fill_1 FILLER_59_179 ();
 sg13g2_decap_8 FILLER_59_185 ();
 sg13g2_decap_8 FILLER_59_192 ();
 sg13g2_fill_2 FILLER_59_199 ();
 sg13g2_decap_4 FILLER_59_221 ();
 sg13g2_fill_2 FILLER_59_225 ();
 sg13g2_decap_8 FILLER_59_250 ();
 sg13g2_fill_2 FILLER_59_257 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_269 ();
 sg13g2_fill_1 FILLER_59_276 ();
 sg13g2_fill_2 FILLER_59_289 ();
 sg13g2_fill_1 FILLER_59_300 ();
 sg13g2_fill_2 FILLER_59_351 ();
 sg13g2_fill_1 FILLER_59_353 ();
 sg13g2_fill_2 FILLER_59_384 ();
 sg13g2_fill_1 FILLER_59_457 ();
 sg13g2_fill_1 FILLER_59_463 ();
 sg13g2_fill_2 FILLER_59_469 ();
 sg13g2_fill_1 FILLER_59_471 ();
 sg13g2_decap_8 FILLER_59_477 ();
 sg13g2_fill_2 FILLER_59_484 ();
 sg13g2_fill_1 FILLER_59_486 ();
 sg13g2_fill_1 FILLER_59_495 ();
 sg13g2_fill_2 FILLER_59_500 ();
 sg13g2_decap_8 FILLER_59_511 ();
 sg13g2_fill_2 FILLER_59_518 ();
 sg13g2_decap_8 FILLER_59_536 ();
 sg13g2_decap_8 FILLER_59_547 ();
 sg13g2_fill_1 FILLER_59_554 ();
 sg13g2_decap_8 FILLER_59_607 ();
 sg13g2_fill_1 FILLER_59_614 ();
 sg13g2_fill_1 FILLER_59_670 ();
 sg13g2_decap_4 FILLER_59_684 ();
 sg13g2_decap_8 FILLER_59_701 ();
 sg13g2_decap_4 FILLER_59_708 ();
 sg13g2_decap_4 FILLER_59_725 ();
 sg13g2_decap_8 FILLER_59_741 ();
 sg13g2_decap_4 FILLER_59_771 ();
 sg13g2_fill_2 FILLER_59_775 ();
 sg13g2_decap_8 FILLER_59_781 ();
 sg13g2_decap_8 FILLER_59_788 ();
 sg13g2_decap_8 FILLER_59_795 ();
 sg13g2_decap_8 FILLER_59_802 ();
 sg13g2_decap_8 FILLER_59_809 ();
 sg13g2_decap_8 FILLER_59_816 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_decap_8 FILLER_59_830 ();
 sg13g2_decap_8 FILLER_59_837 ();
 sg13g2_decap_8 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_851 ();
 sg13g2_decap_4 FILLER_59_858 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_decap_4 FILLER_60_24 ();
 sg13g2_fill_1 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_43 ();
 sg13g2_decap_8 FILLER_60_50 ();
 sg13g2_decap_4 FILLER_60_57 ();
 sg13g2_fill_1 FILLER_60_61 ();
 sg13g2_fill_2 FILLER_60_65 ();
 sg13g2_fill_1 FILLER_60_67 ();
 sg13g2_decap_8 FILLER_60_78 ();
 sg13g2_decap_8 FILLER_60_85 ();
 sg13g2_fill_2 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_109 ();
 sg13g2_fill_1 FILLER_60_111 ();
 sg13g2_fill_2 FILLER_60_122 ();
 sg13g2_decap_4 FILLER_60_137 ();
 sg13g2_fill_2 FILLER_60_141 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_fill_2 FILLER_60_169 ();
 sg13g2_fill_1 FILLER_60_171 ();
 sg13g2_fill_1 FILLER_60_176 ();
 sg13g2_decap_4 FILLER_60_201 ();
 sg13g2_fill_2 FILLER_60_205 ();
 sg13g2_decap_8 FILLER_60_215 ();
 sg13g2_decap_8 FILLER_60_222 ();
 sg13g2_decap_8 FILLER_60_229 ();
 sg13g2_fill_1 FILLER_60_236 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_254 ();
 sg13g2_fill_1 FILLER_60_256 ();
 sg13g2_decap_8 FILLER_60_278 ();
 sg13g2_decap_4 FILLER_60_285 ();
 sg13g2_fill_1 FILLER_60_289 ();
 sg13g2_fill_2 FILLER_60_306 ();
 sg13g2_fill_1 FILLER_60_308 ();
 sg13g2_fill_2 FILLER_60_321 ();
 sg13g2_fill_2 FILLER_60_327 ();
 sg13g2_fill_2 FILLER_60_376 ();
 sg13g2_decap_4 FILLER_60_393 ();
 sg13g2_fill_2 FILLER_60_397 ();
 sg13g2_decap_8 FILLER_60_431 ();
 sg13g2_decap_4 FILLER_60_438 ();
 sg13g2_fill_1 FILLER_60_442 ();
 sg13g2_fill_2 FILLER_60_460 ();
 sg13g2_fill_1 FILLER_60_462 ();
 sg13g2_fill_2 FILLER_60_478 ();
 sg13g2_decap_4 FILLER_60_486 ();
 sg13g2_fill_2 FILLER_60_490 ();
 sg13g2_fill_1 FILLER_60_501 ();
 sg13g2_fill_2 FILLER_60_511 ();
 sg13g2_fill_1 FILLER_60_513 ();
 sg13g2_fill_2 FILLER_60_545 ();
 sg13g2_decap_8 FILLER_60_555 ();
 sg13g2_decap_4 FILLER_60_562 ();
 sg13g2_decap_4 FILLER_60_570 ();
 sg13g2_decap_4 FILLER_60_602 ();
 sg13g2_fill_1 FILLER_60_606 ();
 sg13g2_fill_2 FILLER_60_620 ();
 sg13g2_fill_1 FILLER_60_622 ();
 sg13g2_fill_1 FILLER_60_628 ();
 sg13g2_fill_2 FILLER_60_632 ();
 sg13g2_fill_2 FILLER_60_653 ();
 sg13g2_fill_2 FILLER_60_709 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_fill_2 FILLER_60_731 ();
 sg13g2_fill_1 FILLER_60_733 ();
 sg13g2_decap_8 FILLER_60_738 ();
 sg13g2_decap_4 FILLER_60_745 ();
 sg13g2_fill_2 FILLER_60_752 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_836 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_fill_2 FILLER_61_45 ();
 sg13g2_fill_1 FILLER_61_47 ();
 sg13g2_fill_1 FILLER_61_61 ();
 sg13g2_fill_2 FILLER_61_87 ();
 sg13g2_fill_1 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_116 ();
 sg13g2_fill_1 FILLER_61_118 ();
 sg13g2_decap_4 FILLER_61_135 ();
 sg13g2_fill_1 FILLER_61_139 ();
 sg13g2_decap_8 FILLER_61_158 ();
 sg13g2_decap_8 FILLER_61_165 ();
 sg13g2_fill_2 FILLER_61_172 ();
 sg13g2_fill_2 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_181 ();
 sg13g2_decap_4 FILLER_61_199 ();
 sg13g2_decap_8 FILLER_61_207 ();
 sg13g2_decap_8 FILLER_61_214 ();
 sg13g2_fill_1 FILLER_61_228 ();
 sg13g2_fill_1 FILLER_61_239 ();
 sg13g2_decap_8 FILLER_61_257 ();
 sg13g2_decap_8 FILLER_61_269 ();
 sg13g2_decap_8 FILLER_61_276 ();
 sg13g2_decap_4 FILLER_61_283 ();
 sg13g2_fill_2 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_decap_4 FILLER_61_301 ();
 sg13g2_fill_2 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_321 ();
 sg13g2_fill_1 FILLER_61_328 ();
 sg13g2_decap_8 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_341 ();
 sg13g2_fill_1 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_decap_4 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_368 ();
 sg13g2_decap_4 FILLER_61_445 ();
 sg13g2_fill_1 FILLER_61_449 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_466 ();
 sg13g2_fill_2 FILLER_61_472 ();
 sg13g2_fill_1 FILLER_61_474 ();
 sg13g2_fill_1 FILLER_61_516 ();
 sg13g2_decap_4 FILLER_61_579 ();
 sg13g2_fill_1 FILLER_61_607 ();
 sg13g2_decap_8 FILLER_61_624 ();
 sg13g2_fill_2 FILLER_61_631 ();
 sg13g2_fill_1 FILLER_61_633 ();
 sg13g2_fill_1 FILLER_61_643 ();
 sg13g2_fill_1 FILLER_61_653 ();
 sg13g2_fill_1 FILLER_61_686 ();
 sg13g2_decap_4 FILLER_61_696 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_decap_8 FILLER_61_705 ();
 sg13g2_fill_2 FILLER_61_712 ();
 sg13g2_fill_1 FILLER_61_714 ();
 sg13g2_decap_4 FILLER_61_718 ();
 sg13g2_fill_1 FILLER_61_722 ();
 sg13g2_decap_4 FILLER_61_749 ();
 sg13g2_decap_8 FILLER_61_757 ();
 sg13g2_decap_8 FILLER_61_768 ();
 sg13g2_decap_8 FILLER_61_775 ();
 sg13g2_decap_8 FILLER_61_782 ();
 sg13g2_decap_8 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_796 ();
 sg13g2_decap_8 FILLER_61_803 ();
 sg13g2_decap_8 FILLER_61_810 ();
 sg13g2_decap_8 FILLER_61_817 ();
 sg13g2_decap_8 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_decap_8 FILLER_61_838 ();
 sg13g2_decap_8 FILLER_61_845 ();
 sg13g2_decap_8 FILLER_61_852 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_11 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_fill_2 FILLER_62_25 ();
 sg13g2_decap_4 FILLER_62_48 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_fill_1 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_69 ();
 sg13g2_decap_4 FILLER_62_75 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_4 FILLER_62_91 ();
 sg13g2_fill_2 FILLER_62_95 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_fill_1 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_128 ();
 sg13g2_decap_8 FILLER_62_135 ();
 sg13g2_decap_8 FILLER_62_165 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_decap_4 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_decap_8 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_251 ();
 sg13g2_fill_1 FILLER_62_253 ();
 sg13g2_decap_8 FILLER_62_258 ();
 sg13g2_decap_8 FILLER_62_265 ();
 sg13g2_decap_4 FILLER_62_272 ();
 sg13g2_fill_1 FILLER_62_276 ();
 sg13g2_fill_2 FILLER_62_284 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_fill_1 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_314 ();
 sg13g2_fill_2 FILLER_62_321 ();
 sg13g2_decap_8 FILLER_62_345 ();
 sg13g2_fill_1 FILLER_62_352 ();
 sg13g2_decap_4 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_62_376 ();
 sg13g2_fill_2 FILLER_62_387 ();
 sg13g2_fill_1 FILLER_62_393 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_414 ();
 sg13g2_fill_1 FILLER_62_416 ();
 sg13g2_fill_2 FILLER_62_431 ();
 sg13g2_decap_4 FILLER_62_445 ();
 sg13g2_fill_2 FILLER_62_474 ();
 sg13g2_fill_1 FILLER_62_476 ();
 sg13g2_decap_4 FILLER_62_485 ();
 sg13g2_decap_8 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_499 ();
 sg13g2_fill_1 FILLER_62_501 ();
 sg13g2_fill_1 FILLER_62_528 ();
 sg13g2_decap_8 FILLER_62_572 ();
 sg13g2_fill_2 FILLER_62_587 ();
 sg13g2_decap_8 FILLER_62_605 ();
 sg13g2_decap_4 FILLER_62_612 ();
 sg13g2_fill_2 FILLER_62_673 ();
 sg13g2_decap_4 FILLER_62_716 ();
 sg13g2_fill_1 FILLER_62_720 ();
 sg13g2_fill_1 FILLER_62_753 ();
 sg13g2_decap_8 FILLER_62_763 ();
 sg13g2_decap_8 FILLER_62_770 ();
 sg13g2_decap_8 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_798 ();
 sg13g2_decap_8 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_4 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_45 ();
 sg13g2_fill_2 FILLER_63_60 ();
 sg13g2_fill_2 FILLER_63_84 ();
 sg13g2_fill_1 FILLER_63_86 ();
 sg13g2_decap_4 FILLER_63_118 ();
 sg13g2_fill_2 FILLER_63_122 ();
 sg13g2_decap_8 FILLER_63_150 ();
 sg13g2_decap_8 FILLER_63_157 ();
 sg13g2_fill_1 FILLER_63_179 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_4 FILLER_63_206 ();
 sg13g2_fill_1 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_221 ();
 sg13g2_fill_1 FILLER_63_228 ();
 sg13g2_decap_8 FILLER_63_234 ();
 sg13g2_decap_4 FILLER_63_241 ();
 sg13g2_fill_2 FILLER_63_245 ();
 sg13g2_decap_4 FILLER_63_252 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_284 ();
 sg13g2_fill_2 FILLER_63_298 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_332 ();
 sg13g2_decap_8 FILLER_63_339 ();
 sg13g2_decap_4 FILLER_63_346 ();
 sg13g2_fill_2 FILLER_63_350 ();
 sg13g2_decap_4 FILLER_63_376 ();
 sg13g2_fill_2 FILLER_63_393 ();
 sg13g2_fill_1 FILLER_63_395 ();
 sg13g2_decap_4 FILLER_63_418 ();
 sg13g2_decap_8 FILLER_63_433 ();
 sg13g2_fill_1 FILLER_63_440 ();
 sg13g2_decap_8 FILLER_63_449 ();
 sg13g2_decap_8 FILLER_63_456 ();
 sg13g2_fill_1 FILLER_63_463 ();
 sg13g2_decap_8 FILLER_63_491 ();
 sg13g2_decap_4 FILLER_63_507 ();
 sg13g2_fill_2 FILLER_63_511 ();
 sg13g2_decap_8 FILLER_63_517 ();
 sg13g2_decap_8 FILLER_63_529 ();
 sg13g2_fill_1 FILLER_63_536 ();
 sg13g2_fill_2 FILLER_63_544 ();
 sg13g2_fill_1 FILLER_63_546 ();
 sg13g2_decap_8 FILLER_63_556 ();
 sg13g2_fill_2 FILLER_63_563 ();
 sg13g2_decap_8 FILLER_63_569 ();
 sg13g2_decap_8 FILLER_63_576 ();
 sg13g2_decap_8 FILLER_63_583 ();
 sg13g2_fill_1 FILLER_63_590 ();
 sg13g2_fill_2 FILLER_63_609 ();
 sg13g2_fill_1 FILLER_63_611 ();
 sg13g2_decap_8 FILLER_63_629 ();
 sg13g2_fill_2 FILLER_63_636 ();
 sg13g2_decap_4 FILLER_63_651 ();
 sg13g2_fill_1 FILLER_63_655 ();
 sg13g2_decap_4 FILLER_63_659 ();
 sg13g2_fill_2 FILLER_63_710 ();
 sg13g2_fill_1 FILLER_63_712 ();
 sg13g2_fill_1 FILLER_63_717 ();
 sg13g2_decap_8 FILLER_63_726 ();
 sg13g2_decap_8 FILLER_63_768 ();
 sg13g2_decap_8 FILLER_63_775 ();
 sg13g2_decap_8 FILLER_63_782 ();
 sg13g2_decap_8 FILLER_63_789 ();
 sg13g2_decap_8 FILLER_63_796 ();
 sg13g2_decap_8 FILLER_63_803 ();
 sg13g2_decap_8 FILLER_63_810 ();
 sg13g2_decap_8 FILLER_63_817 ();
 sg13g2_decap_8 FILLER_63_824 ();
 sg13g2_decap_8 FILLER_63_831 ();
 sg13g2_decap_8 FILLER_63_838 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_2 FILLER_64_26 ();
 sg13g2_fill_1 FILLER_64_28 ();
 sg13g2_decap_4 FILLER_64_57 ();
 sg13g2_fill_1 FILLER_64_61 ();
 sg13g2_decap_8 FILLER_64_78 ();
 sg13g2_fill_2 FILLER_64_85 ();
 sg13g2_fill_1 FILLER_64_87 ();
 sg13g2_decap_8 FILLER_64_103 ();
 sg13g2_decap_4 FILLER_64_110 ();
 sg13g2_fill_2 FILLER_64_114 ();
 sg13g2_decap_4 FILLER_64_155 ();
 sg13g2_decap_8 FILLER_64_170 ();
 sg13g2_decap_4 FILLER_64_177 ();
 sg13g2_fill_2 FILLER_64_209 ();
 sg13g2_fill_1 FILLER_64_211 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_fill_1 FILLER_64_273 ();
 sg13g2_decap_4 FILLER_64_279 ();
 sg13g2_fill_1 FILLER_64_283 ();
 sg13g2_decap_8 FILLER_64_289 ();
 sg13g2_fill_2 FILLER_64_296 ();
 sg13g2_fill_1 FILLER_64_298 ();
 sg13g2_decap_4 FILLER_64_303 ();
 sg13g2_fill_1 FILLER_64_307 ();
 sg13g2_decap_8 FILLER_64_318 ();
 sg13g2_decap_4 FILLER_64_325 ();
 sg13g2_fill_2 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_fill_2 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_359 ();
 sg13g2_fill_2 FILLER_64_365 ();
 sg13g2_fill_2 FILLER_64_382 ();
 sg13g2_fill_1 FILLER_64_384 ();
 sg13g2_fill_2 FILLER_64_390 ();
 sg13g2_fill_2 FILLER_64_404 ();
 sg13g2_fill_1 FILLER_64_414 ();
 sg13g2_fill_1 FILLER_64_423 ();
 sg13g2_decap_8 FILLER_64_437 ();
 sg13g2_fill_1 FILLER_64_444 ();
 sg13g2_decap_8 FILLER_64_467 ();
 sg13g2_decap_4 FILLER_64_474 ();
 sg13g2_fill_1 FILLER_64_478 ();
 sg13g2_fill_1 FILLER_64_483 ();
 sg13g2_fill_2 FILLER_64_517 ();
 sg13g2_fill_1 FILLER_64_519 ();
 sg13g2_fill_1 FILLER_64_525 ();
 sg13g2_fill_2 FILLER_64_552 ();
 sg13g2_fill_2 FILLER_64_580 ();
 sg13g2_decap_4 FILLER_64_608 ();
 sg13g2_fill_1 FILLER_64_612 ();
 sg13g2_decap_8 FILLER_64_618 ();
 sg13g2_fill_2 FILLER_64_625 ();
 sg13g2_fill_1 FILLER_64_661 ();
 sg13g2_decap_4 FILLER_64_679 ();
 sg13g2_fill_2 FILLER_64_687 ();
 sg13g2_decap_4 FILLER_64_711 ();
 sg13g2_fill_1 FILLER_64_715 ();
 sg13g2_decap_8 FILLER_64_765 ();
 sg13g2_decap_8 FILLER_64_772 ();
 sg13g2_decap_8 FILLER_64_779 ();
 sg13g2_decap_8 FILLER_64_786 ();
 sg13g2_decap_8 FILLER_64_793 ();
 sg13g2_decap_8 FILLER_64_800 ();
 sg13g2_decap_8 FILLER_64_807 ();
 sg13g2_decap_8 FILLER_64_814 ();
 sg13g2_decap_8 FILLER_64_821 ();
 sg13g2_decap_8 FILLER_64_828 ();
 sg13g2_decap_8 FILLER_64_835 ();
 sg13g2_decap_8 FILLER_64_842 ();
 sg13g2_decap_8 FILLER_64_849 ();
 sg13g2_decap_4 FILLER_64_856 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_41 ();
 sg13g2_fill_2 FILLER_65_48 ();
 sg13g2_fill_1 FILLER_65_55 ();
 sg13g2_decap_8 FILLER_65_65 ();
 sg13g2_fill_2 FILLER_65_76 ();
 sg13g2_decap_4 FILLER_65_86 ();
 sg13g2_fill_1 FILLER_65_90 ();
 sg13g2_decap_8 FILLER_65_107 ();
 sg13g2_fill_2 FILLER_65_114 ();
 sg13g2_fill_2 FILLER_65_124 ();
 sg13g2_decap_8 FILLER_65_129 ();
 sg13g2_decap_8 FILLER_65_136 ();
 sg13g2_decap_4 FILLER_65_143 ();
 sg13g2_decap_8 FILLER_65_152 ();
 sg13g2_decap_8 FILLER_65_159 ();
 sg13g2_decap_4 FILLER_65_178 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_4 FILLER_65_203 ();
 sg13g2_decap_4 FILLER_65_213 ();
 sg13g2_decap_4 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_decap_4 FILLER_65_234 ();
 sg13g2_fill_1 FILLER_65_238 ();
 sg13g2_fill_2 FILLER_65_242 ();
 sg13g2_fill_1 FILLER_65_244 ();
 sg13g2_decap_8 FILLER_65_250 ();
 sg13g2_decap_8 FILLER_65_257 ();
 sg13g2_fill_1 FILLER_65_264 ();
 sg13g2_fill_1 FILLER_65_281 ();
 sg13g2_decap_4 FILLER_65_300 ();
 sg13g2_fill_1 FILLER_65_304 ();
 sg13g2_fill_1 FILLER_65_325 ();
 sg13g2_decap_8 FILLER_65_334 ();
 sg13g2_fill_2 FILLER_65_341 ();
 sg13g2_fill_1 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_356 ();
 sg13g2_decap_4 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_367 ();
 sg13g2_decap_8 FILLER_65_395 ();
 sg13g2_fill_2 FILLER_65_402 ();
 sg13g2_decap_8 FILLER_65_430 ();
 sg13g2_decap_8 FILLER_65_437 ();
 sg13g2_decap_4 FILLER_65_444 ();
 sg13g2_fill_1 FILLER_65_448 ();
 sg13g2_fill_1 FILLER_65_457 ();
 sg13g2_fill_1 FILLER_65_463 ();
 sg13g2_decap_8 FILLER_65_472 ();
 sg13g2_decap_8 FILLER_65_479 ();
 sg13g2_decap_8 FILLER_65_486 ();
 sg13g2_fill_2 FILLER_65_493 ();
 sg13g2_fill_2 FILLER_65_499 ();
 sg13g2_fill_1 FILLER_65_501 ();
 sg13g2_fill_2 FILLER_65_522 ();
 sg13g2_decap_4 FILLER_65_540 ();
 sg13g2_fill_2 FILLER_65_571 ();
 sg13g2_fill_1 FILLER_65_573 ();
 sg13g2_fill_2 FILLER_65_587 ();
 sg13g2_decap_4 FILLER_65_610 ();
 sg13g2_fill_1 FILLER_65_614 ();
 sg13g2_decap_4 FILLER_65_623 ();
 sg13g2_fill_2 FILLER_65_635 ();
 sg13g2_fill_1 FILLER_65_637 ();
 sg13g2_decap_8 FILLER_65_642 ();
 sg13g2_decap_8 FILLER_65_649 ();
 sg13g2_decap_8 FILLER_65_656 ();
 sg13g2_decap_8 FILLER_65_663 ();
 sg13g2_decap_8 FILLER_65_670 ();
 sg13g2_fill_2 FILLER_65_677 ();
 sg13g2_fill_1 FILLER_65_693 ();
 sg13g2_decap_8 FILLER_65_768 ();
 sg13g2_decap_8 FILLER_65_775 ();
 sg13g2_decap_8 FILLER_65_782 ();
 sg13g2_decap_8 FILLER_65_789 ();
 sg13g2_decap_8 FILLER_65_796 ();
 sg13g2_decap_8 FILLER_65_803 ();
 sg13g2_decap_8 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_817 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_831 ();
 sg13g2_decap_8 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_845 ();
 sg13g2_decap_8 FILLER_65_852 ();
 sg13g2_fill_2 FILLER_65_859 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_fill_2 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_113 ();
 sg13g2_fill_1 FILLER_66_115 ();
 sg13g2_decap_8 FILLER_66_129 ();
 sg13g2_decap_8 FILLER_66_136 ();
 sg13g2_decap_8 FILLER_66_149 ();
 sg13g2_fill_1 FILLER_66_156 ();
 sg13g2_decap_4 FILLER_66_182 ();
 sg13g2_fill_2 FILLER_66_186 ();
 sg13g2_decap_4 FILLER_66_197 ();
 sg13g2_fill_2 FILLER_66_201 ();
 sg13g2_fill_1 FILLER_66_219 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_fill_1 FILLER_66_235 ();
 sg13g2_decap_8 FILLER_66_262 ();
 sg13g2_decap_8 FILLER_66_269 ();
 sg13g2_fill_2 FILLER_66_286 ();
 sg13g2_decap_4 FILLER_66_309 ();
 sg13g2_fill_2 FILLER_66_313 ();
 sg13g2_fill_2 FILLER_66_319 ();
 sg13g2_fill_1 FILLER_66_321 ();
 sg13g2_decap_8 FILLER_66_335 ();
 sg13g2_fill_1 FILLER_66_342 ();
 sg13g2_fill_1 FILLER_66_346 ();
 sg13g2_decap_8 FILLER_66_364 ();
 sg13g2_decap_4 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_decap_4 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_423 ();
 sg13g2_fill_1 FILLER_66_427 ();
 sg13g2_decap_8 FILLER_66_433 ();
 sg13g2_fill_2 FILLER_66_440 ();
 sg13g2_fill_1 FILLER_66_442 ();
 sg13g2_fill_2 FILLER_66_460 ();
 sg13g2_fill_1 FILLER_66_462 ();
 sg13g2_fill_1 FILLER_66_471 ();
 sg13g2_fill_2 FILLER_66_491 ();
 sg13g2_fill_1 FILLER_66_493 ();
 sg13g2_decap_8 FILLER_66_511 ();
 sg13g2_decap_4 FILLER_66_518 ();
 sg13g2_decap_8 FILLER_66_531 ();
 sg13g2_decap_8 FILLER_66_538 ();
 sg13g2_fill_1 FILLER_66_545 ();
 sg13g2_fill_1 FILLER_66_561 ();
 sg13g2_decap_4 FILLER_66_588 ();
 sg13g2_fill_2 FILLER_66_625 ();
 sg13g2_fill_1 FILLER_66_627 ();
 sg13g2_fill_2 FILLER_66_654 ();
 sg13g2_decap_8 FILLER_66_673 ();
 sg13g2_fill_2 FILLER_66_680 ();
 sg13g2_fill_2 FILLER_66_686 ();
 sg13g2_fill_1 FILLER_66_688 ();
 sg13g2_fill_2 FILLER_66_711 ();
 sg13g2_fill_1 FILLER_66_713 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_4 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_47 ();
 sg13g2_fill_2 FILLER_67_54 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_60 ();
 sg13g2_fill_1 FILLER_67_62 ();
 sg13g2_decap_8 FILLER_67_68 ();
 sg13g2_fill_2 FILLER_67_85 ();
 sg13g2_fill_1 FILLER_67_87 ();
 sg13g2_fill_1 FILLER_67_92 ();
 sg13g2_fill_2 FILLER_67_97 ();
 sg13g2_fill_1 FILLER_67_99 ();
 sg13g2_decap_4 FILLER_67_121 ();
 sg13g2_decap_4 FILLER_67_143 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_fill_1 FILLER_67_153 ();
 sg13g2_decap_4 FILLER_67_158 ();
 sg13g2_fill_2 FILLER_67_162 ();
 sg13g2_decap_8 FILLER_67_176 ();
 sg13g2_decap_4 FILLER_67_183 ();
 sg13g2_fill_2 FILLER_67_202 ();
 sg13g2_fill_1 FILLER_67_204 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_fill_2 FILLER_67_245 ();
 sg13g2_fill_1 FILLER_67_247 ();
 sg13g2_decap_8 FILLER_67_253 ();
 sg13g2_fill_2 FILLER_67_260 ();
 sg13g2_decap_8 FILLER_67_291 ();
 sg13g2_decap_8 FILLER_67_298 ();
 sg13g2_decap_8 FILLER_67_305 ();
 sg13g2_fill_2 FILLER_67_312 ();
 sg13g2_decap_8 FILLER_67_319 ();
 sg13g2_fill_2 FILLER_67_326 ();
 sg13g2_fill_1 FILLER_67_328 ();
 sg13g2_fill_2 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_344 ();
 sg13g2_decap_8 FILLER_67_353 ();
 sg13g2_fill_2 FILLER_67_360 ();
 sg13g2_fill_1 FILLER_67_362 ();
 sg13g2_fill_1 FILLER_67_386 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_fill_2 FILLER_67_413 ();
 sg13g2_fill_1 FILLER_67_415 ();
 sg13g2_decap_8 FILLER_67_450 ();
 sg13g2_decap_8 FILLER_67_465 ();
 sg13g2_decap_8 FILLER_67_472 ();
 sg13g2_decap_8 FILLER_67_479 ();
 sg13g2_decap_4 FILLER_67_486 ();
 sg13g2_fill_2 FILLER_67_490 ();
 sg13g2_decap_4 FILLER_67_553 ();
 sg13g2_fill_2 FILLER_67_557 ();
 sg13g2_decap_8 FILLER_67_573 ();
 sg13g2_fill_2 FILLER_67_580 ();
 sg13g2_fill_2 FILLER_67_586 ();
 sg13g2_decap_8 FILLER_67_593 ();
 sg13g2_fill_2 FILLER_67_600 ();
 sg13g2_fill_1 FILLER_67_602 ();
 sg13g2_fill_2 FILLER_67_667 ();
 sg13g2_decap_4 FILLER_67_713 ();
 sg13g2_fill_1 FILLER_67_721 ();
 sg13g2_decap_8 FILLER_67_735 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_749 ();
 sg13g2_decap_8 FILLER_67_756 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_8 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_decap_4 FILLER_68_41 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_59 ();
 sg13g2_fill_1 FILLER_68_61 ();
 sg13g2_fill_2 FILLER_68_76 ();
 sg13g2_fill_1 FILLER_68_78 ();
 sg13g2_fill_1 FILLER_68_90 ();
 sg13g2_decap_4 FILLER_68_115 ();
 sg13g2_fill_2 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_139 ();
 sg13g2_decap_8 FILLER_68_146 ();
 sg13g2_decap_4 FILLER_68_153 ();
 sg13g2_fill_1 FILLER_68_169 ();
 sg13g2_fill_1 FILLER_68_175 ();
 sg13g2_decap_4 FILLER_68_191 ();
 sg13g2_fill_2 FILLER_68_202 ();
 sg13g2_fill_2 FILLER_68_209 ();
 sg13g2_fill_1 FILLER_68_216 ();
 sg13g2_decap_8 FILLER_68_222 ();
 sg13g2_decap_4 FILLER_68_229 ();
 sg13g2_fill_1 FILLER_68_241 ();
 sg13g2_decap_8 FILLER_68_247 ();
 sg13g2_decap_4 FILLER_68_254 ();
 sg13g2_fill_2 FILLER_68_258 ();
 sg13g2_fill_2 FILLER_68_272 ();
 sg13g2_fill_1 FILLER_68_274 ();
 sg13g2_decap_8 FILLER_68_293 ();
 sg13g2_fill_2 FILLER_68_300 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_decap_4 FILLER_68_336 ();
 sg13g2_decap_4 FILLER_68_353 ();
 sg13g2_fill_1 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_365 ();
 sg13g2_fill_1 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_411 ();
 sg13g2_decap_8 FILLER_68_418 ();
 sg13g2_decap_8 FILLER_68_425 ();
 sg13g2_decap_8 FILLER_68_432 ();
 sg13g2_decap_8 FILLER_68_439 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_fill_2 FILLER_68_485 ();
 sg13g2_decap_8 FILLER_68_491 ();
 sg13g2_decap_4 FILLER_68_498 ();
 sg13g2_fill_2 FILLER_68_502 ();
 sg13g2_decap_8 FILLER_68_512 ();
 sg13g2_decap_8 FILLER_68_519 ();
 sg13g2_decap_8 FILLER_68_526 ();
 sg13g2_fill_2 FILLER_68_546 ();
 sg13g2_decap_8 FILLER_68_566 ();
 sg13g2_fill_2 FILLER_68_573 ();
 sg13g2_fill_1 FILLER_68_584 ();
 sg13g2_decap_8 FILLER_68_590 ();
 sg13g2_decap_8 FILLER_68_597 ();
 sg13g2_decap_4 FILLER_68_604 ();
 sg13g2_fill_1 FILLER_68_608 ();
 sg13g2_decap_8 FILLER_68_623 ();
 sg13g2_fill_2 FILLER_68_630 ();
 sg13g2_decap_4 FILLER_68_652 ();
 sg13g2_fill_2 FILLER_68_656 ();
 sg13g2_decap_8 FILLER_68_663 ();
 sg13g2_fill_2 FILLER_68_670 ();
 sg13g2_fill_1 FILLER_68_685 ();
 sg13g2_fill_2 FILLER_68_704 ();
 sg13g2_fill_1 FILLER_68_706 ();
 sg13g2_decap_8 FILLER_68_733 ();
 sg13g2_decap_8 FILLER_68_740 ();
 sg13g2_decap_8 FILLER_68_747 ();
 sg13g2_decap_8 FILLER_68_754 ();
 sg13g2_decap_8 FILLER_68_761 ();
 sg13g2_decap_8 FILLER_68_768 ();
 sg13g2_decap_8 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_782 ();
 sg13g2_decap_8 FILLER_68_789 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_810 ();
 sg13g2_decap_8 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_824 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_decap_8 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_852 ();
 sg13g2_fill_2 FILLER_68_859 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_16 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_68 ();
 sg13g2_fill_1 FILLER_69_75 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_117 ();
 sg13g2_fill_2 FILLER_69_124 ();
 sg13g2_fill_1 FILLER_69_126 ();
 sg13g2_decap_4 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_137 ();
 sg13g2_decap_4 FILLER_69_147 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_fill_2 FILLER_69_157 ();
 sg13g2_decap_8 FILLER_69_164 ();
 sg13g2_decap_8 FILLER_69_171 ();
 sg13g2_decap_8 FILLER_69_178 ();
 sg13g2_decap_8 FILLER_69_194 ();
 sg13g2_decap_8 FILLER_69_201 ();
 sg13g2_decap_4 FILLER_69_208 ();
 sg13g2_fill_2 FILLER_69_225 ();
 sg13g2_fill_1 FILLER_69_227 ();
 sg13g2_decap_8 FILLER_69_266 ();
 sg13g2_fill_2 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_299 ();
 sg13g2_decap_4 FILLER_69_326 ();
 sg13g2_fill_2 FILLER_69_330 ();
 sg13g2_fill_2 FILLER_69_348 ();
 sg13g2_fill_1 FILLER_69_362 ();
 sg13g2_fill_2 FILLER_69_376 ();
 sg13g2_decap_4 FILLER_69_383 ();
 sg13g2_fill_1 FILLER_69_387 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_fill_2 FILLER_69_402 ();
 sg13g2_fill_1 FILLER_69_404 ();
 sg13g2_decap_8 FILLER_69_426 ();
 sg13g2_decap_4 FILLER_69_433 ();
 sg13g2_fill_2 FILLER_69_437 ();
 sg13g2_decap_8 FILLER_69_452 ();
 sg13g2_decap_8 FILLER_69_464 ();
 sg13g2_decap_4 FILLER_69_471 ();
 sg13g2_fill_1 FILLER_69_475 ();
 sg13g2_fill_2 FILLER_69_502 ();
 sg13g2_decap_8 FILLER_69_530 ();
 sg13g2_fill_2 FILLER_69_550 ();
 sg13g2_decap_8 FILLER_69_557 ();
 sg13g2_fill_1 FILLER_69_564 ();
 sg13g2_fill_2 FILLER_69_596 ();
 sg13g2_fill_1 FILLER_69_598 ();
 sg13g2_fill_2 FILLER_69_612 ();
 sg13g2_fill_1 FILLER_69_614 ();
 sg13g2_decap_8 FILLER_69_620 ();
 sg13g2_decap_8 FILLER_69_627 ();
 sg13g2_fill_2 FILLER_69_634 ();
 sg13g2_fill_1 FILLER_69_636 ();
 sg13g2_decap_8 FILLER_69_650 ();
 sg13g2_fill_2 FILLER_69_686 ();
 sg13g2_decap_8 FILLER_69_732 ();
 sg13g2_decap_8 FILLER_69_739 ();
 sg13g2_decap_8 FILLER_69_746 ();
 sg13g2_decap_8 FILLER_69_753 ();
 sg13g2_decap_8 FILLER_69_760 ();
 sg13g2_decap_8 FILLER_69_767 ();
 sg13g2_decap_8 FILLER_69_774 ();
 sg13g2_decap_8 FILLER_69_781 ();
 sg13g2_decap_8 FILLER_69_788 ();
 sg13g2_decap_8 FILLER_69_795 ();
 sg13g2_decap_8 FILLER_69_802 ();
 sg13g2_decap_8 FILLER_69_809 ();
 sg13g2_decap_8 FILLER_69_816 ();
 sg13g2_decap_8 FILLER_69_823 ();
 sg13g2_decap_8 FILLER_69_830 ();
 sg13g2_decap_8 FILLER_69_837 ();
 sg13g2_decap_8 FILLER_69_844 ();
 sg13g2_decap_8 FILLER_69_851 ();
 sg13g2_decap_4 FILLER_69_858 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_fill_1 FILLER_70_88 ();
 sg13g2_decap_8 FILLER_70_94 ();
 sg13g2_decap_4 FILLER_70_101 ();
 sg13g2_fill_2 FILLER_70_105 ();
 sg13g2_fill_2 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_146 ();
 sg13g2_fill_1 FILLER_70_148 ();
 sg13g2_fill_1 FILLER_70_162 ();
 sg13g2_fill_2 FILLER_70_177 ();
 sg13g2_decap_4 FILLER_70_188 ();
 sg13g2_fill_2 FILLER_70_204 ();
 sg13g2_decap_8 FILLER_70_215 ();
 sg13g2_fill_2 FILLER_70_227 ();
 sg13g2_decap_8 FILLER_70_247 ();
 sg13g2_decap_4 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_258 ();
 sg13g2_decap_8 FILLER_70_267 ();
 sg13g2_fill_1 FILLER_70_274 ();
 sg13g2_decap_8 FILLER_70_283 ();
 sg13g2_decap_8 FILLER_70_290 ();
 sg13g2_fill_2 FILLER_70_297 ();
 sg13g2_fill_1 FILLER_70_299 ();
 sg13g2_fill_1 FILLER_70_316 ();
 sg13g2_decap_8 FILLER_70_325 ();
 sg13g2_decap_8 FILLER_70_332 ();
 sg13g2_fill_2 FILLER_70_339 ();
 sg13g2_fill_1 FILLER_70_341 ();
 sg13g2_decap_8 FILLER_70_346 ();
 sg13g2_decap_4 FILLER_70_353 ();
 sg13g2_fill_2 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_373 ();
 sg13g2_decap_4 FILLER_70_380 ();
 sg13g2_fill_1 FILLER_70_384 ();
 sg13g2_fill_2 FILLER_70_389 ();
 sg13g2_fill_1 FILLER_70_391 ();
 sg13g2_decap_4 FILLER_70_409 ();
 sg13g2_decap_4 FILLER_70_423 ();
 sg13g2_fill_1 FILLER_70_427 ();
 sg13g2_decap_4 FILLER_70_449 ();
 sg13g2_fill_1 FILLER_70_453 ();
 sg13g2_decap_4 FILLER_70_459 ();
 sg13g2_fill_1 FILLER_70_470 ();
 sg13g2_decap_8 FILLER_70_477 ();
 sg13g2_decap_8 FILLER_70_484 ();
 sg13g2_decap_8 FILLER_70_491 ();
 sg13g2_fill_1 FILLER_70_520 ();
 sg13g2_decap_8 FILLER_70_567 ();
 sg13g2_decap_4 FILLER_70_574 ();
 sg13g2_fill_1 FILLER_70_578 ();
 sg13g2_decap_8 FILLER_70_583 ();
 sg13g2_decap_8 FILLER_70_626 ();
 sg13g2_decap_4 FILLER_70_661 ();
 sg13g2_fill_2 FILLER_70_665 ();
 sg13g2_decap_8 FILLER_70_675 ();
 sg13g2_fill_2 FILLER_70_682 ();
 sg13g2_fill_1 FILLER_70_684 ();
 sg13g2_fill_2 FILLER_70_702 ();
 sg13g2_fill_1 FILLER_70_704 ();
 sg13g2_decap_8 FILLER_70_735 ();
 sg13g2_decap_8 FILLER_70_742 ();
 sg13g2_decap_8 FILLER_70_749 ();
 sg13g2_decap_8 FILLER_70_756 ();
 sg13g2_decap_8 FILLER_70_763 ();
 sg13g2_decap_8 FILLER_70_770 ();
 sg13g2_decap_8 FILLER_70_777 ();
 sg13g2_decap_8 FILLER_70_784 ();
 sg13g2_decap_8 FILLER_70_791 ();
 sg13g2_decap_8 FILLER_70_798 ();
 sg13g2_decap_8 FILLER_70_805 ();
 sg13g2_decap_8 FILLER_70_812 ();
 sg13g2_decap_8 FILLER_70_819 ();
 sg13g2_decap_8 FILLER_70_826 ();
 sg13g2_decap_8 FILLER_70_833 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_fill_2 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_79 ();
 sg13g2_decap_4 FILLER_71_106 ();
 sg13g2_decap_4 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_decap_4 FILLER_71_128 ();
 sg13g2_decap_4 FILLER_71_137 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_fill_1 FILLER_71_175 ();
 sg13g2_fill_2 FILLER_71_191 ();
 sg13g2_fill_1 FILLER_71_193 ();
 sg13g2_fill_2 FILLER_71_205 ();
 sg13g2_fill_1 FILLER_71_207 ();
 sg13g2_decap_4 FILLER_71_233 ();
 sg13g2_fill_2 FILLER_71_240 ();
 sg13g2_fill_1 FILLER_71_242 ();
 sg13g2_decap_8 FILLER_71_248 ();
 sg13g2_decap_8 FILLER_71_255 ();
 sg13g2_fill_2 FILLER_71_262 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_295 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_fill_2 FILLER_71_315 ();
 sg13g2_fill_1 FILLER_71_317 ();
 sg13g2_decap_8 FILLER_71_331 ();
 sg13g2_decap_4 FILLER_71_352 ();
 sg13g2_decap_4 FILLER_71_377 ();
 sg13g2_fill_1 FILLER_71_395 ();
 sg13g2_decap_4 FILLER_71_404 ();
 sg13g2_decap_4 FILLER_71_413 ();
 sg13g2_fill_2 FILLER_71_437 ();
 sg13g2_decap_8 FILLER_71_444 ();
 sg13g2_decap_4 FILLER_71_451 ();
 sg13g2_decap_8 FILLER_71_459 ();
 sg13g2_fill_2 FILLER_71_466 ();
 sg13g2_fill_1 FILLER_71_478 ();
 sg13g2_decap_8 FILLER_71_487 ();
 sg13g2_decap_8 FILLER_71_494 ();
 sg13g2_decap_4 FILLER_71_539 ();
 sg13g2_fill_2 FILLER_71_543 ();
 sg13g2_fill_2 FILLER_71_549 ();
 sg13g2_fill_1 FILLER_71_551 ();
 sg13g2_decap_4 FILLER_71_565 ();
 sg13g2_fill_2 FILLER_71_586 ();
 sg13g2_fill_1 FILLER_71_592 ();
 sg13g2_decap_8 FILLER_71_602 ();
 sg13g2_fill_2 FILLER_71_613 ();
 sg13g2_fill_1 FILLER_71_615 ();
 sg13g2_decap_8 FILLER_71_621 ();
 sg13g2_decap_4 FILLER_71_628 ();
 sg13g2_fill_2 FILLER_71_632 ();
 sg13g2_fill_2 FILLER_71_644 ();
 sg13g2_fill_1 FILLER_71_646 ();
 sg13g2_decap_4 FILLER_71_682 ();
 sg13g2_fill_1 FILLER_71_686 ();
 sg13g2_decap_8 FILLER_71_731 ();
 sg13g2_decap_8 FILLER_71_738 ();
 sg13g2_decap_8 FILLER_71_745 ();
 sg13g2_decap_8 FILLER_71_752 ();
 sg13g2_decap_8 FILLER_71_759 ();
 sg13g2_decap_8 FILLER_71_766 ();
 sg13g2_decap_8 FILLER_71_773 ();
 sg13g2_decap_8 FILLER_71_780 ();
 sg13g2_decap_8 FILLER_71_787 ();
 sg13g2_decap_8 FILLER_71_794 ();
 sg13g2_decap_8 FILLER_71_801 ();
 sg13g2_decap_8 FILLER_71_808 ();
 sg13g2_decap_8 FILLER_71_815 ();
 sg13g2_decap_8 FILLER_71_822 ();
 sg13g2_decap_8 FILLER_71_829 ();
 sg13g2_decap_8 FILLER_71_836 ();
 sg13g2_decap_8 FILLER_71_843 ();
 sg13g2_decap_8 FILLER_71_850 ();
 sg13g2_decap_4 FILLER_71_857 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_77 ();
 sg13g2_fill_1 FILLER_72_79 ();
 sg13g2_fill_1 FILLER_72_85 ();
 sg13g2_fill_1 FILLER_72_96 ();
 sg13g2_fill_2 FILLER_72_102 ();
 sg13g2_fill_2 FILLER_72_113 ();
 sg13g2_fill_1 FILLER_72_115 ();
 sg13g2_decap_8 FILLER_72_141 ();
 sg13g2_decap_4 FILLER_72_148 ();
 sg13g2_fill_1 FILLER_72_152 ();
 sg13g2_decap_8 FILLER_72_159 ();
 sg13g2_decap_8 FILLER_72_166 ();
 sg13g2_fill_2 FILLER_72_173 ();
 sg13g2_decap_8 FILLER_72_199 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_4 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_fill_2 FILLER_72_238 ();
 sg13g2_fill_1 FILLER_72_240 ();
 sg13g2_decap_4 FILLER_72_259 ();
 sg13g2_fill_1 FILLER_72_263 ();
 sg13g2_fill_2 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_302 ();
 sg13g2_decap_8 FILLER_72_309 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_decap_4 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_358 ();
 sg13g2_fill_1 FILLER_72_365 ();
 sg13g2_decap_8 FILLER_72_376 ();
 sg13g2_decap_4 FILLER_72_383 ();
 sg13g2_decap_4 FILLER_72_392 ();
 sg13g2_fill_2 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_72_412 ();
 sg13g2_decap_4 FILLER_72_419 ();
 sg13g2_fill_1 FILLER_72_423 ();
 sg13g2_decap_4 FILLER_72_433 ();
 sg13g2_decap_4 FILLER_72_451 ();
 sg13g2_fill_1 FILLER_72_455 ();
 sg13g2_fill_1 FILLER_72_476 ();
 sg13g2_decap_4 FILLER_72_482 ();
 sg13g2_fill_1 FILLER_72_486 ();
 sg13g2_fill_2 FILLER_72_517 ();
 sg13g2_fill_1 FILLER_72_519 ();
 sg13g2_decap_4 FILLER_72_573 ();
 sg13g2_fill_2 FILLER_72_623 ();
 sg13g2_fill_2 FILLER_72_646 ();
 sg13g2_decap_8 FILLER_72_671 ();
 sg13g2_decap_8 FILLER_72_678 ();
 sg13g2_fill_2 FILLER_72_685 ();
 sg13g2_decap_8 FILLER_72_722 ();
 sg13g2_decap_8 FILLER_72_729 ();
 sg13g2_decap_8 FILLER_72_736 ();
 sg13g2_decap_8 FILLER_72_743 ();
 sg13g2_decap_8 FILLER_72_750 ();
 sg13g2_decap_8 FILLER_72_757 ();
 sg13g2_decap_8 FILLER_72_764 ();
 sg13g2_decap_8 FILLER_72_771 ();
 sg13g2_decap_8 FILLER_72_778 ();
 sg13g2_decap_8 FILLER_72_785 ();
 sg13g2_decap_8 FILLER_72_792 ();
 sg13g2_decap_8 FILLER_72_799 ();
 sg13g2_decap_8 FILLER_72_806 ();
 sg13g2_decap_8 FILLER_72_813 ();
 sg13g2_decap_8 FILLER_72_820 ();
 sg13g2_decap_8 FILLER_72_827 ();
 sg13g2_decap_8 FILLER_72_834 ();
 sg13g2_decap_8 FILLER_72_841 ();
 sg13g2_decap_8 FILLER_72_848 ();
 sg13g2_decap_8 FILLER_72_855 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_fill_2 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_101 ();
 sg13g2_decap_4 FILLER_73_108 ();
 sg13g2_fill_1 FILLER_73_116 ();
 sg13g2_decap_8 FILLER_73_121 ();
 sg13g2_decap_8 FILLER_73_128 ();
 sg13g2_decap_8 FILLER_73_135 ();
 sg13g2_decap_4 FILLER_73_142 ();
 sg13g2_fill_1 FILLER_73_146 ();
 sg13g2_decap_4 FILLER_73_165 ();
 sg13g2_decap_8 FILLER_73_173 ();
 sg13g2_decap_4 FILLER_73_180 ();
 sg13g2_fill_2 FILLER_73_184 ();
 sg13g2_decap_4 FILLER_73_207 ();
 sg13g2_fill_2 FILLER_73_211 ();
 sg13g2_decap_4 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_decap_8 FILLER_73_256 ();
 sg13g2_decap_4 FILLER_73_263 ();
 sg13g2_fill_1 FILLER_73_267 ();
 sg13g2_decap_8 FILLER_73_274 ();
 sg13g2_fill_2 FILLER_73_281 ();
 sg13g2_fill_1 FILLER_73_283 ();
 sg13g2_fill_2 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_302 ();
 sg13g2_fill_2 FILLER_73_309 ();
 sg13g2_fill_1 FILLER_73_311 ();
 sg13g2_decap_8 FILLER_73_321 ();
 sg13g2_decap_8 FILLER_73_333 ();
 sg13g2_fill_2 FILLER_73_340 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_4 FILLER_73_357 ();
 sg13g2_fill_2 FILLER_73_361 ();
 sg13g2_fill_1 FILLER_73_373 ();
 sg13g2_fill_2 FILLER_73_392 ();
 sg13g2_decap_4 FILLER_73_409 ();
 sg13g2_fill_1 FILLER_73_413 ();
 sg13g2_fill_2 FILLER_73_441 ();
 sg13g2_fill_2 FILLER_73_453 ();
 sg13g2_fill_1 FILLER_73_455 ();
 sg13g2_fill_1 FILLER_73_468 ();
 sg13g2_fill_2 FILLER_73_478 ();
 sg13g2_fill_1 FILLER_73_480 ();
 sg13g2_decap_8 FILLER_73_486 ();
 sg13g2_decap_4 FILLER_73_493 ();
 sg13g2_fill_1 FILLER_73_497 ();
 sg13g2_decap_8 FILLER_73_502 ();
 sg13g2_decap_4 FILLER_73_509 ();
 sg13g2_decap_4 FILLER_73_518 ();
 sg13g2_fill_2 FILLER_73_522 ();
 sg13g2_fill_2 FILLER_73_536 ();
 sg13g2_fill_1 FILLER_73_538 ();
 sg13g2_decap_8 FILLER_73_550 ();
 sg13g2_fill_1 FILLER_73_557 ();
 sg13g2_fill_2 FILLER_73_576 ();
 sg13g2_fill_1 FILLER_73_578 ();
 sg13g2_decap_4 FILLER_73_591 ();
 sg13g2_fill_2 FILLER_73_595 ();
 sg13g2_decap_8 FILLER_73_602 ();
 sg13g2_decap_8 FILLER_73_609 ();
 sg13g2_decap_8 FILLER_73_616 ();
 sg13g2_fill_2 FILLER_73_627 ();
 sg13g2_fill_1 FILLER_73_629 ();
 sg13g2_decap_4 FILLER_73_637 ();
 sg13g2_fill_1 FILLER_73_641 ();
 sg13g2_decap_8 FILLER_73_674 ();
 sg13g2_decap_8 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_688 ();
 sg13g2_fill_2 FILLER_73_695 ();
 sg13g2_fill_1 FILLER_73_697 ();
 sg13g2_decap_8 FILLER_73_702 ();
 sg13g2_decap_8 FILLER_73_709 ();
 sg13g2_decap_8 FILLER_73_716 ();
 sg13g2_decap_8 FILLER_73_723 ();
 sg13g2_decap_8 FILLER_73_730 ();
 sg13g2_decap_8 FILLER_73_737 ();
 sg13g2_decap_8 FILLER_73_744 ();
 sg13g2_decap_8 FILLER_73_751 ();
 sg13g2_decap_8 FILLER_73_758 ();
 sg13g2_decap_8 FILLER_73_765 ();
 sg13g2_decap_8 FILLER_73_772 ();
 sg13g2_decap_8 FILLER_73_779 ();
 sg13g2_decap_8 FILLER_73_786 ();
 sg13g2_decap_8 FILLER_73_793 ();
 sg13g2_decap_8 FILLER_73_800 ();
 sg13g2_decap_8 FILLER_73_807 ();
 sg13g2_decap_8 FILLER_73_814 ();
 sg13g2_decap_8 FILLER_73_821 ();
 sg13g2_decap_8 FILLER_73_828 ();
 sg13g2_decap_8 FILLER_73_835 ();
 sg13g2_decap_8 FILLER_73_842 ();
 sg13g2_decap_8 FILLER_73_849 ();
 sg13g2_decap_4 FILLER_73_856 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_4 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_85 ();
 sg13g2_decap_4 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_105 ();
 sg13g2_decap_4 FILLER_74_110 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_148 ();
 sg13g2_fill_2 FILLER_74_165 ();
 sg13g2_decap_8 FILLER_74_179 ();
 sg13g2_decap_4 FILLER_74_186 ();
 sg13g2_fill_1 FILLER_74_190 ();
 sg13g2_fill_1 FILLER_74_195 ();
 sg13g2_decap_8 FILLER_74_209 ();
 sg13g2_decap_4 FILLER_74_216 ();
 sg13g2_fill_2 FILLER_74_220 ();
 sg13g2_decap_8 FILLER_74_232 ();
 sg13g2_fill_2 FILLER_74_239 ();
 sg13g2_fill_1 FILLER_74_241 ();
 sg13g2_decap_8 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_268 ();
 sg13g2_fill_2 FILLER_74_282 ();
 sg13g2_fill_1 FILLER_74_284 ();
 sg13g2_fill_1 FILLER_74_306 ();
 sg13g2_decap_4 FILLER_74_331 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_fill_2 FILLER_74_364 ();
 sg13g2_fill_1 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_fill_2 FILLER_74_399 ();
 sg13g2_fill_1 FILLER_74_401 ();
 sg13g2_decap_8 FILLER_74_411 ();
 sg13g2_decap_4 FILLER_74_418 ();
 sg13g2_decap_8 FILLER_74_431 ();
 sg13g2_decap_8 FILLER_74_438 ();
 sg13g2_decap_8 FILLER_74_445 ();
 sg13g2_decap_8 FILLER_74_494 ();
 sg13g2_decap_8 FILLER_74_501 ();
 sg13g2_decap_4 FILLER_74_524 ();
 sg13g2_fill_2 FILLER_74_541 ();
 sg13g2_fill_2 FILLER_74_552 ();
 sg13g2_fill_1 FILLER_74_554 ();
 sg13g2_fill_2 FILLER_74_568 ();
 sg13g2_fill_1 FILLER_74_570 ();
 sg13g2_fill_1 FILLER_74_619 ();
 sg13g2_decap_8 FILLER_74_649 ();
 sg13g2_decap_8 FILLER_74_656 ();
 sg13g2_decap_8 FILLER_74_663 ();
 sg13g2_decap_8 FILLER_74_670 ();
 sg13g2_decap_8 FILLER_74_677 ();
 sg13g2_decap_8 FILLER_74_684 ();
 sg13g2_decap_8 FILLER_74_691 ();
 sg13g2_decap_8 FILLER_74_698 ();
 sg13g2_decap_8 FILLER_74_705 ();
 sg13g2_decap_8 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_719 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_740 ();
 sg13g2_decap_8 FILLER_74_747 ();
 sg13g2_decap_8 FILLER_74_754 ();
 sg13g2_decap_8 FILLER_74_761 ();
 sg13g2_decap_8 FILLER_74_768 ();
 sg13g2_decap_8 FILLER_74_775 ();
 sg13g2_decap_8 FILLER_74_782 ();
 sg13g2_decap_8 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_796 ();
 sg13g2_decap_8 FILLER_74_803 ();
 sg13g2_decap_8 FILLER_74_810 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_8 FILLER_74_824 ();
 sg13g2_decap_8 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_4 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_117 ();
 sg13g2_decap_8 FILLER_75_124 ();
 sg13g2_fill_1 FILLER_75_131 ();
 sg13g2_fill_1 FILLER_75_153 ();
 sg13g2_decap_8 FILLER_75_171 ();
 sg13g2_decap_4 FILLER_75_178 ();
 sg13g2_fill_1 FILLER_75_182 ();
 sg13g2_fill_2 FILLER_75_191 ();
 sg13g2_fill_1 FILLER_75_193 ();
 sg13g2_fill_2 FILLER_75_211 ();
 sg13g2_fill_1 FILLER_75_213 ();
 sg13g2_decap_8 FILLER_75_240 ();
 sg13g2_decap_8 FILLER_75_247 ();
 sg13g2_decap_8 FILLER_75_254 ();
 sg13g2_decap_8 FILLER_75_261 ();
 sg13g2_fill_1 FILLER_75_268 ();
 sg13g2_fill_1 FILLER_75_275 ();
 sg13g2_fill_2 FILLER_75_285 ();
 sg13g2_fill_1 FILLER_75_287 ();
 sg13g2_fill_2 FILLER_75_300 ();
 sg13g2_fill_1 FILLER_75_302 ();
 sg13g2_decap_8 FILLER_75_309 ();
 sg13g2_fill_2 FILLER_75_316 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_fill_2 FILLER_75_335 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_decap_8 FILLER_75_354 ();
 sg13g2_fill_2 FILLER_75_361 ();
 sg13g2_decap_8 FILLER_75_369 ();
 sg13g2_decap_8 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_396 ();
 sg13g2_fill_2 FILLER_75_403 ();
 sg13g2_fill_1 FILLER_75_405 ();
 sg13g2_fill_1 FILLER_75_413 ();
 sg13g2_fill_2 FILLER_75_421 ();
 sg13g2_fill_1 FILLER_75_423 ();
 sg13g2_fill_2 FILLER_75_429 ();
 sg13g2_decap_4 FILLER_75_436 ();
 sg13g2_decap_8 FILLER_75_453 ();
 sg13g2_decap_8 FILLER_75_460 ();
 sg13g2_decap_4 FILLER_75_467 ();
 sg13g2_fill_2 FILLER_75_477 ();
 sg13g2_fill_1 FILLER_75_479 ();
 sg13g2_decap_8 FILLER_75_489 ();
 sg13g2_decap_8 FILLER_75_496 ();
 sg13g2_decap_8 FILLER_75_503 ();
 sg13g2_fill_2 FILLER_75_510 ();
 sg13g2_decap_8 FILLER_75_516 ();
 sg13g2_decap_4 FILLER_75_523 ();
 sg13g2_decap_8 FILLER_75_553 ();
 sg13g2_fill_2 FILLER_75_560 ();
 sg13g2_fill_1 FILLER_75_562 ();
 sg13g2_decap_8 FILLER_75_589 ();
 sg13g2_fill_2 FILLER_75_596 ();
 sg13g2_decap_8 FILLER_75_603 ();
 sg13g2_decap_8 FILLER_75_610 ();
 sg13g2_decap_4 FILLER_75_617 ();
 sg13g2_fill_2 FILLER_75_621 ();
 sg13g2_decap_8 FILLER_75_636 ();
 sg13g2_decap_8 FILLER_75_643 ();
 sg13g2_decap_8 FILLER_75_650 ();
 sg13g2_decap_8 FILLER_75_657 ();
 sg13g2_decap_8 FILLER_75_664 ();
 sg13g2_decap_8 FILLER_75_671 ();
 sg13g2_decap_8 FILLER_75_678 ();
 sg13g2_decap_8 FILLER_75_685 ();
 sg13g2_decap_8 FILLER_75_692 ();
 sg13g2_decap_8 FILLER_75_699 ();
 sg13g2_decap_8 FILLER_75_706 ();
 sg13g2_decap_8 FILLER_75_713 ();
 sg13g2_decap_8 FILLER_75_720 ();
 sg13g2_decap_8 FILLER_75_727 ();
 sg13g2_decap_8 FILLER_75_734 ();
 sg13g2_decap_8 FILLER_75_741 ();
 sg13g2_decap_8 FILLER_75_748 ();
 sg13g2_decap_8 FILLER_75_755 ();
 sg13g2_decap_8 FILLER_75_762 ();
 sg13g2_decap_8 FILLER_75_769 ();
 sg13g2_decap_8 FILLER_75_776 ();
 sg13g2_decap_8 FILLER_75_783 ();
 sg13g2_decap_8 FILLER_75_790 ();
 sg13g2_decap_8 FILLER_75_797 ();
 sg13g2_decap_8 FILLER_75_804 ();
 sg13g2_decap_8 FILLER_75_811 ();
 sg13g2_decap_8 FILLER_75_818 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_839 ();
 sg13g2_decap_8 FILLER_75_846 ();
 sg13g2_decap_8 FILLER_75_853 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_93 ();
 sg13g2_fill_1 FILLER_76_103 ();
 sg13g2_decap_4 FILLER_76_114 ();
 sg13g2_fill_1 FILLER_76_118 ();
 sg13g2_decap_8 FILLER_76_123 ();
 sg13g2_decap_8 FILLER_76_130 ();
 sg13g2_fill_2 FILLER_76_137 ();
 sg13g2_fill_1 FILLER_76_144 ();
 sg13g2_decap_8 FILLER_76_171 ();
 sg13g2_fill_1 FILLER_76_178 ();
 sg13g2_decap_8 FILLER_76_187 ();
 sg13g2_fill_1 FILLER_76_194 ();
 sg13g2_decap_4 FILLER_76_207 ();
 sg13g2_decap_4 FILLER_76_226 ();
 sg13g2_fill_1 FILLER_76_230 ();
 sg13g2_decap_8 FILLER_76_244 ();
 sg13g2_fill_2 FILLER_76_251 ();
 sg13g2_decap_8 FILLER_76_257 ();
 sg13g2_decap_8 FILLER_76_264 ();
 sg13g2_fill_2 FILLER_76_281 ();
 sg13g2_fill_2 FILLER_76_302 ();
 sg13g2_fill_1 FILLER_76_304 ();
 sg13g2_decap_4 FILLER_76_313 ();
 sg13g2_fill_1 FILLER_76_317 ();
 sg13g2_fill_2 FILLER_76_323 ();
 sg13g2_decap_4 FILLER_76_330 ();
 sg13g2_fill_2 FILLER_76_334 ();
 sg13g2_decap_4 FILLER_76_370 ();
 sg13g2_fill_2 FILLER_76_374 ();
 sg13g2_decap_8 FILLER_76_403 ();
 sg13g2_fill_1 FILLER_76_410 ();
 sg13g2_decap_4 FILLER_76_416 ();
 sg13g2_fill_1 FILLER_76_420 ();
 sg13g2_fill_1 FILLER_76_425 ();
 sg13g2_decap_8 FILLER_76_430 ();
 sg13g2_fill_2 FILLER_76_437 ();
 sg13g2_fill_1 FILLER_76_439 ();
 sg13g2_fill_2 FILLER_76_460 ();
 sg13g2_fill_1 FILLER_76_462 ();
 sg13g2_decap_8 FILLER_76_478 ();
 sg13g2_decap_8 FILLER_76_497 ();
 sg13g2_decap_8 FILLER_76_504 ();
 sg13g2_decap_8 FILLER_76_511 ();
 sg13g2_decap_8 FILLER_76_518 ();
 sg13g2_decap_8 FILLER_76_525 ();
 sg13g2_decap_8 FILLER_76_532 ();
 sg13g2_decap_8 FILLER_76_539 ();
 sg13g2_decap_8 FILLER_76_546 ();
 sg13g2_decap_8 FILLER_76_553 ();
 sg13g2_decap_8 FILLER_76_560 ();
 sg13g2_decap_8 FILLER_76_567 ();
 sg13g2_decap_8 FILLER_76_578 ();
 sg13g2_decap_8 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_592 ();
 sg13g2_decap_4 FILLER_76_599 ();
 sg13g2_fill_1 FILLER_76_603 ();
 sg13g2_decap_8 FILLER_76_630 ();
 sg13g2_decap_8 FILLER_76_637 ();
 sg13g2_decap_8 FILLER_76_644 ();
 sg13g2_decap_8 FILLER_76_651 ();
 sg13g2_decap_8 FILLER_76_658 ();
 sg13g2_decap_8 FILLER_76_665 ();
 sg13g2_decap_8 FILLER_76_672 ();
 sg13g2_decap_8 FILLER_76_679 ();
 sg13g2_decap_8 FILLER_76_686 ();
 sg13g2_decap_8 FILLER_76_693 ();
 sg13g2_decap_8 FILLER_76_700 ();
 sg13g2_decap_8 FILLER_76_707 ();
 sg13g2_decap_8 FILLER_76_714 ();
 sg13g2_decap_8 FILLER_76_721 ();
 sg13g2_decap_8 FILLER_76_728 ();
 sg13g2_decap_8 FILLER_76_735 ();
 sg13g2_decap_8 FILLER_76_742 ();
 sg13g2_decap_8 FILLER_76_749 ();
 sg13g2_decap_8 FILLER_76_756 ();
 sg13g2_decap_8 FILLER_76_763 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_decap_8 FILLER_76_791 ();
 sg13g2_decap_8 FILLER_76_798 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_8 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_decap_8 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_76_847 ();
 sg13g2_decap_8 FILLER_76_854 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_4 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_95 ();
 sg13g2_fill_2 FILLER_77_107 ();
 sg13g2_fill_1 FILLER_77_135 ();
 sg13g2_fill_2 FILLER_77_141 ();
 sg13g2_fill_1 FILLER_77_143 ();
 sg13g2_fill_1 FILLER_77_153 ();
 sg13g2_decap_4 FILLER_77_171 ();
 sg13g2_fill_1 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_199 ();
 sg13g2_decap_4 FILLER_77_206 ();
 sg13g2_fill_1 FILLER_77_210 ();
 sg13g2_fill_2 FILLER_77_226 ();
 sg13g2_fill_1 FILLER_77_228 ();
 sg13g2_decap_8 FILLER_77_235 ();
 sg13g2_fill_2 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_274 ();
 sg13g2_decap_8 FILLER_77_283 ();
 sg13g2_fill_2 FILLER_77_290 ();
 sg13g2_decap_8 FILLER_77_316 ();
 sg13g2_fill_1 FILLER_77_323 ();
 sg13g2_fill_2 FILLER_77_337 ();
 sg13g2_decap_4 FILLER_77_349 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_364 ();
 sg13g2_decap_4 FILLER_77_371 ();
 sg13g2_fill_2 FILLER_77_375 ();
 sg13g2_fill_2 FILLER_77_386 ();
 sg13g2_decap_4 FILLER_77_392 ();
 sg13g2_fill_1 FILLER_77_404 ();
 sg13g2_decap_8 FILLER_77_410 ();
 sg13g2_decap_8 FILLER_77_431 ();
 sg13g2_decap_4 FILLER_77_456 ();
 sg13g2_fill_2 FILLER_77_460 ();
 sg13g2_fill_2 FILLER_77_476 ();
 sg13g2_decap_8 FILLER_77_484 ();
 sg13g2_decap_8 FILLER_77_491 ();
 sg13g2_decap_8 FILLER_77_498 ();
 sg13g2_decap_8 FILLER_77_505 ();
 sg13g2_decap_8 FILLER_77_512 ();
 sg13g2_decap_8 FILLER_77_519 ();
 sg13g2_decap_8 FILLER_77_526 ();
 sg13g2_decap_8 FILLER_77_533 ();
 sg13g2_decap_8 FILLER_77_540 ();
 sg13g2_decap_8 FILLER_77_547 ();
 sg13g2_decap_8 FILLER_77_554 ();
 sg13g2_decap_8 FILLER_77_561 ();
 sg13g2_decap_8 FILLER_77_568 ();
 sg13g2_decap_8 FILLER_77_575 ();
 sg13g2_decap_8 FILLER_77_582 ();
 sg13g2_decap_8 FILLER_77_589 ();
 sg13g2_decap_8 FILLER_77_596 ();
 sg13g2_decap_8 FILLER_77_603 ();
 sg13g2_decap_4 FILLER_77_610 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_decap_8 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_632 ();
 sg13g2_decap_8 FILLER_77_639 ();
 sg13g2_decap_8 FILLER_77_646 ();
 sg13g2_decap_8 FILLER_77_653 ();
 sg13g2_decap_8 FILLER_77_660 ();
 sg13g2_decap_8 FILLER_77_667 ();
 sg13g2_decap_8 FILLER_77_674 ();
 sg13g2_decap_8 FILLER_77_681 ();
 sg13g2_decap_8 FILLER_77_688 ();
 sg13g2_decap_8 FILLER_77_695 ();
 sg13g2_decap_8 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_709 ();
 sg13g2_decap_8 FILLER_77_716 ();
 sg13g2_decap_8 FILLER_77_723 ();
 sg13g2_decap_8 FILLER_77_730 ();
 sg13g2_decap_8 FILLER_77_737 ();
 sg13g2_decap_8 FILLER_77_744 ();
 sg13g2_decap_8 FILLER_77_751 ();
 sg13g2_decap_8 FILLER_77_758 ();
 sg13g2_decap_8 FILLER_77_765 ();
 sg13g2_decap_8 FILLER_77_772 ();
 sg13g2_decap_8 FILLER_77_779 ();
 sg13g2_decap_8 FILLER_77_786 ();
 sg13g2_decap_8 FILLER_77_793 ();
 sg13g2_decap_8 FILLER_77_800 ();
 sg13g2_decap_8 FILLER_77_807 ();
 sg13g2_decap_8 FILLER_77_814 ();
 sg13g2_decap_8 FILLER_77_821 ();
 sg13g2_decap_8 FILLER_77_828 ();
 sg13g2_decap_8 FILLER_77_835 ();
 sg13g2_decap_8 FILLER_77_842 ();
 sg13g2_decap_8 FILLER_77_849 ();
 sg13g2_decap_4 FILLER_77_856 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_4 FILLER_78_77 ();
 sg13g2_fill_2 FILLER_78_81 ();
 sg13g2_decap_8 FILLER_78_109 ();
 sg13g2_decap_8 FILLER_78_116 ();
 sg13g2_decap_4 FILLER_78_123 ();
 sg13g2_fill_1 FILLER_78_138 ();
 sg13g2_fill_2 FILLER_78_144 ();
 sg13g2_fill_1 FILLER_78_146 ();
 sg13g2_fill_1 FILLER_78_156 ();
 sg13g2_decap_8 FILLER_78_162 ();
 sg13g2_decap_8 FILLER_78_169 ();
 sg13g2_decap_8 FILLER_78_176 ();
 sg13g2_fill_2 FILLER_78_183 ();
 sg13g2_fill_1 FILLER_78_185 ();
 sg13g2_fill_1 FILLER_78_195 ();
 sg13g2_decap_8 FILLER_78_206 ();
 sg13g2_decap_4 FILLER_78_213 ();
 sg13g2_fill_1 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_229 ();
 sg13g2_decap_8 FILLER_78_236 ();
 sg13g2_decap_4 FILLER_78_243 ();
 sg13g2_fill_1 FILLER_78_247 ();
 sg13g2_decap_8 FILLER_78_254 ();
 sg13g2_decap_8 FILLER_78_261 ();
 sg13g2_fill_2 FILLER_78_268 ();
 sg13g2_fill_1 FILLER_78_270 ();
 sg13g2_fill_2 FILLER_78_284 ();
 sg13g2_fill_1 FILLER_78_286 ();
 sg13g2_decap_8 FILLER_78_293 ();
 sg13g2_fill_2 FILLER_78_300 ();
 sg13g2_decap_8 FILLER_78_307 ();
 sg13g2_decap_4 FILLER_78_314 ();
 sg13g2_fill_1 FILLER_78_318 ();
 sg13g2_decap_4 FILLER_78_338 ();
 sg13g2_fill_1 FILLER_78_342 ();
 sg13g2_decap_8 FILLER_78_372 ();
 sg13g2_decap_4 FILLER_78_379 ();
 sg13g2_fill_1 FILLER_78_383 ();
 sg13g2_fill_2 FILLER_78_399 ();
 sg13g2_fill_1 FILLER_78_401 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_428 ();
 sg13g2_decap_4 FILLER_78_435 ();
 sg13g2_fill_2 FILLER_78_439 ();
 sg13g2_fill_2 FILLER_78_452 ();
 sg13g2_decap_4 FILLER_78_467 ();
 sg13g2_decap_8 FILLER_78_480 ();
 sg13g2_decap_8 FILLER_78_487 ();
 sg13g2_decap_8 FILLER_78_494 ();
 sg13g2_decap_8 FILLER_78_501 ();
 sg13g2_decap_8 FILLER_78_508 ();
 sg13g2_decap_8 FILLER_78_515 ();
 sg13g2_decap_8 FILLER_78_522 ();
 sg13g2_decap_8 FILLER_78_529 ();
 sg13g2_decap_8 FILLER_78_536 ();
 sg13g2_decap_8 FILLER_78_543 ();
 sg13g2_decap_8 FILLER_78_550 ();
 sg13g2_decap_8 FILLER_78_557 ();
 sg13g2_decap_8 FILLER_78_564 ();
 sg13g2_decap_8 FILLER_78_571 ();
 sg13g2_decap_8 FILLER_78_578 ();
 sg13g2_decap_8 FILLER_78_585 ();
 sg13g2_decap_8 FILLER_78_592 ();
 sg13g2_decap_8 FILLER_78_599 ();
 sg13g2_decap_8 FILLER_78_606 ();
 sg13g2_decap_8 FILLER_78_613 ();
 sg13g2_decap_8 FILLER_78_620 ();
 sg13g2_decap_8 FILLER_78_627 ();
 sg13g2_decap_8 FILLER_78_634 ();
 sg13g2_decap_8 FILLER_78_641 ();
 sg13g2_decap_8 FILLER_78_648 ();
 sg13g2_decap_8 FILLER_78_655 ();
 sg13g2_decap_8 FILLER_78_662 ();
 sg13g2_decap_8 FILLER_78_669 ();
 sg13g2_decap_8 FILLER_78_676 ();
 sg13g2_decap_8 FILLER_78_683 ();
 sg13g2_decap_8 FILLER_78_690 ();
 sg13g2_decap_8 FILLER_78_697 ();
 sg13g2_decap_8 FILLER_78_704 ();
 sg13g2_decap_8 FILLER_78_711 ();
 sg13g2_decap_8 FILLER_78_718 ();
 sg13g2_decap_8 FILLER_78_725 ();
 sg13g2_decap_8 FILLER_78_732 ();
 sg13g2_decap_8 FILLER_78_739 ();
 sg13g2_decap_8 FILLER_78_746 ();
 sg13g2_decap_8 FILLER_78_753 ();
 sg13g2_decap_8 FILLER_78_760 ();
 sg13g2_decap_8 FILLER_78_767 ();
 sg13g2_decap_8 FILLER_78_774 ();
 sg13g2_decap_8 FILLER_78_781 ();
 sg13g2_decap_8 FILLER_78_788 ();
 sg13g2_decap_8 FILLER_78_795 ();
 sg13g2_decap_8 FILLER_78_802 ();
 sg13g2_decap_8 FILLER_78_809 ();
 sg13g2_decap_8 FILLER_78_816 ();
 sg13g2_decap_8 FILLER_78_823 ();
 sg13g2_decap_8 FILLER_78_830 ();
 sg13g2_decap_8 FILLER_78_837 ();
 sg13g2_decap_8 FILLER_78_844 ();
 sg13g2_decap_8 FILLER_78_851 ();
 sg13g2_decap_4 FILLER_78_858 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_91 ();
 sg13g2_fill_1 FILLER_79_93 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_fill_2 FILLER_79_105 ();
 sg13g2_fill_1 FILLER_79_107 ();
 sg13g2_decap_8 FILLER_79_160 ();
 sg13g2_decap_8 FILLER_79_167 ();
 sg13g2_fill_1 FILLER_79_174 ();
 sg13g2_decap_8 FILLER_79_227 ();
 sg13g2_decap_4 FILLER_79_234 ();
 sg13g2_decap_4 FILLER_79_268 ();
 sg13g2_fill_1 FILLER_79_272 ();
 sg13g2_fill_2 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_289 ();
 sg13g2_fill_2 FILLER_79_297 ();
 sg13g2_fill_2 FILLER_79_310 ();
 sg13g2_fill_2 FILLER_79_320 ();
 sg13g2_fill_1 FILLER_79_322 ();
 sg13g2_fill_1 FILLER_79_339 ();
 sg13g2_fill_2 FILLER_79_351 ();
 sg13g2_fill_1 FILLER_79_353 ();
 sg13g2_fill_2 FILLER_79_359 ();
 sg13g2_fill_2 FILLER_79_370 ();
 sg13g2_fill_1 FILLER_79_372 ();
 sg13g2_fill_2 FILLER_79_396 ();
 sg13g2_fill_1 FILLER_79_398 ();
 sg13g2_fill_1 FILLER_79_417 ();
 sg13g2_decap_4 FILLER_79_429 ();
 sg13g2_fill_1 FILLER_79_441 ();
 sg13g2_fill_2 FILLER_79_450 ();
 sg13g2_fill_1 FILLER_79_452 ();
 sg13g2_fill_1 FILLER_79_463 ();
 sg13g2_decap_8 FILLER_79_484 ();
 sg13g2_decap_8 FILLER_79_491 ();
 sg13g2_decap_8 FILLER_79_498 ();
 sg13g2_decap_8 FILLER_79_505 ();
 sg13g2_decap_8 FILLER_79_512 ();
 sg13g2_decap_8 FILLER_79_519 ();
 sg13g2_decap_8 FILLER_79_526 ();
 sg13g2_decap_8 FILLER_79_533 ();
 sg13g2_decap_8 FILLER_79_540 ();
 sg13g2_decap_8 FILLER_79_547 ();
 sg13g2_decap_8 FILLER_79_554 ();
 sg13g2_decap_8 FILLER_79_561 ();
 sg13g2_decap_8 FILLER_79_568 ();
 sg13g2_decap_8 FILLER_79_575 ();
 sg13g2_decap_8 FILLER_79_582 ();
 sg13g2_decap_8 FILLER_79_589 ();
 sg13g2_decap_8 FILLER_79_596 ();
 sg13g2_decap_8 FILLER_79_603 ();
 sg13g2_decap_8 FILLER_79_610 ();
 sg13g2_decap_8 FILLER_79_617 ();
 sg13g2_decap_8 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_631 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_659 ();
 sg13g2_decap_8 FILLER_79_666 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_687 ();
 sg13g2_decap_8 FILLER_79_694 ();
 sg13g2_decap_8 FILLER_79_701 ();
 sg13g2_decap_8 FILLER_79_708 ();
 sg13g2_decap_8 FILLER_79_715 ();
 sg13g2_decap_8 FILLER_79_722 ();
 sg13g2_decap_8 FILLER_79_729 ();
 sg13g2_decap_8 FILLER_79_736 ();
 sg13g2_decap_8 FILLER_79_743 ();
 sg13g2_decap_8 FILLER_79_750 ();
 sg13g2_decap_8 FILLER_79_757 ();
 sg13g2_decap_8 FILLER_79_764 ();
 sg13g2_decap_8 FILLER_79_771 ();
 sg13g2_decap_8 FILLER_79_778 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_fill_1 FILLER_80_140 ();
 sg13g2_fill_2 FILLER_80_149 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_fill_2 FILLER_80_180 ();
 sg13g2_fill_2 FILLER_80_191 ();
 sg13g2_fill_1 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_4 FILLER_80_206 ();
 sg13g2_fill_2 FILLER_80_210 ();
 sg13g2_decap_8 FILLER_80_216 ();
 sg13g2_decap_8 FILLER_80_223 ();
 sg13g2_decap_8 FILLER_80_230 ();
 sg13g2_decap_8 FILLER_80_237 ();
 sg13g2_decap_4 FILLER_80_244 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_decap_4 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_295 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_fill_2 FILLER_80_315 ();
 sg13g2_fill_2 FILLER_80_322 ();
 sg13g2_fill_1 FILLER_80_324 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_347 ();
 sg13g2_fill_2 FILLER_80_351 ();
 sg13g2_decap_8 FILLER_80_369 ();
 sg13g2_decap_8 FILLER_80_376 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_407 ();
 sg13g2_fill_1 FILLER_80_409 ();
 sg13g2_fill_1 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_425 ();
 sg13g2_decap_8 FILLER_80_432 ();
 sg13g2_fill_2 FILLER_80_439 ();
 sg13g2_decap_8 FILLER_80_454 ();
 sg13g2_decap_8 FILLER_80_461 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_536 ();
 sg13g2_decap_8 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_550 ();
 sg13g2_decap_8 FILLER_80_557 ();
 sg13g2_decap_8 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_decap_8 FILLER_80_851 ();
 sg13g2_decap_4 FILLER_80_858 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net164;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule
